module fake_netlist_6_3150_n_2917 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_356, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2917);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_356;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2917;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_1009;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_1371;
wire n_873;
wire n_1285;
wire n_2886;
wire n_1985;
wire n_2838;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_943;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_638;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_699;
wire n_1986;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_1801;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2810;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1317;
wire n_1082;
wire n_2733;
wire n_2824;
wire n_593;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_738;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_705;
wire n_2134;
wire n_1176;
wire n_1004;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_777;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_745;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_623;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_1837;
wire n_831;
wire n_2218;
wire n_2788;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_642;
wire n_995;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_1390;
wire n_906;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_956;
wire n_2276;
wire n_960;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_621;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_609;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2900;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2904;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_1352;
wire n_579;
wire n_2789;
wire n_2872;
wire n_937;
wire n_2257;
wire n_2017;
wire n_1682;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_1548;
wire n_799;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_737;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_1962;
wire n_1236;
wire n_786;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_2062;
wire n_660;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_817;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_2140;
wire n_988;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_1583;
wire n_832;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1848;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_2906;
wire n_1303;
wire n_761;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_1973;
wire n_708;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_779;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_771;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_1260;
wire n_2055;
wire n_1819;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_2899;
wire n_1322;
wire n_640;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2912;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_562),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_257),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_76),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_353),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_156),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_4),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_515),
.Y(n_581)
);

CKINVDCx14_ASAP7_75t_R g582 ( 
.A(n_81),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_469),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_423),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_496),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_218),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_216),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_528),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_509),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_524),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_507),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_541),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_290),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_315),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_469),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_341),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_84),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_495),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_516),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_57),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_182),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_419),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_434),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_226),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_431),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_283),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_81),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_218),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_470),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_527),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_305),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_450),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_442),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_177),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_471),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_388),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_355),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_46),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_129),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_103),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_129),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_19),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_153),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_280),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_64),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_310),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_549),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_205),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_354),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_349),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_342),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_209),
.Y(n_632)
);

CKINVDCx16_ASAP7_75t_R g633 ( 
.A(n_35),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_573),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_530),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_58),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_490),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_137),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_446),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_316),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_192),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_220),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_430),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_185),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_216),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_211),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_138),
.Y(n_647)
);

CKINVDCx16_ASAP7_75t_R g648 ( 
.A(n_445),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_108),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_539),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_517),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_371),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_482),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_137),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_396),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_21),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_223),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_332),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_538),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_58),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_60),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_135),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_393),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_330),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_341),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_447),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_0),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_540),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_458),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_520),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_30),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_421),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_339),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_570),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_207),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_78),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_401),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_574),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_99),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_310),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_458),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_143),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_298),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_15),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_211),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_90),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_56),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_428),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_68),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_429),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_173),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_307),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_16),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_31),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_326),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_253),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_462),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_39),
.Y(n_698)
);

CKINVDCx16_ASAP7_75t_R g699 ( 
.A(n_550),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_367),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_552),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_365),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_112),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_551),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_105),
.Y(n_705)
);

BUFx2_ASAP7_75t_SL g706 ( 
.A(n_449),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_367),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_489),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_365),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_111),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_464),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_174),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_190),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_510),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_460),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_560),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_99),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_240),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_252),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_478),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_477),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_340),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_555),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_74),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_497),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_486),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_31),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_499),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_9),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_361),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_565),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_330),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_559),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_231),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_495),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_571),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_71),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_180),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_494),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_373),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_423),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_513),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_345),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_475),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_273),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_312),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_473),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_163),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_198),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_172),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_88),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_449),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_500),
.Y(n_753)
);

BUFx5_ASAP7_75t_L g754 ( 
.A(n_516),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_299),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_521),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_83),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_532),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_405),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_533),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_487),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_167),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_1),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_513),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_368),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_388),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_359),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_389),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_353),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_39),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_55),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_558),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_362),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_436),
.Y(n_774)
);

INVxp33_ASAP7_75t_SL g775 ( 
.A(n_27),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_57),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_510),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_38),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_202),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_375),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_142),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_42),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_443),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_518),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_321),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_383),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_52),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_186),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_65),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_297),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_564),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_337),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_425),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_548),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_369),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_501),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_143),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_107),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_213),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_136),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_561),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_523),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_148),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_501),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_521),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_404),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_22),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_511),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_303),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_273),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_87),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_556),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_123),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_68),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_360),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_17),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_419),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_72),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_442),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_254),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_94),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_242),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_519),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_290),
.Y(n_824)
);

BUFx5_ASAP7_75t_L g825 ( 
.A(n_284),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_300),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_529),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_56),
.Y(n_828)
);

CKINVDCx14_ASAP7_75t_R g829 ( 
.A(n_483),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_488),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_446),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_110),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_404),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_308),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_441),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_306),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_212),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_277),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_491),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_85),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_254),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_547),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_140),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_535),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_144),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_567),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_142),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_396),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_269),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_485),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_506),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_450),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_505),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_363),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_139),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_161),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_536),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_5),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_206),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_52),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_544),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_493),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_363),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_54),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_546),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_127),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_563),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_379),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_22),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_82),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_122),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_514),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_277),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_237),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_515),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_8),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_566),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_20),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_160),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_110),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_477),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_74),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_468),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_398),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_299),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_3),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_355),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_21),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_500),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_84),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_401),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_235),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_219),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_456),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_239),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_207),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_160),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_118),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_148),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_232),
.Y(n_900)
);

HB1xp67_ASAP7_75t_SL g901 ( 
.A(n_116),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_12),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_487),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_471),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_157),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_537),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_508),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_75),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_489),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_305),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_455),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_45),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_542),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_178),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_30),
.Y(n_915)
);

BUFx2_ASAP7_75t_SL g916 ( 
.A(n_153),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_306),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_189),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_190),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_204),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_569),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_543),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_29),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_368),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_545),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_411),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_452),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_534),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_40),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_173),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_184),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_152),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_102),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_251),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_320),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_260),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_83),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_498),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_44),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_172),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_93),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_17),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_270),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_152),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_301),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_504),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_395),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_104),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_381),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_337),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_175),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_436),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_553),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_409),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_470),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_531),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_333),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_10),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_161),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_525),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_287),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_42),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_557),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_511),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_106),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_59),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_335),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_300),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_61),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_9),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_263),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_145),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_526),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_492),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_522),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_473),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_505),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_512),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_251),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_209),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_86),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_526),
.Y(n_982)
);

CKINVDCx14_ASAP7_75t_R g983 ( 
.A(n_502),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_345),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_45),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_5),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_302),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_360),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_233),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_274),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_315),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_568),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_75),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_400),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_435),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_572),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_503),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_498),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_288),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_200),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_476),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_53),
.Y(n_1002)
);

BUFx2_ASAP7_75t_R g1003 ( 
.A(n_393),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_425),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_312),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_114),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_236),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_28),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_295),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_70),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_554),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_72),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_85),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_582),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_754),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_754),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_754),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_581),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_754),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_754),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_592),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_581),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_616),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_754),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_754),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_754),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_668),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_754),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_825),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_825),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_825),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_825),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_829),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_825),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_825),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_825),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_825),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_825),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_657),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_983),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_616),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_633),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_633),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_914),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_914),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_704),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_877),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_704),
.Y(n_1048)
);

INVxp67_ASAP7_75t_SL g1049 ( 
.A(n_635),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_648),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_716),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_648),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_658),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_992),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_716),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_723),
.Y(n_1056)
);

BUFx2_ASAP7_75t_SL g1057 ( 
.A(n_791),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_723),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_1011),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_760),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_760),
.Y(n_1061)
);

INVxp33_ASAP7_75t_SL g1062 ( 
.A(n_700),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_794),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_658),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_755),
.Y(n_1065)
);

INVxp67_ASAP7_75t_L g1066 ( 
.A(n_752),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_794),
.Y(n_1067)
);

INVxp67_ASAP7_75t_SL g1068 ( 
.A(n_658),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_842),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_842),
.Y(n_1070)
);

CKINVDCx16_ASAP7_75t_R g1071 ( 
.A(n_755),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_857),
.Y(n_1072)
);

CKINVDCx16_ASAP7_75t_R g1073 ( 
.A(n_810),
.Y(n_1073)
);

INVxp33_ASAP7_75t_SL g1074 ( 
.A(n_809),
.Y(n_1074)
);

INVxp33_ASAP7_75t_SL g1075 ( 
.A(n_706),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_857),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_913),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_810),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_658),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_657),
.Y(n_1080)
);

INVxp67_ASAP7_75t_SL g1081 ( 
.A(n_657),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_913),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_921),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_921),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_922),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_657),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_657),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_901),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_1042),
.Y(n_1089)
);

AND2x2_ASAP7_75t_SL g1090 ( 
.A(n_1021),
.B(n_699),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1080),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1039),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1080),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1039),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1086),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_1021),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_1042),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1018),
.A2(n_606),
.B1(n_626),
.B2(n_625),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1081),
.B(n_657),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_1053),
.B(n_791),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_1021),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1086),
.Y(n_1102)
);

INVx5_ASAP7_75t_L g1103 ( 
.A(n_1021),
.Y(n_1103)
);

XNOR2xp5_ASAP7_75t_L g1104 ( 
.A(n_1043),
.B(n_1050),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1087),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_1021),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1053),
.B(n_865),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1087),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1068),
.B(n_672),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1043),
.Y(n_1110)
);

CKINVDCx16_ASAP7_75t_R g1111 ( 
.A(n_1071),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_1023),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_1024),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1057),
.B(n_672),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1064),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_1064),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1027),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1015),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1057),
.B(n_672),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1024),
.A2(n_592),
.B(n_922),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1016),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1025),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_1047),
.Y(n_1123)
);

CKINVDCx6p67_ASAP7_75t_R g1124 ( 
.A(n_1073),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1025),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1017),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1026),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1079),
.Y(n_1128)
);

CKINVDCx11_ASAP7_75t_R g1129 ( 
.A(n_1054),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1019),
.B(n_672),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1079),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1026),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1020),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1062),
.A2(n_1002),
.B1(n_664),
.B2(n_671),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1028),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_1056),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1028),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1056),
.B(n_865),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_1029),
.Y(n_1139)
);

BUFx8_ASAP7_75t_L g1140 ( 
.A(n_1022),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1029),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1059),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1030),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_1030),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1031),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1031),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1050),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1046),
.B(n_615),
.Y(n_1148)
);

NOR2x1_ASAP7_75t_L g1149 ( 
.A(n_1032),
.B(n_963),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1032),
.B(n_963),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1123),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_R g1152 ( 
.A(n_1117),
.B(n_1014),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_1129),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1142),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1111),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_1111),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1110),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1124),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_R g1159 ( 
.A(n_1124),
.B(n_1014),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1124),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1140),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1132),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1140),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1091),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1140),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1110),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1109),
.B(n_1048),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1140),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1112),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1112),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_1104),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1104),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1091),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1091),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1089),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1089),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1093),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1093),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1097),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1097),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1147),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_1147),
.Y(n_1182)
);

BUFx10_ASAP7_75t_L g1183 ( 
.A(n_1090),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_R g1184 ( 
.A(n_1090),
.B(n_1033),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1093),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_1134),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1132),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1118),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1090),
.B(n_1109),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1099),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1118),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1118),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1098),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1121),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1121),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_1134),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_R g1197 ( 
.A(n_1114),
.B(n_1033),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1121),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1126),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_R g1200 ( 
.A(n_1114),
.B(n_1040),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1094),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1098),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_1119),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_1119),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1096),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1138),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1150),
.B(n_1070),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1126),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1190),
.B(n_1139),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_1207),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1162),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1152),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1207),
.Y(n_1213)
);

AO22x2_ASAP7_75t_L g1214 ( 
.A1(n_1189),
.A2(n_1044),
.B1(n_1045),
.B2(n_918),
.Y(n_1214)
);

AND2x6_ASAP7_75t_L g1215 ( 
.A(n_1190),
.B(n_1150),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1207),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1164),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1164),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1207),
.Y(n_1219)
);

INVx5_ASAP7_75t_L g1220 ( 
.A(n_1205),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1167),
.B(n_1138),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1173),
.Y(n_1222)
);

BUFx10_ASAP7_75t_L g1223 ( 
.A(n_1158),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1205),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1151),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1167),
.B(n_1150),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1187),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_1158),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1154),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1203),
.B(n_1052),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1167),
.B(n_1139),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1201),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1204),
.A2(n_1150),
.B1(n_1138),
.B2(n_1139),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1173),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1170),
.B(n_1138),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1201),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1206),
.B(n_699),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1174),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1155),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1169),
.B(n_1052),
.Y(n_1240)
);

OR2x6_ASAP7_75t_L g1241 ( 
.A(n_1163),
.B(n_706),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1183),
.A2(n_1150),
.B1(n_1139),
.B2(n_1062),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1174),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1170),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1177),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1183),
.A2(n_1074),
.B1(n_1149),
.B2(n_1049),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1177),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1205),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1206),
.B(n_1065),
.Y(n_1249)
);

INVxp67_ASAP7_75t_SL g1250 ( 
.A(n_1188),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1191),
.B(n_1148),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1183),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1192),
.B(n_1148),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1178),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1197),
.B(n_1148),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1181),
.B(n_1065),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1178),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1194),
.B(n_1113),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1195),
.B(n_1100),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1198),
.B(n_1199),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1208),
.B(n_1113),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1184),
.B(n_1088),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1157),
.B(n_1078),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1200),
.B(n_1040),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1185),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1159),
.B(n_1075),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1185),
.B(n_1100),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1166),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1193),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1163),
.B(n_1100),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1193),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1154),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1153),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1182),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1175),
.B(n_1113),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1175),
.B(n_1113),
.Y(n_1276)
);

AND2x6_ASAP7_75t_L g1277 ( 
.A(n_1161),
.B(n_1149),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1176),
.Y(n_1278)
);

BUFx10_ASAP7_75t_L g1279 ( 
.A(n_1160),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1176),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1179),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1179),
.B(n_1075),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1156),
.B(n_1100),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1180),
.B(n_1127),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1180),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1202),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1244),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1225),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1221),
.B(n_1127),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1255),
.B(n_1160),
.Y(n_1290)
);

NAND2xp33_ASAP7_75t_SL g1291 ( 
.A(n_1212),
.B(n_1161),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1274),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1226),
.A2(n_622),
.B1(n_647),
.B2(n_610),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1216),
.B(n_1165),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1231),
.A2(n_1103),
.B(n_1096),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1225),
.B(n_1022),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1221),
.B(n_1211),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1251),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1217),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1235),
.B(n_1078),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1269),
.B(n_1074),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1235),
.B(n_1041),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_L g1303 ( 
.A(n_1215),
.B(n_1165),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1269),
.B(n_1186),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1217),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1251),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1218),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1255),
.B(n_1066),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1213),
.B(n_1168),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1244),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1211),
.B(n_1127),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1251),
.B(n_1127),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1218),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1226),
.A2(n_1196),
.B1(n_1126),
.B2(n_1133),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1253),
.B(n_1099),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1226),
.A2(n_1133),
.B1(n_1168),
.B2(n_1107),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1268),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1219),
.A2(n_1133),
.B1(n_1107),
.B2(n_1100),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1222),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1253),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1213),
.A2(n_1107),
.B1(n_627),
.B2(n_634),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1253),
.B(n_1135),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1209),
.B(n_1135),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1213),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1227),
.B(n_1276),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1213),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1267),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1213),
.B(n_1136),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1222),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1215),
.A2(n_622),
.B1(n_647),
.B2(n_610),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1275),
.B(n_1135),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1268),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1271),
.B(n_775),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1284),
.B(n_1141),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1233),
.A2(n_679),
.B1(n_695),
.B2(n_652),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1267),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1271),
.A2(n_973),
.B(n_885),
.C(n_1130),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1250),
.B(n_1141),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1210),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1274),
.B(n_916),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1234),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1210),
.A2(n_1107),
.B1(n_650),
.B2(n_659),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1210),
.B(n_1136),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1259),
.B(n_1141),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1267),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_1281),
.B(n_1239),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1237),
.B(n_1003),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1215),
.A2(n_1214),
.B1(n_622),
.B2(n_647),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1215),
.A2(n_837),
.B1(n_875),
.B2(n_610),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1242),
.B(n_1136),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1278),
.A2(n_675),
.B1(n_690),
.B2(n_590),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1259),
.B(n_1143),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1281),
.B(n_916),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1259),
.B(n_1143),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1243),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1239),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1282),
.B(n_707),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1234),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1245),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1243),
.B(n_1143),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1245),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1254),
.B(n_1145),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1283),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1254),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1215),
.A2(n_1107),
.B1(n_674),
.B2(n_678),
.Y(n_1365)
);

INVx8_ASAP7_75t_L g1366 ( 
.A(n_1277),
.Y(n_1366)
);

NAND2xp33_ASAP7_75t_L g1367 ( 
.A(n_1215),
.B(n_575),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1286),
.B(n_1172),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1240),
.Y(n_1369)
);

OR2x6_ASAP7_75t_L g1370 ( 
.A(n_1283),
.B(n_590),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1286),
.B(n_1278),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1212),
.Y(n_1372)
);

NOR3xp33_ASAP7_75t_L g1373 ( 
.A(n_1280),
.B(n_1172),
.C(n_702),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1265),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1257),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1252),
.B(n_1136),
.Y(n_1376)
);

INVxp67_ASAP7_75t_SL g1377 ( 
.A(n_1224),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1265),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1257),
.B(n_1145),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1214),
.A2(n_875),
.B1(n_909),
.B2(n_837),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1232),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1236),
.B(n_1145),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1252),
.B(n_1136),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1256),
.B(n_1171),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1252),
.B(n_1136),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1262),
.B(n_712),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1238),
.B(n_1146),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1249),
.B(n_719),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1247),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1325),
.B(n_1246),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1355),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1363),
.B(n_1283),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1297),
.B(n_1214),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1323),
.A2(n_1248),
.B(n_1224),
.Y(n_1394)
);

CKINVDCx10_ASAP7_75t_R g1395 ( 
.A(n_1296),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1308),
.B(n_1280),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1330),
.A2(n_1214),
.B1(n_1285),
.B2(n_1272),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1326),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1364),
.Y(n_1399)
);

OAI21xp33_ASAP7_75t_L g1400 ( 
.A1(n_1388),
.A2(n_1230),
.B(n_1229),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1315),
.B(n_1277),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1324),
.B(n_1277),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1298),
.B(n_1270),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1302),
.B(n_1229),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1326),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1300),
.B(n_1272),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1304),
.A2(n_1277),
.B1(n_1270),
.B2(n_1264),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1292),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1339),
.A2(n_1248),
.B(n_1220),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1375),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1330),
.A2(n_1263),
.B1(n_1241),
.B2(n_764),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1369),
.B(n_1270),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1317),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1369),
.B(n_1279),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1288),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1287),
.B(n_1263),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1333),
.A2(n_1266),
.B(n_1260),
.C(n_1261),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1299),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1324),
.B(n_1277),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1289),
.A2(n_1220),
.B(n_1258),
.Y(n_1420)
);

INVx11_ASAP7_75t_L g1421 ( 
.A(n_1292),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1333),
.B(n_1371),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1331),
.A2(n_1120),
.B(n_1130),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1338),
.A2(n_1220),
.B(n_1103),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1287),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1317),
.Y(n_1426)
);

O2A1O1Ixp5_ASAP7_75t_L g1427 ( 
.A1(n_1350),
.A2(n_1055),
.B(n_1058),
.C(n_1051),
.Y(n_1427)
);

BUFx4f_ASAP7_75t_L g1428 ( 
.A(n_1346),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1326),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1301),
.B(n_1223),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1305),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1334),
.B(n_1277),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1304),
.B(n_1223),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1310),
.B(n_1223),
.Y(n_1434)
);

INVxp67_ASAP7_75t_SL g1435 ( 
.A(n_1326),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1301),
.A2(n_768),
.B(n_883),
.C(n_666),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1344),
.A2(n_1220),
.B(n_1103),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1352),
.A2(n_1220),
.B(n_1103),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1337),
.A2(n_927),
.B(n_896),
.C(n_1241),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1386),
.B(n_1228),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1310),
.B(n_1228),
.Y(n_1441)
);

AOI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1376),
.A2(n_1120),
.B(n_1108),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1354),
.A2(n_1103),
.B(n_1096),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1377),
.A2(n_1103),
.B(n_1096),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1332),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1386),
.B(n_1228),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1377),
.A2(n_1322),
.B(n_1367),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1312),
.A2(n_1103),
.B(n_1096),
.Y(n_1448)
);

BUFx4f_ASAP7_75t_L g1449 ( 
.A(n_1346),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_L g1450 ( 
.A(n_1366),
.B(n_1349),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1357),
.B(n_1368),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1349),
.A2(n_1106),
.B(n_1096),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1307),
.B(n_1146),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1311),
.A2(n_1106),
.B(n_1096),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1343),
.A2(n_1106),
.B(n_1146),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1313),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1319),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1314),
.B(n_1279),
.Y(n_1458)
);

OAI21xp33_ASAP7_75t_L g1459 ( 
.A1(n_1357),
.A2(n_1347),
.B(n_1335),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1290),
.A2(n_1351),
.B(n_1373),
.C(n_1353),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1383),
.A2(n_1106),
.B(n_1101),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1385),
.A2(n_1106),
.B(n_1101),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1329),
.B(n_1116),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1360),
.A2(n_1106),
.B(n_1101),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1348),
.A2(n_1120),
.B(n_1035),
.Y(n_1465)
);

OR2x2_ASAP7_75t_SL g1466 ( 
.A(n_1347),
.B(n_577),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1362),
.A2(n_1106),
.B(n_1122),
.Y(n_1467)
);

AOI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1379),
.A2(n_1108),
.B(n_1092),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1341),
.B(n_1116),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1327),
.A2(n_1125),
.B(n_1122),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1358),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1359),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1384),
.B(n_1279),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1361),
.B(n_1116),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1374),
.Y(n_1475)
);

NOR3xp33_ASAP7_75t_L g1476 ( 
.A(n_1373),
.B(n_1273),
.C(n_646),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1378),
.B(n_1092),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_SL g1478 ( 
.A(n_1372),
.B(n_1273),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1296),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1306),
.B(n_1136),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1320),
.A2(n_1345),
.B1(n_1336),
.B2(n_1309),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1348),
.A2(n_1241),
.B1(n_686),
.B2(n_744),
.Y(n_1482)
);

NOR2xp67_ASAP7_75t_L g1483 ( 
.A(n_1294),
.B(n_701),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1382),
.A2(n_1035),
.B(n_1034),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1381),
.B(n_1122),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1346),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1392),
.B(n_1294),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1391),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1422),
.B(n_1380),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1459),
.B(n_1451),
.Y(n_1490)
);

O2A1O1Ixp5_ASAP7_75t_L g1491 ( 
.A1(n_1458),
.A2(n_1295),
.B(n_1328),
.C(n_1389),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1399),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1460),
.A2(n_1351),
.B(n_1353),
.C(n_1296),
.Y(n_1493)
);

NAND2x1p5_ASAP7_75t_L g1494 ( 
.A(n_1415),
.B(n_1356),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1482),
.A2(n_1293),
.B1(n_1380),
.B2(n_1353),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1397),
.A2(n_1340),
.B(n_1370),
.C(n_1241),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1450),
.A2(n_1303),
.B(n_1366),
.Y(n_1497)
);

AO21x1_ASAP7_75t_L g1498 ( 
.A1(n_1432),
.A2(n_1393),
.B(n_1401),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1398),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1447),
.A2(n_1366),
.B(n_1387),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1410),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1404),
.B(n_1291),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1397),
.A2(n_1340),
.B(n_1370),
.C(n_675),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1396),
.B(n_1370),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1390),
.B(n_1446),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1400),
.A2(n_1316),
.B(n_1365),
.C(n_1342),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1394),
.A2(n_1293),
.B(n_1318),
.Y(n_1507)
);

OR2x6_ASAP7_75t_L g1508 ( 
.A(n_1408),
.B(n_1340),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1398),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1430),
.B(n_1321),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1406),
.B(n_742),
.Y(n_1511)
);

INVx5_ASAP7_75t_L g1512 ( 
.A(n_1398),
.Y(n_1512)
);

AO32x1_ASAP7_75t_L g1513 ( 
.A1(n_1411),
.A2(n_762),
.A3(n_796),
.B1(n_745),
.B2(n_690),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1408),
.B(n_745),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1408),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1431),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1432),
.A2(n_1125),
.B(n_1122),
.Y(n_1517)
);

AOI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1423),
.A2(n_1128),
.B(n_1115),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1418),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_SL g1520 ( 
.A1(n_1417),
.A2(n_796),
.B(n_800),
.C(n_762),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1440),
.B(n_1060),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1420),
.A2(n_1125),
.B(n_1122),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1413),
.B(n_1061),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1393),
.A2(n_782),
.B1(n_784),
.B2(n_774),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1466),
.A2(n_803),
.B1(n_841),
.B2(n_798),
.Y(n_1525)
);

INVx5_ASAP7_75t_L g1526 ( 
.A(n_1405),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1456),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1411),
.A2(n_1407),
.B1(n_1449),
.B2(n_1428),
.Y(n_1528)
);

O2A1O1Ixp33_ASAP7_75t_SL g1529 ( 
.A1(n_1402),
.A2(n_911),
.B(n_918),
.C(n_800),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1419),
.A2(n_1125),
.B(n_1122),
.Y(n_1530)
);

NOR2x1_ASAP7_75t_L g1531 ( 
.A(n_1405),
.B(n_872),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1425),
.Y(n_1532)
);

A2O1A1Ixp33_ASAP7_75t_SL g1533 ( 
.A1(n_1434),
.A2(n_1067),
.B(n_1069),
.C(n_1063),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1421),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1478),
.B(n_890),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1439),
.A2(n_655),
.B(n_722),
.C(n_615),
.Y(n_1536)
);

O2A1O1Ixp5_ASAP7_75t_L g1537 ( 
.A1(n_1433),
.A2(n_1076),
.B(n_1077),
.C(n_1072),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1426),
.B(n_1412),
.Y(n_1538)
);

INVx5_ASAP7_75t_L g1539 ( 
.A(n_1429),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1416),
.B(n_1473),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1465),
.A2(n_1137),
.B(n_1125),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_L g1542 ( 
.A(n_1436),
.B(n_1083),
.C(n_1082),
.Y(n_1542)
);

CKINVDCx6p67_ASAP7_75t_R g1543 ( 
.A(n_1395),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1465),
.A2(n_1137),
.B(n_1125),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1392),
.B(n_1084),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1481),
.A2(n_1428),
.B1(n_1449),
.B2(n_1435),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1457),
.Y(n_1547)
);

O2A1O1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1476),
.A2(n_1414),
.B(n_1479),
.C(n_1441),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1403),
.B(n_1085),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1409),
.A2(n_1137),
.B(n_1144),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_SL g1551 ( 
.A(n_1486),
.B(n_977),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1475),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1445),
.B(n_1486),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1471),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1429),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1403),
.B(n_893),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1472),
.A2(n_919),
.B1(n_946),
.B2(n_934),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1485),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1424),
.A2(n_1137),
.B(n_1144),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1483),
.B(n_624),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1485),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1463),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1463),
.B(n_577),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1477),
.B(n_714),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1484),
.A2(n_1137),
.B(n_1144),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1484),
.A2(n_1137),
.B(n_1144),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1477),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1469),
.B(n_729),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1427),
.B(n_974),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1469),
.B(n_730),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1442),
.A2(n_1128),
.B(n_1115),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1474),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1474),
.A2(n_1453),
.B1(n_1480),
.B2(n_1470),
.Y(n_1573)
);

OR2x4_ASAP7_75t_L g1574 ( 
.A(n_1453),
.B(n_588),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1461),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1437),
.B(n_978),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1468),
.Y(n_1577)
);

BUFx2_ASAP7_75t_SL g1578 ( 
.A(n_1462),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1455),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1452),
.B(n_586),
.Y(n_1580)
);

BUFx12f_ASAP7_75t_L g1581 ( 
.A(n_1464),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_R g1582 ( 
.A(n_1448),
.B(n_731),
.Y(n_1582)
);

NOR2x1_ASAP7_75t_L g1583 ( 
.A(n_1444),
.B(n_615),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1467),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1454),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1443),
.Y(n_1586)
);

A2O1A1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1438),
.A2(n_722),
.B(n_741),
.C(n_655),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1490),
.A2(n_911),
.B1(n_722),
.B2(n_741),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1488),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1532),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1487),
.B(n_655),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1504),
.B(n_1540),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1494),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1508),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1571),
.A2(n_1131),
.B(n_1095),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1508),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1495),
.A2(n_769),
.B1(n_781),
.B2(n_741),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1493),
.B(n_578),
.C(n_576),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1497),
.A2(n_1131),
.B(n_736),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1496),
.A2(n_781),
.B(n_788),
.C(n_769),
.Y(n_1600)
);

O2A1O1Ixp5_ASAP7_75t_L g1601 ( 
.A1(n_1498),
.A2(n_588),
.B(n_600),
.C(n_597),
.Y(n_1601)
);

A2O1A1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1503),
.A2(n_1506),
.B(n_1505),
.C(n_1495),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1564),
.B(n_767),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1500),
.A2(n_1507),
.B(n_1541),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1489),
.A2(n_1095),
.B(n_1094),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1515),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1567),
.B(n_597),
.Y(n_1607)
);

A2O1A1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1528),
.A2(n_781),
.B(n_788),
.C(n_769),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1562),
.B(n_600),
.Y(n_1609)
);

NAND3x1_ASAP7_75t_L g1610 ( 
.A(n_1531),
.B(n_607),
.C(n_601),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1551),
.B(n_733),
.Y(n_1611)
);

OA21x2_ASAP7_75t_L g1612 ( 
.A1(n_1518),
.A2(n_1036),
.B(n_1034),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1522),
.A2(n_1095),
.B(n_1094),
.Y(n_1613)
);

AOI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1530),
.A2(n_1037),
.B(n_1036),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1517),
.A2(n_1105),
.B(n_1102),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_SL g1616 ( 
.A1(n_1528),
.A2(n_875),
.B(n_837),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1535),
.B(n_820),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1544),
.A2(n_772),
.B(n_758),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1487),
.B(n_788),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1508),
.Y(n_1620)
);

AO31x2_ASAP7_75t_L g1621 ( 
.A1(n_1577),
.A2(n_994),
.A3(n_1008),
.B(n_909),
.Y(n_1621)
);

AO32x2_ASAP7_75t_L g1622 ( 
.A1(n_1524),
.A2(n_617),
.A3(n_595),
.B1(n_586),
.B2(n_882),
.Y(n_1622)
);

NOR3xp33_ASAP7_75t_L g1623 ( 
.A(n_1525),
.B(n_853),
.C(n_849),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1546),
.B(n_909),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1501),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1585),
.A2(n_1105),
.B(n_1102),
.Y(n_1626)
);

AO31x2_ASAP7_75t_L g1627 ( 
.A1(n_1586),
.A2(n_1008),
.A3(n_994),
.B(n_602),
.Y(n_1627)
);

AOI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1576),
.A2(n_1038),
.B(n_1037),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1492),
.Y(n_1629)
);

OAI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1573),
.A2(n_1038),
.B(n_1008),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1548),
.A2(n_931),
.B(n_951),
.C(n_882),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1510),
.A2(n_812),
.B(n_801),
.Y(n_1632)
);

NOR4xp25_ASAP7_75t_L g1633 ( 
.A(n_1524),
.B(n_607),
.C(n_611),
.D(n_601),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1568),
.B(n_866),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1565),
.A2(n_846),
.B(n_844),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1516),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1570),
.B(n_910),
.Y(n_1637)
);

BUFx2_ASAP7_75t_R g1638 ( 
.A(n_1511),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1566),
.A2(n_867),
.B(n_861),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1559),
.A2(n_994),
.B(n_613),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1491),
.A2(n_613),
.B(n_611),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1538),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1584),
.A2(n_925),
.B(n_906),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1521),
.B(n_932),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1556),
.B(n_964),
.Y(n_1645)
);

A2O1A1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1536),
.A2(n_931),
.B(n_951),
.C(n_882),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1499),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1554),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1499),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1551),
.B(n_1525),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1520),
.A2(n_953),
.B(n_928),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1553),
.B(n_931),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1579),
.A2(n_996),
.B(n_956),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1550),
.A2(n_628),
.B(n_619),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1569),
.A2(n_1137),
.B(n_739),
.Y(n_1655)
);

NAND3x1_ASAP7_75t_L g1656 ( 
.A(n_1560),
.B(n_628),
.C(n_619),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1563),
.B(n_586),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1583),
.A2(n_1558),
.B(n_1537),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1587),
.A2(n_630),
.B(n_629),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1558),
.A2(n_1547),
.B(n_1580),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1563),
.B(n_579),
.Y(n_1661)
);

CKINVDCx20_ASAP7_75t_R g1662 ( 
.A(n_1543),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1575),
.A2(n_739),
.B(n_602),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1555),
.Y(n_1664)
);

AO31x2_ASAP7_75t_L g1665 ( 
.A1(n_1519),
.A2(n_884),
.A3(n_917),
.B(n_748),
.Y(n_1665)
);

OA21x2_ASAP7_75t_L g1666 ( 
.A1(n_1542),
.A2(n_630),
.B(n_629),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1527),
.A2(n_639),
.B(n_638),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1562),
.A2(n_884),
.B(n_748),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1557),
.A2(n_584),
.B1(n_585),
.B2(n_583),
.C(n_580),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1604),
.A2(n_1529),
.B(n_1502),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1642),
.B(n_1552),
.Y(n_1671)
);

INVx6_ASAP7_75t_L g1672 ( 
.A(n_1593),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1594),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1592),
.B(n_1557),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1629),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1606),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1601),
.A2(n_1542),
.B(n_1545),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1615),
.A2(n_1578),
.B(n_1549),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1650),
.A2(n_1574),
.B1(n_1514),
.B2(n_1523),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1660),
.B(n_1562),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1627),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1614),
.A2(n_1581),
.B(n_1572),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1633),
.B(n_1572),
.Y(n_1683)
);

AO32x2_ASAP7_75t_L g1684 ( 
.A1(n_1597),
.A2(n_1513),
.A3(n_1533),
.B1(n_1534),
.B2(n_1582),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1647),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1630),
.A2(n_1572),
.B(n_639),
.Y(n_1686)
);

OR2x6_ASAP7_75t_L g1687 ( 
.A(n_1624),
.B(n_1514),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1636),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1613),
.A2(n_642),
.B(n_638),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1602),
.A2(n_1513),
.B(n_1512),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1623),
.A2(n_595),
.B1(n_617),
.B2(n_586),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1626),
.A2(n_645),
.B(n_642),
.Y(n_1692)
);

OA21x2_ASAP7_75t_L g1693 ( 
.A1(n_1641),
.A2(n_649),
.B(n_645),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1589),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1625),
.Y(n_1695)
);

AOI221x1_ASAP7_75t_L g1696 ( 
.A1(n_1663),
.A2(n_649),
.B1(n_676),
.B2(n_663),
.C(n_651),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1621),
.Y(n_1697)
);

INVx5_ASAP7_75t_L g1698 ( 
.A(n_1624),
.Y(n_1698)
);

AO21x2_ASAP7_75t_L g1699 ( 
.A1(n_1641),
.A2(n_1513),
.B(n_663),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1600),
.A2(n_1633),
.B(n_1631),
.C(n_1608),
.Y(n_1700)
);

BUFx12f_ASAP7_75t_L g1701 ( 
.A(n_1591),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1596),
.B(n_1526),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1648),
.B(n_1555),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1621),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1598),
.A2(n_1514),
.B(n_1561),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1621),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1598),
.A2(n_980),
.B(n_993),
.C(n_951),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1617),
.A2(n_617),
.B1(n_595),
.B2(n_980),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1653),
.A2(n_1539),
.B(n_1526),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1640),
.A2(n_676),
.B(n_651),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1664),
.B(n_1509),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1649),
.Y(n_1712)
);

AO31x2_ASAP7_75t_L g1713 ( 
.A1(n_1646),
.A2(n_949),
.A3(n_917),
.B(n_677),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1665),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1620),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1665),
.B(n_1526),
.Y(n_1716)
);

O2A1O1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1645),
.A2(n_1588),
.B(n_1611),
.C(n_1624),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1665),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1627),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1637),
.B(n_1509),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1627),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1609),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1609),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_SL g1724 ( 
.A(n_1662),
.B(n_1534),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1595),
.A2(n_688),
.B(n_682),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1605),
.A2(n_1512),
.B(n_1539),
.Y(n_1726)
);

OA21x2_ASAP7_75t_L g1727 ( 
.A1(n_1654),
.A2(n_689),
.B(n_688),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1607),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1681),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1728),
.B(n_1603),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1678),
.A2(n_1658),
.B(n_1667),
.Y(n_1731)
);

AO21x2_ASAP7_75t_L g1732 ( 
.A1(n_1714),
.A2(n_1616),
.B(n_1605),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1722),
.B(n_1607),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1708),
.A2(n_1638),
.B1(n_1610),
.B2(n_1656),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1707),
.A2(n_1618),
.B(n_1635),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1680),
.B(n_1668),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1697),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1698),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1680),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1681),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1675),
.B(n_1622),
.Y(n_1741)
);

BUFx12f_ASAP7_75t_L g1742 ( 
.A(n_1701),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1723),
.B(n_1634),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1673),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1717),
.A2(n_1588),
.B(n_1659),
.C(n_1597),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1671),
.B(n_1644),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1678),
.A2(n_1612),
.B(n_1628),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1693),
.A2(n_1632),
.B(n_1639),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1719),
.Y(n_1749)
);

OA21x2_ASAP7_75t_L g1750 ( 
.A1(n_1718),
.A2(n_1659),
.B(n_1655),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1719),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1693),
.A2(n_1599),
.B(n_1643),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1715),
.Y(n_1753)
);

BUFx8_ASAP7_75t_L g1754 ( 
.A(n_1701),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1721),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1704),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1680),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1688),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1674),
.B(n_1590),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1693),
.A2(n_1666),
.B(n_1612),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1726),
.A2(n_1666),
.B(n_1651),
.Y(n_1761)
);

OAI21x1_ASAP7_75t_L g1762 ( 
.A1(n_1670),
.A2(n_692),
.B(n_689),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1706),
.Y(n_1763)
);

CKINVDCx11_ASAP7_75t_R g1764 ( 
.A(n_1676),
.Y(n_1764)
);

OAI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1689),
.A2(n_694),
.B(n_692),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1691),
.A2(n_1657),
.B1(n_1619),
.B2(n_1591),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1694),
.B(n_1652),
.Y(n_1767)
);

NAND2x1_ASAP7_75t_L g1768 ( 
.A(n_1716),
.B(n_1509),
.Y(n_1768)
);

OA21x2_ASAP7_75t_L g1769 ( 
.A1(n_1721),
.A2(n_696),
.B(n_694),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1715),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1702),
.Y(n_1771)
);

OA21x2_ASAP7_75t_L g1772 ( 
.A1(n_1690),
.A2(n_697),
.B(n_696),
.Y(n_1772)
);

AO21x2_ASAP7_75t_L g1773 ( 
.A1(n_1683),
.A2(n_1661),
.B(n_1652),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1695),
.Y(n_1774)
);

OAI21x1_ASAP7_75t_L g1775 ( 
.A1(n_1689),
.A2(n_698),
.B(n_697),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1725),
.A2(n_703),
.B(n_698),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1685),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1774),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1739),
.B(n_1711),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1774),
.Y(n_1780)
);

OA21x2_ASAP7_75t_L g1781 ( 
.A1(n_1731),
.A2(n_1725),
.B(n_1716),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1739),
.B(n_1757),
.Y(n_1782)
);

BUFx4f_ASAP7_75t_SL g1783 ( 
.A(n_1742),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1777),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1741),
.B(n_1712),
.Y(n_1785)
);

CKINVDCx20_ASAP7_75t_R g1786 ( 
.A(n_1764),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1729),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1744),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1739),
.B(n_1684),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1739),
.Y(n_1790)
);

AO21x2_ASAP7_75t_L g1791 ( 
.A1(n_1760),
.A2(n_1699),
.B(n_1707),
.Y(n_1791)
);

AO21x2_ASAP7_75t_L g1792 ( 
.A1(n_1737),
.A2(n_1699),
.B(n_1679),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1758),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1757),
.B(n_1684),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1757),
.B(n_1684),
.Y(n_1795)
);

OAI21x1_ASAP7_75t_L g1796 ( 
.A1(n_1747),
.A2(n_1731),
.B(n_1761),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1737),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1756),
.Y(n_1798)
);

BUFx2_ASAP7_75t_SL g1799 ( 
.A(n_1753),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1756),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1763),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1763),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1757),
.B(n_1684),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1769),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1769),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1769),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1729),
.Y(n_1807)
);

BUFx3_ASAP7_75t_L g1808 ( 
.A(n_1757),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1729),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1769),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1740),
.B(n_1713),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1757),
.B(n_1713),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1740),
.B(n_1713),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1741),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1740),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1749),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1749),
.B(n_1713),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1749),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1751),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1751),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1751),
.Y(n_1821)
);

AOI21x1_ASAP7_75t_L g1822 ( 
.A1(n_1772),
.A2(n_1716),
.B(n_1727),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1755),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1755),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1755),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1747),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1736),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1771),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1742),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1771),
.Y(n_1830)
);

CKINVDCx11_ASAP7_75t_R g1831 ( 
.A(n_1742),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1814),
.B(n_1773),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_SL g1833 ( 
.A1(n_1783),
.A2(n_1734),
.B1(n_1698),
.B2(n_1772),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1793),
.B(n_1773),
.Y(n_1834)
);

OA21x2_ASAP7_75t_L g1835 ( 
.A1(n_1796),
.A2(n_1762),
.B(n_1752),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1797),
.Y(n_1836)
);

OAI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1783),
.A2(n_1698),
.B1(n_1766),
.B2(n_1687),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1797),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1792),
.A2(n_1773),
.B1(n_1736),
.B2(n_1691),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1782),
.B(n_1771),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1786),
.A2(n_1745),
.B1(n_1766),
.B2(n_1679),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1782),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1792),
.A2(n_1736),
.B1(n_1708),
.B2(n_1687),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1792),
.A2(n_1736),
.B1(n_1687),
.B2(n_1698),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1792),
.A2(n_1748),
.B(n_1735),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1794),
.A2(n_904),
.B1(n_833),
.B2(n_814),
.C(n_715),
.Y(n_1846)
);

AOI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1815),
.A2(n_1768),
.B(n_1730),
.Y(n_1847)
);

AOI21x1_ASAP7_75t_L g1848 ( 
.A1(n_1815),
.A2(n_1768),
.B(n_1743),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1792),
.A2(n_1735),
.B1(n_1705),
.B2(n_1772),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1790),
.Y(n_1850)
);

OAI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1786),
.A2(n_1772),
.B1(n_1738),
.B2(n_1696),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1782),
.B(n_1753),
.Y(n_1852)
);

OAI31xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1788),
.A2(n_1762),
.A3(n_1622),
.B(n_1709),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1790),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1814),
.B(n_1770),
.Y(n_1855)
);

BUFx4f_ASAP7_75t_SL g1856 ( 
.A(n_1788),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1787),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1827),
.B(n_1770),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_SL g1859 ( 
.A1(n_1794),
.A2(n_1754),
.B1(n_1738),
.B2(n_1759),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1798),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1831),
.A2(n_1677),
.B1(n_1619),
.B2(n_1702),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1798),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1829),
.B(n_1746),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1836),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1857),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1834),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1836),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1842),
.B(n_1794),
.Y(n_1868)
);

NOR2x1_ASAP7_75t_SL g1869 ( 
.A(n_1847),
.B(n_1799),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1847),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1841),
.A2(n_1827),
.B1(n_1791),
.B2(n_1831),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1834),
.B(n_1799),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1857),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1857),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1838),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1838),
.B(n_1793),
.Y(n_1876)
);

BUFx3_ASAP7_75t_L g1877 ( 
.A(n_1856),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1860),
.B(n_1785),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1842),
.B(n_1795),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1860),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1850),
.B(n_1790),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1848),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1850),
.B(n_1795),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1848),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1862),
.B(n_1832),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1832),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1841),
.A2(n_1784),
.B1(n_1767),
.B2(n_1733),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1854),
.B(n_1790),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1833),
.B(n_1784),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1862),
.B(n_1785),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1854),
.B(n_1795),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1855),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1855),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1858),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1890),
.B(n_1779),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1883),
.B(n_1891),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1864),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1864),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1875),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1887),
.B(n_1853),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1887),
.B(n_1853),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1875),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1870),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1867),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1869),
.B(n_1827),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1867),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1883),
.B(n_1840),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1865),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1890),
.B(n_1779),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1880),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1883),
.B(n_1840),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1891),
.B(n_1858),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1865),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1880),
.Y(n_1914)
);

BUFx3_ASAP7_75t_L g1915 ( 
.A(n_1877),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1876),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1876),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1891),
.B(n_1852),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1877),
.B(n_1863),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1866),
.B(n_1846),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1868),
.B(n_1852),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1868),
.B(n_1803),
.Y(n_1922)
);

AND2x4_ASAP7_75t_SL g1923 ( 
.A(n_1881),
.B(n_1843),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1892),
.B(n_1846),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1869),
.B(n_1827),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1865),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1866),
.B(n_1778),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_SL g1928 ( 
.A(n_1915),
.B(n_1877),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1915),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1900),
.A2(n_1889),
.B1(n_1871),
.B2(n_1837),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1897),
.Y(n_1931)
);

AOI33xp33_ASAP7_75t_L g1932 ( 
.A1(n_1923),
.A2(n_1849),
.A3(n_1839),
.B1(n_1851),
.B2(n_709),
.B3(n_715),
.Y(n_1932)
);

AND2x4_ASAP7_75t_SL g1933 ( 
.A(n_1919),
.B(n_1907),
.Y(n_1933)
);

OAI33xp33_ASAP7_75t_L g1934 ( 
.A1(n_1901),
.A2(n_1920),
.A3(n_1924),
.B1(n_1899),
.B2(n_1898),
.B3(n_1902),
.Y(n_1934)
);

AOI33xp33_ASAP7_75t_L g1935 ( 
.A1(n_1923),
.A2(n_1896),
.A3(n_1917),
.B1(n_1916),
.B2(n_709),
.B3(n_717),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1915),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1920),
.A2(n_1845),
.B1(n_1870),
.B2(n_1844),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1923),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1907),
.B(n_1911),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1911),
.B(n_1892),
.Y(n_1940)
);

AND2x4_ASAP7_75t_SL g1941 ( 
.A(n_1896),
.B(n_1881),
.Y(n_1941)
);

INVxp67_ASAP7_75t_SL g1942 ( 
.A(n_1903),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1904),
.Y(n_1943)
);

AOI221xp5_ASAP7_75t_L g1944 ( 
.A1(n_1916),
.A2(n_1870),
.B1(n_720),
.B2(n_721),
.C(n_717),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1903),
.A2(n_1870),
.B1(n_1791),
.B2(n_1861),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1918),
.B(n_1893),
.Y(n_1946)
);

OAI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1917),
.A2(n_1859),
.B1(n_1872),
.B2(n_1870),
.C(n_1882),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1895),
.B(n_1909),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1895),
.B(n_1894),
.Y(n_1949)
);

NAND4xp25_ASAP7_75t_SL g1950 ( 
.A(n_1918),
.B(n_1872),
.C(n_1879),
.D(n_1868),
.Y(n_1950)
);

AO21x2_ASAP7_75t_L g1951 ( 
.A1(n_1898),
.A2(n_1884),
.B(n_1882),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1904),
.Y(n_1952)
);

OAI321xp33_ASAP7_75t_L g1953 ( 
.A1(n_1899),
.A2(n_1870),
.A3(n_1882),
.B1(n_1884),
.B2(n_1886),
.C(n_1885),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_R g1954 ( 
.A(n_1903),
.B(n_1724),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1906),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1906),
.Y(n_1956)
);

OA21x2_ASAP7_75t_L g1957 ( 
.A1(n_1908),
.A2(n_1884),
.B(n_1874),
.Y(n_1957)
);

INVxp67_ASAP7_75t_SL g1958 ( 
.A(n_1903),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1931),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1935),
.B(n_1912),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1957),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1939),
.B(n_1909),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1933),
.B(n_1912),
.Y(n_1963)
);

AND2x4_ASAP7_75t_SL g1964 ( 
.A(n_1929),
.B(n_1905),
.Y(n_1964)
);

AOI211x1_ASAP7_75t_L g1965 ( 
.A1(n_1947),
.A2(n_1902),
.B(n_1927),
.C(n_1914),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1936),
.B(n_1922),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1938),
.B(n_1922),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1931),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1941),
.B(n_1921),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1943),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1952),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1957),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1928),
.B(n_1929),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1955),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1957),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1929),
.B(n_1921),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1956),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1929),
.B(n_1932),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1940),
.B(n_1905),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1946),
.B(n_1905),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1942),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1934),
.A2(n_1927),
.B(n_1905),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1942),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1951),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1958),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1958),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1948),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1951),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1954),
.B(n_1925),
.Y(n_1989)
);

BUFx2_ASAP7_75t_L g1990 ( 
.A(n_1954),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1937),
.B(n_1925),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1944),
.B(n_1894),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1949),
.B(n_1910),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1937),
.B(n_1925),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1930),
.B(n_1910),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1945),
.B(n_1925),
.Y(n_1996)
);

INVxp67_ASAP7_75t_SL g1997 ( 
.A(n_1945),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1953),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1950),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1931),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1931),
.Y(n_2001)
);

AND2x2_ASAP7_75t_SL g2002 ( 
.A(n_1932),
.B(n_1870),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1997),
.A2(n_1914),
.B1(n_1881),
.B2(n_1888),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1960),
.B(n_1894),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_2002),
.B(n_1893),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1976),
.B(n_1881),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1966),
.B(n_1881),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1986),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_2002),
.B(n_1878),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_2001),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1984),
.Y(n_2011)
);

INVx4_ASAP7_75t_L g2012 ( 
.A(n_1984),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1966),
.B(n_1888),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1987),
.B(n_1878),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1981),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1976),
.B(n_1888),
.Y(n_2016)
);

INVx1_ASAP7_75t_SL g2017 ( 
.A(n_1973),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1973),
.B(n_1888),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1981),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_2002),
.B(n_1879),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1987),
.B(n_1885),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1983),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1990),
.B(n_1879),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1962),
.B(n_1886),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1962),
.B(n_1886),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1967),
.B(n_1888),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1983),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1978),
.B(n_1992),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1990),
.B(n_1995),
.Y(n_2029)
);

INVx1_ASAP7_75t_SL g2030 ( 
.A(n_1967),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1965),
.B(n_1754),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1963),
.B(n_1908),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1985),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1985),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1998),
.B(n_1908),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1959),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1999),
.B(n_1676),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1998),
.B(n_1913),
.Y(n_2038)
);

BUFx2_ASAP7_75t_L g2039 ( 
.A(n_1963),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1984),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1969),
.B(n_1913),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1969),
.B(n_1913),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1959),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1999),
.B(n_1926),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1991),
.B(n_1926),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1991),
.B(n_1926),
.Y(n_2046)
);

INVxp67_ASAP7_75t_L g2047 ( 
.A(n_1968),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1994),
.B(n_1873),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1995),
.B(n_1779),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1968),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1994),
.B(n_1873),
.Y(n_2051)
);

NOR2x1_ASAP7_75t_L g2052 ( 
.A(n_1988),
.B(n_980),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1995),
.B(n_703),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1995),
.B(n_1873),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2000),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1999),
.B(n_1874),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1989),
.B(n_1874),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1989),
.B(n_1979),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_2000),
.B(n_1982),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1970),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_1993),
.B(n_1720),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1965),
.B(n_720),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1970),
.B(n_721),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1979),
.B(n_1808),
.Y(n_2064)
);

AND2x2_ASAP7_75t_SL g2065 ( 
.A(n_1988),
.B(n_1996),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1980),
.B(n_1803),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_2039),
.Y(n_2067)
);

NOR2xp67_ASAP7_75t_L g2068 ( 
.A(n_2029),
.B(n_1993),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2040),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2030),
.B(n_2017),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2023),
.B(n_2010),
.Y(n_2071)
);

NAND3xp33_ASAP7_75t_L g2072 ( 
.A(n_2059),
.B(n_1974),
.C(n_1971),
.Y(n_2072)
);

INVxp67_ASAP7_75t_L g2073 ( 
.A(n_2058),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_2035),
.B(n_1971),
.Y(n_2074)
);

OAI32xp33_ASAP7_75t_L g2075 ( 
.A1(n_2059),
.A2(n_2031),
.A3(n_2009),
.B1(n_2062),
.B2(n_2020),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2040),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2011),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2011),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2015),
.Y(n_2079)
);

OAI32xp33_ASAP7_75t_L g2080 ( 
.A1(n_2031),
.A2(n_1996),
.A3(n_1975),
.B1(n_1972),
.B2(n_1961),
.Y(n_2080)
);

AND2x4_ASAP7_75t_L g2081 ( 
.A(n_2058),
.B(n_1964),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2019),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2022),
.Y(n_2083)
);

INVxp67_ASAP7_75t_SL g2084 ( 
.A(n_2047),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2027),
.Y(n_2085)
);

NAND3xp33_ASAP7_75t_SL g2086 ( 
.A(n_2028),
.B(n_1975),
.C(n_1961),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2033),
.Y(n_2087)
);

AND2x4_ASAP7_75t_L g2088 ( 
.A(n_2008),
.B(n_1964),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2018),
.B(n_1980),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2044),
.B(n_1974),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2034),
.Y(n_2091)
);

INVx1_ASAP7_75t_SL g2092 ( 
.A(n_2018),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2006),
.B(n_1964),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_2047),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_SL g2095 ( 
.A1(n_2065),
.A2(n_1972),
.B1(n_1975),
.B2(n_1961),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2016),
.B(n_1977),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2012),
.Y(n_2097)
);

OAI32xp33_ASAP7_75t_L g2098 ( 
.A1(n_2005),
.A2(n_1972),
.A3(n_1977),
.B1(n_1803),
.B2(n_1808),
.Y(n_2098)
);

OAI22xp33_ASAP7_75t_L g2099 ( 
.A1(n_2003),
.A2(n_1808),
.B1(n_1830),
.B2(n_1828),
.Y(n_2099)
);

INVxp67_ASAP7_75t_L g2100 ( 
.A(n_2037),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2007),
.Y(n_2101)
);

INVx2_ASAP7_75t_SL g2102 ( 
.A(n_2007),
.Y(n_2102)
);

AND2x4_ASAP7_75t_SL g2103 ( 
.A(n_2037),
.B(n_1754),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2012),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_2053),
.B(n_1754),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2012),
.Y(n_2106)
);

INVx1_ASAP7_75t_SL g2107 ( 
.A(n_2032),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_2045),
.Y(n_2108)
);

AOI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2065),
.A2(n_1672),
.B1(n_1812),
.B2(n_1789),
.Y(n_2109)
);

O2A1O1Ixp5_ASAP7_75t_L g2110 ( 
.A1(n_2036),
.A2(n_726),
.B(n_727),
.C(n_724),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2056),
.B(n_724),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2013),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2043),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2050),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2013),
.Y(n_2115)
);

AOI21xp33_ASAP7_75t_SL g2116 ( 
.A1(n_2004),
.A2(n_727),
.B(n_726),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_2038),
.B(n_738),
.Y(n_2117)
);

AOI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_2026),
.A2(n_2042),
.B1(n_2041),
.B2(n_2064),
.Y(n_2118)
);

O2A1O1Ixp33_ASAP7_75t_L g2119 ( 
.A1(n_2052),
.A2(n_771),
.B(n_777),
.C(n_738),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2055),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2056),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2045),
.B(n_2046),
.Y(n_2122)
);

AOI21xp33_ASAP7_75t_L g2123 ( 
.A1(n_2054),
.A2(n_777),
.B(n_771),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_2049),
.A2(n_2014),
.B1(n_2021),
.B2(n_2061),
.Y(n_2124)
);

AO22x1_ASAP7_75t_L g2125 ( 
.A1(n_2046),
.A2(n_1622),
.B1(n_1702),
.B2(n_828),
.Y(n_2125)
);

INVx1_ASAP7_75t_SL g2126 ( 
.A(n_2048),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2066),
.B(n_1808),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2060),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2066),
.Y(n_2129)
);

AOI32xp33_ASAP7_75t_L g2130 ( 
.A1(n_2048),
.A2(n_2051),
.A3(n_2057),
.B1(n_2063),
.B2(n_2025),
.Y(n_2130)
);

INVx5_ASAP7_75t_L g2131 ( 
.A(n_2057),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2024),
.A2(n_2051),
.B1(n_1828),
.B2(n_1830),
.Y(n_2132)
);

NOR2x1_ASAP7_75t_L g2133 ( 
.A(n_2052),
.B(n_993),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2040),
.Y(n_2134)
);

OA21x2_ASAP7_75t_L g2135 ( 
.A1(n_2062),
.A2(n_783),
.B(n_779),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2017),
.B(n_779),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2040),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_2007),
.Y(n_2138)
);

NAND4xp75_ASAP7_75t_L g2139 ( 
.A(n_2065),
.B(n_1669),
.C(n_790),
.D(n_807),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2039),
.B(n_1672),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2039),
.B(n_1672),
.Y(n_2141)
);

AO21x1_ASAP7_75t_L g2142 ( 
.A1(n_2012),
.A2(n_790),
.B(n_783),
.Y(n_2142)
);

AOI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2059),
.A2(n_1812),
.B1(n_1789),
.B2(n_807),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2039),
.B(n_1789),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2039),
.B(n_804),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2040),
.Y(n_2146)
);

OAI32xp33_ASAP7_75t_L g2147 ( 
.A1(n_2059),
.A2(n_815),
.A3(n_828),
.B1(n_814),
.B2(n_804),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2040),
.Y(n_2148)
);

NAND4xp25_ASAP7_75t_SL g2149 ( 
.A(n_2030),
.B(n_833),
.C(n_834),
.D(n_815),
.Y(n_2149)
);

BUFx2_ASAP7_75t_L g2150 ( 
.A(n_2039),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2040),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_2059),
.A2(n_1791),
.B1(n_1835),
.B2(n_1738),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2059),
.A2(n_1780),
.B1(n_1778),
.B2(n_1800),
.Y(n_2153)
);

AOI321xp33_ASAP7_75t_L g2154 ( 
.A1(n_2075),
.A2(n_1700),
.A3(n_835),
.B1(n_851),
.B2(n_858),
.C(n_854),
.Y(n_2154)
);

AOI222xp33_ASAP7_75t_L g2155 ( 
.A1(n_2086),
.A2(n_835),
.B1(n_851),
.B2(n_858),
.C1(n_854),
.C2(n_834),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2108),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2150),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2069),
.Y(n_2158)
);

NOR2x1_ASAP7_75t_L g2159 ( 
.A(n_2133),
.B(n_993),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2069),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2092),
.B(n_860),
.Y(n_2161)
);

INVx2_ASAP7_75t_SL g2162 ( 
.A(n_2131),
.Y(n_2162)
);

INVx1_ASAP7_75t_SL g2163 ( 
.A(n_2081),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_2131),
.Y(n_2164)
);

AOI211xp5_ASAP7_75t_SL g2165 ( 
.A1(n_2073),
.A2(n_864),
.B(n_868),
.C(n_860),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2143),
.A2(n_868),
.B1(n_876),
.B2(n_864),
.Y(n_2166)
);

OAI21xp33_ASAP7_75t_L g2167 ( 
.A1(n_2089),
.A2(n_1812),
.B(n_879),
.Y(n_2167)
);

AOI31xp33_ASAP7_75t_L g2168 ( 
.A1(n_2142),
.A2(n_879),
.A3(n_881),
.B(n_876),
.Y(n_2168)
);

NOR2xp67_ASAP7_75t_SL g2169 ( 
.A(n_2139),
.B(n_881),
.Y(n_2169)
);

NAND3xp33_ASAP7_75t_L g2170 ( 
.A(n_2072),
.B(n_892),
.C(n_889),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2067),
.B(n_889),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2102),
.B(n_892),
.Y(n_2172)
);

INVxp67_ASAP7_75t_L g2173 ( 
.A(n_2081),
.Y(n_2173)
);

INVxp67_ASAP7_75t_L g2174 ( 
.A(n_2122),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_2100),
.B(n_897),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2068),
.B(n_897),
.Y(n_2176)
);

AOI22xp33_ASAP7_75t_SL g2177 ( 
.A1(n_2080),
.A2(n_617),
.B1(n_595),
.B2(n_1738),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2151),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_2118),
.A2(n_1780),
.B1(n_903),
.B2(n_904),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2070),
.A2(n_903),
.B1(n_912),
.B2(n_898),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2151),
.Y(n_2181)
);

AOI22xp5_ASAP7_75t_L g2182 ( 
.A1(n_2084),
.A2(n_912),
.B1(n_920),
.B2(n_898),
.Y(n_2182)
);

NAND2xp33_ASAP7_75t_SL g2183 ( 
.A(n_2138),
.B(n_593),
.Y(n_2183)
);

INVxp67_ASAP7_75t_L g2184 ( 
.A(n_2094),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2121),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2093),
.B(n_920),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2138),
.B(n_2107),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2121),
.Y(n_2188)
);

AOI221xp5_ASAP7_75t_L g2189 ( 
.A1(n_2147),
.A2(n_942),
.B1(n_945),
.B2(n_939),
.C(n_936),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2126),
.B(n_936),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_2103),
.Y(n_2191)
);

INVxp33_ASAP7_75t_L g2192 ( 
.A(n_2105),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2153),
.A2(n_942),
.B(n_939),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2076),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2071),
.B(n_945),
.Y(n_2195)
);

O2A1O1Ixp5_ASAP7_75t_L g2196 ( 
.A1(n_2098),
.A2(n_954),
.B(n_961),
.C(n_957),
.Y(n_2196)
);

AOI211xp5_ASAP7_75t_L g2197 ( 
.A1(n_2116),
.A2(n_954),
.B(n_961),
.C(n_957),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2134),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2088),
.B(n_966),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2137),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2146),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2101),
.B(n_966),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2112),
.B(n_971),
.Y(n_2203)
);

BUFx3_ASAP7_75t_L g2204 ( 
.A(n_2088),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2115),
.B(n_971),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2140),
.B(n_2141),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2148),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_2131),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2129),
.Y(n_2209)
);

NOR4xp25_ASAP7_75t_L g2210 ( 
.A(n_2077),
.B(n_975),
.C(n_982),
.D(n_979),
.Y(n_2210)
);

AOI211xp5_ASAP7_75t_L g2211 ( 
.A1(n_2124),
.A2(n_975),
.B(n_982),
.C(n_979),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2078),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2090),
.Y(n_2213)
);

AOI22xp33_ASAP7_75t_L g2214 ( 
.A1(n_2152),
.A2(n_1791),
.B1(n_1835),
.B2(n_986),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2074),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2113),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2113),
.Y(n_2217)
);

NOR4xp25_ASAP7_75t_SL g2218 ( 
.A(n_2097),
.B(n_589),
.C(n_591),
.D(n_587),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2104),
.Y(n_2219)
);

O2A1O1Ixp5_ASAP7_75t_SL g2220 ( 
.A1(n_2106),
.A2(n_987),
.B(n_1004),
.C(n_986),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2096),
.B(n_2130),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2145),
.Y(n_2222)
);

INVxp67_ASAP7_75t_L g2223 ( 
.A(n_2136),
.Y(n_2223)
);

AND2x4_ASAP7_75t_L g2224 ( 
.A(n_2114),
.B(n_987),
.Y(n_2224)
);

OR2x2_ASAP7_75t_L g2225 ( 
.A(n_2149),
.B(n_1004),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2117),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2111),
.Y(n_2227)
);

OAI21xp33_ASAP7_75t_L g2228 ( 
.A1(n_2109),
.A2(n_1006),
.B(n_949),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2120),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2135),
.B(n_1006),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2144),
.B(n_594),
.Y(n_2231)
);

AOI221x1_ASAP7_75t_SL g2232 ( 
.A1(n_2079),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.C(n_3),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2082),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2083),
.Y(n_2234)
);

AOI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_2095),
.A2(n_599),
.B1(n_603),
.B2(n_598),
.C(n_596),
.Y(n_2235)
);

AOI221xp5_ASAP7_75t_L g2236 ( 
.A1(n_2085),
.A2(n_608),
.B1(n_609),
.B2(n_605),
.C(n_604),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2127),
.B(n_612),
.Y(n_2237)
);

NAND3xp33_ASAP7_75t_L g2238 ( 
.A(n_2110),
.B(n_686),
.C(n_672),
.Y(n_2238)
);

OAI221xp5_ASAP7_75t_L g2239 ( 
.A1(n_2119),
.A2(n_2091),
.B1(n_2087),
.B2(n_2128),
.C(n_2135),
.Y(n_2239)
);

OAI21xp33_ASAP7_75t_L g2240 ( 
.A1(n_2123),
.A2(n_618),
.B(n_614),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2132),
.B(n_620),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2125),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_2099),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2131),
.Y(n_2244)
);

AOI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2086),
.A2(n_661),
.B1(n_680),
.B2(n_640),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2089),
.B(n_621),
.Y(n_2246)
);

A2O1A1Ixp33_ASAP7_75t_L g2247 ( 
.A1(n_2143),
.A2(n_631),
.B(n_632),
.C(n_623),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2108),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_SL g2249 ( 
.A(n_2150),
.B(n_1512),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2108),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2108),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2150),
.B(n_636),
.Y(n_2252)
);

OAI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2143),
.A2(n_1801),
.B1(n_1802),
.B2(n_1800),
.Y(n_2253)
);

INVxp67_ASAP7_75t_L g2254 ( 
.A(n_2150),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2108),
.Y(n_2255)
);

NOR4xp25_ASAP7_75t_L g2256 ( 
.A(n_2086),
.B(n_6),
.C(n_2),
.D(n_4),
.Y(n_2256)
);

OAI221xp5_ASAP7_75t_L g2257 ( 
.A1(n_2143),
.A2(n_643),
.B1(n_644),
.B2(n_641),
.C(n_637),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2108),
.Y(n_2258)
);

AOI221xp5_ASAP7_75t_L g2259 ( 
.A1(n_2075),
.A2(n_656),
.B1(n_660),
.B2(n_654),
.C(n_653),
.Y(n_2259)
);

AOI322xp5_ASAP7_75t_L g2260 ( 
.A1(n_2086),
.A2(n_669),
.A3(n_665),
.B1(n_670),
.B2(n_673),
.C1(n_667),
.C2(n_662),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2131),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2150),
.B(n_681),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2108),
.Y(n_2263)
);

OR2x2_ASAP7_75t_L g2264 ( 
.A(n_2150),
.B(n_6),
.Y(n_2264)
);

NAND2x1_ASAP7_75t_L g2265 ( 
.A(n_2081),
.B(n_1835),
.Y(n_2265)
);

OAI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_2143),
.A2(n_1802),
.B1(n_1801),
.B2(n_1826),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2150),
.B(n_683),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2108),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2108),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2150),
.B(n_684),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2108),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2150),
.B(n_685),
.Y(n_2272)
);

AOI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2086),
.A2(n_740),
.B1(n_753),
.B2(n_713),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2089),
.B(n_687),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_2100),
.B(n_691),
.Y(n_2275)
);

HB1xp67_ASAP7_75t_L g2276 ( 
.A(n_2131),
.Y(n_2276)
);

XOR2x2_ASAP7_75t_L g2277 ( 
.A(n_2139),
.B(n_7),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2089),
.B(n_693),
.Y(n_2278)
);

INVx1_ASAP7_75t_SL g2279 ( 
.A(n_2150),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2150),
.B(n_705),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_2150),
.B(n_7),
.Y(n_2281)
);

NOR2x1_ASAP7_75t_SL g2282 ( 
.A(n_2131),
.B(n_672),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2108),
.Y(n_2283)
);

INVx1_ASAP7_75t_SL g2284 ( 
.A(n_2150),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_SL g2285 ( 
.A(n_2150),
.B(n_710),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_2081),
.B(n_1826),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2108),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_2100),
.B(n_708),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2150),
.B(n_711),
.Y(n_2289)
);

AOI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_2086),
.A2(n_1791),
.B1(n_1835),
.B2(n_1796),
.Y(n_2290)
);

OAI22xp33_ASAP7_75t_L g2291 ( 
.A1(n_2143),
.A2(n_1805),
.B1(n_1806),
.B2(n_1804),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2150),
.B(n_718),
.Y(n_2292)
);

AOI221xp5_ASAP7_75t_L g2293 ( 
.A1(n_2075),
.A2(n_728),
.B1(n_734),
.B2(n_732),
.C(n_725),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_2150),
.B(n_8),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2089),
.B(n_735),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2131),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2108),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2108),
.Y(n_2298)
);

AOI21xp33_ASAP7_75t_L g2299 ( 
.A1(n_2070),
.A2(n_743),
.B(n_737),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2108),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2089),
.B(n_746),
.Y(n_2301)
);

O2A1O1Ixp33_ASAP7_75t_L g2302 ( 
.A1(n_2147),
.A2(n_1826),
.B(n_1677),
.C(n_12),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2089),
.B(n_747),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2164),
.Y(n_2304)
);

OR2x2_ASAP7_75t_L g2305 ( 
.A(n_2279),
.B(n_10),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2208),
.Y(n_2306)
);

INVx2_ASAP7_75t_SL g2307 ( 
.A(n_2204),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2163),
.B(n_749),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2276),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2264),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2281),
.Y(n_2311)
);

NAND3xp33_ASAP7_75t_SL g2312 ( 
.A(n_2256),
.B(n_751),
.C(n_750),
.Y(n_2312)
);

AOI21xp33_ASAP7_75t_L g2313 ( 
.A1(n_2192),
.A2(n_757),
.B(n_756),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2294),
.Y(n_2314)
);

INVx1_ASAP7_75t_SL g2315 ( 
.A(n_2284),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_2173),
.B(n_759),
.Y(n_2316)
);

AND2x4_ASAP7_75t_L g2317 ( 
.A(n_2162),
.B(n_11),
.Y(n_2317)
);

OAI21xp33_ASAP7_75t_SL g2318 ( 
.A1(n_2245),
.A2(n_1796),
.B(n_1826),
.Y(n_2318)
);

AOI321xp33_ASAP7_75t_L g2319 ( 
.A1(n_2221),
.A2(n_1703),
.A3(n_14),
.B1(n_16),
.B2(n_11),
.C(n_13),
.Y(n_2319)
);

OAI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2254),
.A2(n_763),
.B1(n_765),
.B2(n_761),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_SL g2321 ( 
.A1(n_2243),
.A2(n_2157),
.B1(n_2285),
.B2(n_2191),
.Y(n_2321)
);

OAI22xp5_ASAP7_75t_SL g2322 ( 
.A1(n_2177),
.A2(n_770),
.B1(n_773),
.B2(n_766),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2187),
.Y(n_2323)
);

OA21x2_ASAP7_75t_L g2324 ( 
.A1(n_2245),
.A2(n_778),
.B(n_776),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2158),
.Y(n_2325)
);

NAND4xp25_ASAP7_75t_SL g2326 ( 
.A(n_2273),
.B(n_1805),
.C(n_1806),
.D(n_1804),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2160),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_2184),
.B(n_780),
.Y(n_2328)
);

BUFx2_ASAP7_75t_SL g2329 ( 
.A(n_2244),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2206),
.B(n_785),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2174),
.B(n_786),
.Y(n_2331)
);

INVx3_ASAP7_75t_L g2332 ( 
.A(n_2261),
.Y(n_2332)
);

OAI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2273),
.A2(n_789),
.B1(n_792),
.B2(n_787),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2178),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2181),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_SL g2336 ( 
.A(n_2222),
.B(n_793),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2156),
.B(n_795),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2296),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2248),
.Y(n_2339)
);

AOI21xp33_ASAP7_75t_SL g2340 ( 
.A1(n_2168),
.A2(n_13),
.B(n_14),
.Y(n_2340)
);

OAI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2243),
.A2(n_1811),
.B1(n_1810),
.B2(n_799),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2250),
.Y(n_2342)
);

OAI22xp5_ASAP7_75t_L g2343 ( 
.A1(n_2251),
.A2(n_802),
.B1(n_805),
.B2(n_797),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2282),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2255),
.B(n_806),
.Y(n_2345)
);

INVxp67_ASAP7_75t_SL g2346 ( 
.A(n_2159),
.Y(n_2346)
);

OAI22xp33_ASAP7_75t_SL g2347 ( 
.A1(n_2249),
.A2(n_811),
.B1(n_813),
.B2(n_808),
.Y(n_2347)
);

AOI221xp5_ASAP7_75t_L g2348 ( 
.A1(n_2210),
.A2(n_816),
.B1(n_821),
.B2(n_819),
.C(n_818),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2258),
.B(n_822),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2263),
.B(n_823),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_2223),
.B(n_824),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2268),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2269),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2271),
.B(n_826),
.Y(n_2354)
);

AO22x1_ASAP7_75t_L g2355 ( 
.A1(n_2283),
.A2(n_830),
.B1(n_831),
.B2(n_827),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2287),
.B(n_832),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2297),
.Y(n_2357)
);

OR2x2_ASAP7_75t_L g2358 ( 
.A(n_2298),
.B(n_15),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2300),
.B(n_836),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2185),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2209),
.B(n_838),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2226),
.B(n_839),
.Y(n_2362)
);

A2O1A1Ixp33_ASAP7_75t_L g2363 ( 
.A1(n_2232),
.A2(n_843),
.B(n_845),
.C(n_840),
.Y(n_2363)
);

OAI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_2260),
.A2(n_880),
.B(n_862),
.Y(n_2364)
);

AO22x1_ASAP7_75t_L g2365 ( 
.A1(n_2215),
.A2(n_848),
.B1(n_850),
.B2(n_847),
.Y(n_2365)
);

NAND3xp33_ASAP7_75t_SL g2366 ( 
.A(n_2154),
.B(n_855),
.C(n_852),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_2188),
.Y(n_2367)
);

OAI322xp33_ASAP7_75t_L g2368 ( 
.A1(n_2194),
.A2(n_856),
.A3(n_869),
.B1(n_859),
.B2(n_871),
.C1(n_870),
.C2(n_863),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2198),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2242),
.B(n_686),
.Y(n_2370)
);

AOI211xp5_ASAP7_75t_L g2371 ( 
.A1(n_2259),
.A2(n_915),
.B(n_937),
.C(n_894),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2200),
.Y(n_2372)
);

INVxp67_ASAP7_75t_SL g2373 ( 
.A(n_2176),
.Y(n_2373)
);

O2A1O1Ixp33_ASAP7_75t_L g2374 ( 
.A1(n_2155),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2213),
.A2(n_878),
.B1(n_886),
.B2(n_873),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2201),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2246),
.B(n_887),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2186),
.Y(n_2378)
);

AOI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_2207),
.A2(n_895),
.B1(n_899),
.B2(n_891),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2219),
.Y(n_2380)
);

XNOR2xp5_ASAP7_75t_L g2381 ( 
.A(n_2277),
.B(n_18),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2274),
.B(n_2278),
.Y(n_2382)
);

AOI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_2167),
.A2(n_902),
.B1(n_905),
.B2(n_900),
.Y(n_2383)
);

OAI21xp33_ASAP7_75t_L g2384 ( 
.A1(n_2228),
.A2(n_908),
.B(n_907),
.Y(n_2384)
);

AOI322xp5_ASAP7_75t_L g2385 ( 
.A1(n_2293),
.A2(n_929),
.A3(n_924),
.B1(n_930),
.B2(n_933),
.C1(n_926),
.C2(n_923),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2225),
.Y(n_2386)
);

OAI21xp33_ASAP7_75t_L g2387 ( 
.A1(n_2227),
.A2(n_938),
.B(n_935),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2295),
.B(n_940),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2301),
.B(n_941),
.Y(n_2389)
);

AOI22xp5_ASAP7_75t_L g2390 ( 
.A1(n_2183),
.A2(n_2212),
.B1(n_2179),
.B2(n_2303),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2231),
.B(n_943),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2237),
.B(n_947),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_2216),
.Y(n_2393)
);

OAI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2166),
.A2(n_948),
.B1(n_955),
.B2(n_952),
.Y(n_2394)
);

OAI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2166),
.A2(n_958),
.B1(n_960),
.B2(n_959),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2202),
.B(n_962),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2199),
.Y(n_2397)
);

OR2x2_ASAP7_75t_L g2398 ( 
.A(n_2252),
.B(n_23),
.Y(n_2398)
);

OAI22xp5_ASAP7_75t_L g2399 ( 
.A1(n_2257),
.A2(n_2247),
.B1(n_2235),
.B2(n_2218),
.Y(n_2399)
);

INVxp67_ASAP7_75t_L g2400 ( 
.A(n_2169),
.Y(n_2400)
);

OR2x2_ASAP7_75t_L g2401 ( 
.A(n_2262),
.B(n_23),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2165),
.B(n_965),
.Y(n_2402)
);

XOR2x2_ASAP7_75t_L g2403 ( 
.A(n_2238),
.B(n_24),
.Y(n_2403)
);

NAND2x1_ASAP7_75t_L g2404 ( 
.A(n_2217),
.B(n_2229),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2253),
.A2(n_2288),
.B1(n_2275),
.B2(n_2266),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2175),
.B(n_2203),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2190),
.Y(n_2407)
);

OAI22xp33_ASAP7_75t_L g2408 ( 
.A1(n_2239),
.A2(n_1811),
.B1(n_1810),
.B2(n_968),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2161),
.Y(n_2409)
);

AOI31xp33_ASAP7_75t_L g2410 ( 
.A1(n_2211),
.A2(n_969),
.A3(n_970),
.B(n_967),
.Y(n_2410)
);

OA21x2_ASAP7_75t_L g2411 ( 
.A1(n_2196),
.A2(n_976),
.B(n_972),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2265),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2267),
.B(n_24),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2270),
.B(n_25),
.Y(n_2414)
);

NOR2x1_ASAP7_75t_L g2415 ( 
.A(n_2170),
.B(n_686),
.Y(n_2415)
);

O2A1O1Ixp33_ASAP7_75t_L g2416 ( 
.A1(n_2233),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_2416)
);

OAI32xp33_ASAP7_75t_L g2417 ( 
.A1(n_2234),
.A2(n_985),
.A3(n_988),
.B1(n_984),
.B2(n_981),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2195),
.B(n_2197),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2272),
.B(n_26),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2224),
.Y(n_2420)
);

OAI321xp33_ASAP7_75t_L g2421 ( 
.A1(n_2290),
.A2(n_874),
.A3(n_744),
.B1(n_888),
.B2(n_817),
.C(n_686),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2214),
.A2(n_989),
.B1(n_991),
.B2(n_990),
.Y(n_2422)
);

OAI211xp5_ASAP7_75t_SL g2423 ( 
.A1(n_2321),
.A2(n_2236),
.B(n_2289),
.C(n_2280),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2307),
.B(n_2292),
.Y(n_2424)
);

AOI22xp33_ASAP7_75t_SL g2425 ( 
.A1(n_2315),
.A2(n_2171),
.B1(n_2241),
.B2(n_2180),
.Y(n_2425)
);

O2A1O1Ixp33_ASAP7_75t_SL g2426 ( 
.A1(n_2404),
.A2(n_2230),
.B(n_2299),
.C(n_2172),
.Y(n_2426)
);

OR2x2_ASAP7_75t_L g2427 ( 
.A(n_2305),
.B(n_2205),
.Y(n_2427)
);

OAI21xp33_ASAP7_75t_L g2428 ( 
.A1(n_2323),
.A2(n_2286),
.B(n_2302),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2332),
.Y(n_2429)
);

AOI211xp5_ASAP7_75t_SL g2430 ( 
.A1(n_2347),
.A2(n_2291),
.B(n_2240),
.C(n_2193),
.Y(n_2430)
);

O2A1O1Ixp33_ASAP7_75t_L g2431 ( 
.A1(n_2312),
.A2(n_2240),
.B(n_2189),
.C(n_2224),
.Y(n_2431)
);

NAND4xp25_ASAP7_75t_L g2432 ( 
.A(n_2319),
.B(n_2182),
.C(n_2220),
.D(n_32),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2332),
.B(n_2182),
.Y(n_2433)
);

NOR3xp33_ASAP7_75t_L g2434 ( 
.A(n_2399),
.B(n_997),
.C(n_995),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2304),
.B(n_2306),
.Y(n_2435)
);

A2O1A1Ixp33_ASAP7_75t_L g2436 ( 
.A1(n_2416),
.A2(n_999),
.B(n_1000),
.C(n_998),
.Y(n_2436)
);

OAI22xp5_ASAP7_75t_L g2437 ( 
.A1(n_2400),
.A2(n_1009),
.B1(n_1007),
.B2(n_1005),
.Y(n_2437)
);

AOI221xp5_ASAP7_75t_L g2438 ( 
.A1(n_2341),
.A2(n_1012),
.B1(n_1010),
.B2(n_1013),
.C(n_817),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2309),
.B(n_28),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2317),
.Y(n_2440)
);

NOR2xp67_ASAP7_75t_L g2441 ( 
.A(n_2367),
.B(n_2393),
.Y(n_2441)
);

AOI211x1_ASAP7_75t_L g2442 ( 
.A1(n_2355),
.A2(n_1822),
.B(n_33),
.C(n_29),
.Y(n_2442)
);

A2O1A1Ixp33_ASAP7_75t_L g2443 ( 
.A1(n_2374),
.A2(n_744),
.B(n_817),
.C(n_686),
.Y(n_2443)
);

NAND3xp33_ASAP7_75t_SL g2444 ( 
.A(n_2336),
.B(n_34),
.C(n_33),
.Y(n_2444)
);

AOI21xp33_ASAP7_75t_L g2445 ( 
.A1(n_2310),
.A2(n_817),
.B(n_744),
.Y(n_2445)
);

AOI222xp33_ASAP7_75t_L g2446 ( 
.A1(n_2322),
.A2(n_888),
.B1(n_817),
.B2(n_944),
.C1(n_874),
.C2(n_744),
.Y(n_2446)
);

OAI221xp5_ASAP7_75t_L g2447 ( 
.A1(n_2338),
.A2(n_2342),
.B1(n_2353),
.B2(n_2352),
.C(n_2339),
.Y(n_2447)
);

OAI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_2357),
.A2(n_2314),
.B(n_2311),
.Y(n_2448)
);

AOI322xp5_ASAP7_75t_L g2449 ( 
.A1(n_2366),
.A2(n_1817),
.A3(n_1813),
.B1(n_1816),
.B2(n_1815),
.C1(n_1820),
.C2(n_944),
.Y(n_2449)
);

NAND3xp33_ASAP7_75t_L g2450 ( 
.A(n_2380),
.B(n_817),
.C(n_744),
.Y(n_2450)
);

O2A1O1Ixp33_ASAP7_75t_L g2451 ( 
.A1(n_2363),
.A2(n_35),
.B(n_32),
.C(n_34),
.Y(n_2451)
);

INVx3_ASAP7_75t_L g2452 ( 
.A(n_2317),
.Y(n_2452)
);

AND4x1_ASAP7_75t_L g2453 ( 
.A(n_2371),
.B(n_38),
.C(n_36),
.D(n_37),
.Y(n_2453)
);

OAI221xp5_ASAP7_75t_L g2454 ( 
.A1(n_2390),
.A2(n_2329),
.B1(n_2405),
.B2(n_2346),
.C(n_2386),
.Y(n_2454)
);

OAI21xp33_ASAP7_75t_SL g2455 ( 
.A1(n_2412),
.A2(n_1824),
.B(n_1823),
.Y(n_2455)
);

NAND4xp25_ASAP7_75t_L g2456 ( 
.A(n_2418),
.B(n_40),
.C(n_36),
.D(n_37),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2382),
.B(n_41),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2358),
.Y(n_2458)
);

NOR3xp33_ASAP7_75t_SL g2459 ( 
.A(n_2408),
.B(n_41),
.C(n_43),
.Y(n_2459)
);

O2A1O1Ixp33_ASAP7_75t_L g2460 ( 
.A1(n_2340),
.A2(n_46),
.B(n_43),
.C(n_44),
.Y(n_2460)
);

NAND4xp25_ASAP7_75t_L g2461 ( 
.A(n_2406),
.B(n_49),
.C(n_47),
.D(n_48),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2420),
.Y(n_2462)
);

A2O1A1Ixp33_ASAP7_75t_L g2463 ( 
.A1(n_2328),
.A2(n_888),
.B(n_944),
.C(n_874),
.Y(n_2463)
);

AOI211x1_ASAP7_75t_SL g2464 ( 
.A1(n_2370),
.A2(n_888),
.B(n_944),
.C(n_874),
.Y(n_2464)
);

OAI311xp33_ASAP7_75t_L g2465 ( 
.A1(n_2369),
.A2(n_49),
.A3(n_47),
.B1(n_48),
.C1(n_50),
.Y(n_2465)
);

NOR3xp33_ASAP7_75t_L g2466 ( 
.A(n_2365),
.B(n_1682),
.C(n_1776),
.Y(n_2466)
);

NOR3xp33_ASAP7_75t_L g2467 ( 
.A(n_2373),
.B(n_1776),
.C(n_1686),
.Y(n_2467)
);

OAI321xp33_ASAP7_75t_L g2468 ( 
.A1(n_2372),
.A2(n_950),
.A3(n_888),
.B1(n_1001),
.B2(n_944),
.C(n_874),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2381),
.B(n_50),
.Y(n_2469)
);

OAI33xp33_ASAP7_75t_L g2470 ( 
.A1(n_2325),
.A2(n_54),
.A3(n_59),
.B1(n_51),
.B2(n_53),
.B3(n_55),
.Y(n_2470)
);

AOI21xp5_ASAP7_75t_L g2471 ( 
.A1(n_2402),
.A2(n_888),
.B(n_874),
.Y(n_2471)
);

OAI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_2378),
.A2(n_1811),
.B1(n_1823),
.B2(n_1821),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_L g2473 ( 
.A(n_2407),
.B(n_51),
.Y(n_2473)
);

OAI21xp5_ASAP7_75t_SL g2474 ( 
.A1(n_2376),
.A2(n_2409),
.B(n_2316),
.Y(n_2474)
);

NAND4xp75_ASAP7_75t_L g2475 ( 
.A(n_2415),
.B(n_62),
.C(n_60),
.D(n_61),
.Y(n_2475)
);

AOI21xp5_ASAP7_75t_L g2476 ( 
.A1(n_2377),
.A2(n_950),
.B(n_944),
.Y(n_2476)
);

AOI221xp5_ASAP7_75t_L g2477 ( 
.A1(n_2327),
.A2(n_1001),
.B1(n_950),
.B2(n_64),
.C(n_62),
.Y(n_2477)
);

AOI221xp5_ASAP7_75t_L g2478 ( 
.A1(n_2334),
.A2(n_1001),
.B1(n_950),
.B2(n_66),
.C(n_63),
.Y(n_2478)
);

AOI211x1_ASAP7_75t_L g2479 ( 
.A1(n_2417),
.A2(n_1822),
.B(n_66),
.C(n_63),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2344),
.B(n_950),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2330),
.Y(n_2481)
);

AOI21x1_ASAP7_75t_L g2482 ( 
.A1(n_2360),
.A2(n_65),
.B(n_67),
.Y(n_2482)
);

AOI211xp5_ASAP7_75t_SL g2483 ( 
.A1(n_2421),
.A2(n_70),
.B(n_67),
.C(n_69),
.Y(n_2483)
);

AOI221xp5_ASAP7_75t_L g2484 ( 
.A1(n_2335),
.A2(n_1001),
.B1(n_950),
.B2(n_73),
.C(n_69),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2398),
.Y(n_2485)
);

NOR2xp67_ASAP7_75t_L g2486 ( 
.A(n_2326),
.B(n_71),
.Y(n_2486)
);

OAI21xp33_ASAP7_75t_L g2487 ( 
.A1(n_2397),
.A2(n_1817),
.B(n_1813),
.Y(n_2487)
);

AOI322xp5_ASAP7_75t_L g2488 ( 
.A1(n_2415),
.A2(n_1813),
.A3(n_1817),
.B1(n_1816),
.B2(n_1820),
.C1(n_1001),
.C2(n_1821),
.Y(n_2488)
);

AOI211xp5_ASAP7_75t_L g2489 ( 
.A1(n_2308),
.A2(n_1001),
.B(n_77),
.C(n_73),
.Y(n_2489)
);

OAI221xp5_ASAP7_75t_L g2490 ( 
.A1(n_2387),
.A2(n_1677),
.B1(n_78),
.B2(n_76),
.C(n_77),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2401),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2388),
.B(n_79),
.Y(n_2492)
);

AOI21xp33_ASAP7_75t_SL g2493 ( 
.A1(n_2411),
.A2(n_79),
.B(n_80),
.Y(n_2493)
);

NOR2x1_ASAP7_75t_L g2494 ( 
.A(n_2411),
.B(n_80),
.Y(n_2494)
);

OAI21xp5_ASAP7_75t_L g2495 ( 
.A1(n_2403),
.A2(n_1775),
.B(n_1765),
.Y(n_2495)
);

AOI211xp5_ASAP7_75t_SL g2496 ( 
.A1(n_2410),
.A2(n_87),
.B(n_82),
.C(n_86),
.Y(n_2496)
);

AOI211xp5_ASAP7_75t_L g2497 ( 
.A1(n_2422),
.A2(n_90),
.B(n_88),
.C(n_89),
.Y(n_2497)
);

AOI22xp5_ASAP7_75t_SL g2498 ( 
.A1(n_2324),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_2498)
);

O2A1O1Ixp33_ASAP7_75t_SL g2499 ( 
.A1(n_2337),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_2499)
);

OAI221xp5_ASAP7_75t_L g2500 ( 
.A1(n_2375),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.C(n_97),
.Y(n_2500)
);

NOR3xp33_ASAP7_75t_L g2501 ( 
.A(n_2345),
.B(n_1686),
.C(n_1765),
.Y(n_2501)
);

NOR3xp33_ASAP7_75t_L g2502 ( 
.A(n_2354),
.B(n_2356),
.C(n_2368),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_2348),
.B(n_1539),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2396),
.B(n_95),
.Y(n_2504)
);

AOI221xp5_ASAP7_75t_L g2505 ( 
.A1(n_2333),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.C(n_100),
.Y(n_2505)
);

AOI22xp5_ASAP7_75t_L g2506 ( 
.A1(n_2362),
.A2(n_1825),
.B1(n_1824),
.B2(n_1787),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2413),
.B(n_98),
.Y(n_2507)
);

AOI22xp33_ASAP7_75t_SL g2508 ( 
.A1(n_2331),
.A2(n_1750),
.B1(n_1781),
.B2(n_1820),
.Y(n_2508)
);

NAND4xp75_ASAP7_75t_L g2509 ( 
.A(n_2324),
.B(n_2350),
.C(n_2359),
.D(n_2349),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2389),
.A2(n_1775),
.B(n_1727),
.Y(n_2510)
);

XNOR2xp5_ASAP7_75t_L g2511 ( 
.A(n_2383),
.B(n_2414),
.Y(n_2511)
);

AOI221xp5_ASAP7_75t_L g2512 ( 
.A1(n_2343),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.C(n_103),
.Y(n_2512)
);

NAND3xp33_ASAP7_75t_L g2513 ( 
.A(n_2385),
.B(n_101),
.C(n_104),
.Y(n_2513)
);

OAI211xp5_ASAP7_75t_L g2514 ( 
.A1(n_2379),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_2514)
);

AOI22xp33_ASAP7_75t_SL g2515 ( 
.A1(n_2361),
.A2(n_1750),
.B1(n_1781),
.B2(n_1825),
.Y(n_2515)
);

INVx1_ASAP7_75t_SL g2516 ( 
.A(n_2419),
.Y(n_2516)
);

A2O1A1Ixp33_ASAP7_75t_L g2517 ( 
.A1(n_2351),
.A2(n_111),
.B(n_108),
.C(n_109),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2391),
.Y(n_2518)
);

OAI21xp5_ASAP7_75t_L g2519 ( 
.A1(n_2392),
.A2(n_1710),
.B(n_1692),
.Y(n_2519)
);

A2O1A1Ixp33_ASAP7_75t_L g2520 ( 
.A1(n_2384),
.A2(n_113),
.B(n_109),
.C(n_112),
.Y(n_2520)
);

AOI21xp5_ASAP7_75t_L g2521 ( 
.A1(n_2313),
.A2(n_1727),
.B(n_113),
.Y(n_2521)
);

NOR3xp33_ASAP7_75t_L g2522 ( 
.A(n_2320),
.B(n_114),
.C(n_115),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2394),
.B(n_115),
.Y(n_2523)
);

AOI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_2318),
.A2(n_2395),
.B1(n_2364),
.B2(n_1819),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2332),
.Y(n_2525)
);

NAND3xp33_ASAP7_75t_L g2526 ( 
.A(n_2319),
.B(n_116),
.C(n_117),
.Y(n_2526)
);

AOI311xp33_ASAP7_75t_L g2527 ( 
.A1(n_2323),
.A2(n_119),
.A3(n_117),
.B(n_118),
.C(n_120),
.Y(n_2527)
);

OAI21xp5_ASAP7_75t_L g2528 ( 
.A1(n_2321),
.A2(n_1710),
.B(n_119),
.Y(n_2528)
);

AOI221xp5_ASAP7_75t_L g2529 ( 
.A1(n_2341),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.C(n_123),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2332),
.Y(n_2530)
);

A2O1A1Ixp33_ASAP7_75t_L g2531 ( 
.A1(n_2319),
.A2(n_125),
.B(n_121),
.C(n_124),
.Y(n_2531)
);

OAI211xp5_ASAP7_75t_SL g2532 ( 
.A1(n_2321),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_2532)
);

OAI22xp33_ASAP7_75t_SL g2533 ( 
.A1(n_2404),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_2533)
);

OAI22xp5_ASAP7_75t_L g2534 ( 
.A1(n_2315),
.A2(n_1819),
.B1(n_1787),
.B2(n_1809),
.Y(n_2534)
);

OAI211xp5_ASAP7_75t_L g2535 ( 
.A1(n_2319),
.A2(n_131),
.B(n_128),
.C(n_130),
.Y(n_2535)
);

AOI21xp5_ASAP7_75t_L g2536 ( 
.A1(n_2312),
.A2(n_130),
.B(n_131),
.Y(n_2536)
);

AOI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_2312),
.A2(n_132),
.B(n_133),
.Y(n_2537)
);

AOI221xp5_ASAP7_75t_L g2538 ( 
.A1(n_2341),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_2538)
);

AOI21xp33_ASAP7_75t_L g2539 ( 
.A1(n_2315),
.A2(n_134),
.B(n_136),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2307),
.B(n_138),
.Y(n_2540)
);

AOI221xp5_ASAP7_75t_L g2541 ( 
.A1(n_2341),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.C(n_144),
.Y(n_2541)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2542 ( 
.A1(n_2319),
.A2(n_146),
.B(n_141),
.C(n_145),
.D(n_147),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2307),
.B(n_146),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2315),
.B(n_147),
.Y(n_2544)
);

O2A1O1Ixp5_ASAP7_75t_L g2545 ( 
.A1(n_2404),
.A2(n_1822),
.B(n_1819),
.C(n_1787),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2332),
.Y(n_2546)
);

AND4x1_ASAP7_75t_L g2547 ( 
.A(n_2336),
.B(n_151),
.C(n_149),
.D(n_150),
.Y(n_2547)
);

A2O1A1Ixp33_ASAP7_75t_L g2548 ( 
.A1(n_2319),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2307),
.B(n_154),
.Y(n_2549)
);

OAI211xp5_ASAP7_75t_L g2550 ( 
.A1(n_2319),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_2550)
);

OAI221xp5_ASAP7_75t_L g2551 ( 
.A1(n_2321),
.A2(n_158),
.B1(n_155),
.B2(n_157),
.C(n_159),
.Y(n_2551)
);

OAI221xp5_ASAP7_75t_SL g2552 ( 
.A1(n_2315),
.A2(n_162),
.B1(n_158),
.B2(n_159),
.C(n_163),
.Y(n_2552)
);

NOR3xp33_ASAP7_75t_SL g2553 ( 
.A(n_2341),
.B(n_162),
.C(n_164),
.Y(n_2553)
);

OAI21xp33_ASAP7_75t_L g2554 ( 
.A1(n_2321),
.A2(n_1819),
.B(n_1809),
.Y(n_2554)
);

AOI221xp5_ASAP7_75t_L g2555 ( 
.A1(n_2341),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_167),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2315),
.A2(n_1807),
.B1(n_1818),
.B2(n_1809),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2307),
.B(n_165),
.Y(n_2557)
);

OAI21xp5_ASAP7_75t_SL g2558 ( 
.A1(n_2321),
.A2(n_166),
.B(n_168),
.Y(n_2558)
);

OAI21xp5_ASAP7_75t_L g2559 ( 
.A1(n_2321),
.A2(n_168),
.B(n_169),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2307),
.B(n_169),
.Y(n_2560)
);

AOI31xp33_ASAP7_75t_L g2561 ( 
.A1(n_2315),
.A2(n_174),
.A3(n_170),
.B(n_171),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2307),
.B(n_170),
.Y(n_2562)
);

OAI21xp5_ASAP7_75t_SL g2563 ( 
.A1(n_2321),
.A2(n_171),
.B(n_175),
.Y(n_2563)
);

OAI221xp5_ASAP7_75t_SL g2564 ( 
.A1(n_2315),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.C(n_179),
.Y(n_2564)
);

INVxp67_ASAP7_75t_L g2565 ( 
.A(n_2329),
.Y(n_2565)
);

OAI211xp5_ASAP7_75t_L g2566 ( 
.A1(n_2319),
.A2(n_180),
.B(n_176),
.C(n_179),
.Y(n_2566)
);

O2A1O1Ixp5_ASAP7_75t_L g2567 ( 
.A1(n_2404),
.A2(n_1818),
.B(n_1807),
.C(n_183),
.Y(n_2567)
);

AOI32xp33_ASAP7_75t_L g2568 ( 
.A1(n_2315),
.A2(n_183),
.A3(n_181),
.B1(n_182),
.B2(n_184),
.Y(n_2568)
);

NOR2xp67_ASAP7_75t_L g2569 ( 
.A(n_2307),
.B(n_181),
.Y(n_2569)
);

OAI21xp33_ASAP7_75t_SL g2570 ( 
.A1(n_2315),
.A2(n_1818),
.B(n_1807),
.Y(n_2570)
);

OAI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2315),
.A2(n_1781),
.B1(n_1750),
.B2(n_187),
.Y(n_2571)
);

OAI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_2565),
.A2(n_2542),
.B(n_2526),
.Y(n_2572)
);

OAI211xp5_ASAP7_75t_L g2573 ( 
.A1(n_2558),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2452),
.Y(n_2574)
);

INVxp67_ASAP7_75t_L g2575 ( 
.A(n_2452),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2569),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2440),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2441),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2429),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2546),
.Y(n_2580)
);

OAI221xp5_ASAP7_75t_L g2581 ( 
.A1(n_2563),
.A2(n_191),
.B1(n_188),
.B2(n_189),
.C(n_192),
.Y(n_2581)
);

AOI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_2535),
.A2(n_1781),
.B1(n_1750),
.B2(n_1732),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2525),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2530),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2457),
.Y(n_2585)
);

AOI222xp33_ASAP7_75t_L g2586 ( 
.A1(n_2428),
.A2(n_193),
.B1(n_195),
.B2(n_188),
.C1(n_191),
.C2(n_194),
.Y(n_2586)
);

NOR2x1_ASAP7_75t_L g2587 ( 
.A(n_2561),
.B(n_193),
.Y(n_2587)
);

OAI31xp33_ASAP7_75t_L g2588 ( 
.A1(n_2550),
.A2(n_196),
.A3(n_194),
.B(n_195),
.Y(n_2588)
);

OAI221xp5_ASAP7_75t_L g2589 ( 
.A1(n_2559),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_2589)
);

AOI221xp5_ASAP7_75t_L g2590 ( 
.A1(n_2454),
.A2(n_200),
.B1(n_197),
.B2(n_199),
.C(n_201),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2482),
.Y(n_2591)
);

OAI311xp33_ASAP7_75t_L g2592 ( 
.A1(n_2448),
.A2(n_203),
.A3(n_201),
.B1(n_202),
.C1(n_204),
.Y(n_2592)
);

AOI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_2566),
.A2(n_1781),
.B1(n_1732),
.B2(n_206),
.Y(n_2593)
);

NOR3xp33_ASAP7_75t_L g2594 ( 
.A(n_2423),
.B(n_203),
.C(n_205),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2532),
.B(n_208),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2561),
.B(n_2568),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2531),
.B(n_208),
.Y(n_2597)
);

NOR4xp25_ASAP7_75t_L g2598 ( 
.A(n_2447),
.B(n_213),
.C(n_210),
.D(n_212),
.Y(n_2598)
);

AOI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2544),
.A2(n_1781),
.B1(n_1732),
.B2(n_215),
.Y(n_2599)
);

OAI211xp5_ASAP7_75t_L g2600 ( 
.A1(n_2435),
.A2(n_215),
.B(n_210),
.C(n_214),
.Y(n_2600)
);

NOR2xp33_ASAP7_75t_L g2601 ( 
.A(n_2551),
.B(n_214),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2433),
.Y(n_2602)
);

AOI21xp5_ASAP7_75t_L g2603 ( 
.A1(n_2426),
.A2(n_217),
.B(n_219),
.Y(n_2603)
);

AOI221xp5_ASAP7_75t_L g2604 ( 
.A1(n_2479),
.A2(n_221),
.B1(n_217),
.B2(n_220),
.C(n_222),
.Y(n_2604)
);

OA22x2_ASAP7_75t_L g2605 ( 
.A1(n_2524),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_2605)
);

AOI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2469),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2462),
.A2(n_227),
.B1(n_224),
.B2(n_225),
.Y(n_2607)
);

OAI211xp5_ASAP7_75t_L g2608 ( 
.A1(n_2432),
.A2(n_229),
.B(n_227),
.C(n_228),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2548),
.B(n_228),
.Y(n_2609)
);

INVx3_ASAP7_75t_L g2610 ( 
.A(n_2547),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2516),
.B(n_229),
.Y(n_2611)
);

AOI21xp33_ASAP7_75t_L g2612 ( 
.A1(n_2431),
.A2(n_230),
.B(n_231),
.Y(n_2612)
);

OAI22xp5_ASAP7_75t_L g2613 ( 
.A1(n_2425),
.A2(n_233),
.B1(n_230),
.B2(n_232),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2540),
.Y(n_2614)
);

AOI211xp5_ASAP7_75t_L g2615 ( 
.A1(n_2465),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_2615)
);

NAND4xp25_ASAP7_75t_L g2616 ( 
.A(n_2430),
.B(n_238),
.C(n_234),
.D(n_237),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2543),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2549),
.Y(n_2618)
);

OAI211xp5_ASAP7_75t_L g2619 ( 
.A1(n_2474),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_2619)
);

OAI222xp33_ASAP7_75t_L g2620 ( 
.A1(n_2516),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.C1(n_244),
.C2(n_245),
.Y(n_2620)
);

OAI22xp33_ASAP7_75t_L g2621 ( 
.A1(n_2496),
.A2(n_2483),
.B1(n_2560),
.B2(n_2557),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2562),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2486),
.B(n_241),
.Y(n_2623)
);

OAI21xp33_ASAP7_75t_SL g2624 ( 
.A1(n_2494),
.A2(n_243),
.B(n_244),
.Y(n_2624)
);

AOI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2444),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_2625)
);

NOR2xp33_ASAP7_75t_SL g2626 ( 
.A(n_2552),
.B(n_246),
.Y(n_2626)
);

AND4x1_ASAP7_75t_L g2627 ( 
.A(n_2527),
.B(n_2489),
.C(n_2553),
.D(n_2464),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2439),
.Y(n_2628)
);

AOI22xp5_ASAP7_75t_L g2629 ( 
.A1(n_2502),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_2629)
);

OAI21xp5_ASAP7_75t_L g2630 ( 
.A1(n_2536),
.A2(n_248),
.B(n_249),
.Y(n_2630)
);

O2A1O1Ixp33_ASAP7_75t_L g2631 ( 
.A1(n_2533),
.A2(n_253),
.B(n_250),
.C(n_252),
.Y(n_2631)
);

AOI22xp33_ASAP7_75t_SL g2632 ( 
.A1(n_2458),
.A2(n_256),
.B1(n_250),
.B2(n_255),
.Y(n_2632)
);

AOI221xp5_ASAP7_75t_L g2633 ( 
.A1(n_2528),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.C(n_258),
.Y(n_2633)
);

AOI22xp5_ASAP7_75t_L g2634 ( 
.A1(n_2485),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_2564),
.B(n_259),
.Y(n_2635)
);

OAI21xp33_ASAP7_75t_L g2636 ( 
.A1(n_2424),
.A2(n_261),
.B(n_262),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2499),
.Y(n_2637)
);

NOR2x1_ASAP7_75t_L g2638 ( 
.A(n_2475),
.B(n_261),
.Y(n_2638)
);

OAI211xp5_ASAP7_75t_L g2639 ( 
.A1(n_2442),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_2639)
);

A2O1A1Ixp33_ASAP7_75t_L g2640 ( 
.A1(n_2498),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_2640)
);

AOI221xp5_ASAP7_75t_L g2641 ( 
.A1(n_2451),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.C(n_268),
.Y(n_2641)
);

OAI32xp33_ASAP7_75t_L g2642 ( 
.A1(n_2481),
.A2(n_269),
.A3(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2507),
.B(n_271),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_SL g2644 ( 
.A(n_2493),
.B(n_2460),
.Y(n_2644)
);

O2A1O1Ixp5_ASAP7_75t_SL g2645 ( 
.A1(n_2480),
.A2(n_274),
.B(n_271),
.C(n_272),
.Y(n_2645)
);

INVx2_ASAP7_75t_SL g2646 ( 
.A(n_2427),
.Y(n_2646)
);

OAI322xp33_ASAP7_75t_L g2647 ( 
.A1(n_2491),
.A2(n_272),
.A3(n_275),
.B1(n_276),
.B2(n_278),
.C1(n_279),
.C2(n_280),
.Y(n_2647)
);

AOI322xp5_ASAP7_75t_L g2648 ( 
.A1(n_2459),
.A2(n_275),
.A3(n_276),
.B1(n_278),
.B2(n_279),
.C1(n_281),
.C2(n_282),
.Y(n_2648)
);

INVx3_ASAP7_75t_L g2649 ( 
.A(n_2453),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_L g2650 ( 
.A(n_2456),
.B(n_281),
.Y(n_2650)
);

OAI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2537),
.A2(n_282),
.B(n_283),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2509),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_SL g2653 ( 
.A1(n_2436),
.A2(n_284),
.B(n_285),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2492),
.Y(n_2654)
);

AOI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2522),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_2655)
);

AOI31xp33_ASAP7_75t_L g2656 ( 
.A1(n_2513),
.A2(n_289),
.A3(n_286),
.B(n_288),
.Y(n_2656)
);

AOI221xp5_ASAP7_75t_L g2657 ( 
.A1(n_2539),
.A2(n_2554),
.B1(n_2443),
.B2(n_2470),
.C(n_2567),
.Y(n_2657)
);

O2A1O1Ixp33_ASAP7_75t_L g2658 ( 
.A1(n_2517),
.A2(n_292),
.B(n_289),
.C(n_291),
.Y(n_2658)
);

INVx1_ASAP7_75t_SL g2659 ( 
.A(n_2504),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2587),
.B(n_2574),
.Y(n_2660)
);

OAI21xp33_ASAP7_75t_L g2661 ( 
.A1(n_2626),
.A2(n_2511),
.B(n_2518),
.Y(n_2661)
);

NOR3xp33_ASAP7_75t_SL g2662 ( 
.A(n_2572),
.B(n_2468),
.C(n_2514),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2610),
.Y(n_2663)
);

AOI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2652),
.A2(n_2434),
.B1(n_2466),
.B2(n_2461),
.Y(n_2664)
);

AOI221xp5_ASAP7_75t_L g2665 ( 
.A1(n_2598),
.A2(n_2612),
.B1(n_2590),
.B2(n_2594),
.C(n_2616),
.Y(n_2665)
);

AOI221xp5_ASAP7_75t_L g2666 ( 
.A1(n_2575),
.A2(n_2445),
.B1(n_2438),
.B2(n_2495),
.C(n_2478),
.Y(n_2666)
);

AOI21xp33_ASAP7_75t_L g2667 ( 
.A1(n_2578),
.A2(n_2446),
.B(n_2490),
.Y(n_2667)
);

OAI21xp33_ASAP7_75t_SL g2668 ( 
.A1(n_2637),
.A2(n_2449),
.B(n_2488),
.Y(n_2668)
);

OAI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2624),
.A2(n_2638),
.B(n_2603),
.Y(n_2669)
);

INVxp67_ASAP7_75t_L g2670 ( 
.A(n_2595),
.Y(n_2670)
);

AOI21xp5_ASAP7_75t_L g2671 ( 
.A1(n_2644),
.A2(n_2596),
.B(n_2576),
.Y(n_2671)
);

AOI21xp33_ASAP7_75t_SL g2672 ( 
.A1(n_2605),
.A2(n_2503),
.B(n_2437),
.Y(n_2672)
);

NAND4xp25_ASAP7_75t_L g2673 ( 
.A(n_2657),
.B(n_2588),
.C(n_2610),
.D(n_2649),
.Y(n_2673)
);

NAND3xp33_ASAP7_75t_SL g2674 ( 
.A(n_2615),
.B(n_2538),
.C(n_2529),
.Y(n_2674)
);

AOI22xp5_ASAP7_75t_L g2675 ( 
.A1(n_2649),
.A2(n_2608),
.B1(n_2650),
.B2(n_2635),
.Y(n_2675)
);

NOR2x1_ASAP7_75t_L g2676 ( 
.A(n_2620),
.B(n_2473),
.Y(n_2676)
);

CKINVDCx5p33_ASAP7_75t_R g2677 ( 
.A(n_2646),
.Y(n_2677)
);

AOI21xp33_ASAP7_75t_SL g2678 ( 
.A1(n_2656),
.A2(n_2500),
.B(n_2523),
.Y(n_2678)
);

AOI21xp33_ASAP7_75t_SL g2679 ( 
.A1(n_2621),
.A2(n_2520),
.B(n_2450),
.Y(n_2679)
);

AOI21xp33_ASAP7_75t_L g2680 ( 
.A1(n_2577),
.A2(n_2463),
.B(n_2477),
.Y(n_2680)
);

AOI22xp33_ASAP7_75t_SL g2681 ( 
.A1(n_2639),
.A2(n_2570),
.B1(n_2571),
.B2(n_2455),
.Y(n_2681)
);

AOI211xp5_ASAP7_75t_L g2682 ( 
.A1(n_2592),
.A2(n_2613),
.B(n_2619),
.C(n_2600),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2611),
.Y(n_2683)
);

NAND2x1_ASAP7_75t_SL g2684 ( 
.A(n_2591),
.B(n_2506),
.Y(n_2684)
);

XNOR2x2_ASAP7_75t_L g2685 ( 
.A(n_2623),
.B(n_2484),
.Y(n_2685)
);

AOI21xp33_ASAP7_75t_L g2686 ( 
.A1(n_2585),
.A2(n_2471),
.B(n_2476),
.Y(n_2686)
);

AOI21xp33_ASAP7_75t_L g2687 ( 
.A1(n_2583),
.A2(n_2497),
.B(n_2521),
.Y(n_2687)
);

NOR2x1_ASAP7_75t_L g2688 ( 
.A(n_2647),
.B(n_2512),
.Y(n_2688)
);

XNOR2xp5_ASAP7_75t_L g2689 ( 
.A(n_2627),
.B(n_2505),
.Y(n_2689)
);

AOI22xp5_ASAP7_75t_L g2690 ( 
.A1(n_2601),
.A2(n_2541),
.B1(n_2555),
.B2(n_2467),
.Y(n_2690)
);

AOI221xp5_ASAP7_75t_L g2691 ( 
.A1(n_2604),
.A2(n_2534),
.B1(n_2487),
.B2(n_2501),
.C(n_2510),
.Y(n_2691)
);

OAI22xp5_ASAP7_75t_SL g2692 ( 
.A1(n_2581),
.A2(n_2508),
.B1(n_2515),
.B2(n_2556),
.Y(n_2692)
);

AOI21xp5_ASAP7_75t_L g2693 ( 
.A1(n_2631),
.A2(n_2545),
.B(n_2519),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2648),
.B(n_2472),
.Y(n_2694)
);

AOI221xp5_ASAP7_75t_L g2695 ( 
.A1(n_2579),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.C(n_294),
.Y(n_2695)
);

AOI21xp33_ASAP7_75t_L g2696 ( 
.A1(n_2584),
.A2(n_293),
.B(n_294),
.Y(n_2696)
);

OAI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2593),
.A2(n_295),
.B(n_296),
.Y(n_2697)
);

AOI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2573),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_2698)
);

OAI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_2625),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_2699)
);

A2O1A1Ixp33_ASAP7_75t_L g2700 ( 
.A1(n_2658),
.A2(n_308),
.B(n_304),
.C(n_307),
.Y(n_2700)
);

BUFx2_ASAP7_75t_L g2701 ( 
.A(n_2640),
.Y(n_2701)
);

AOI222xp33_ASAP7_75t_L g2702 ( 
.A1(n_2580),
.A2(n_304),
.B1(n_309),
.B2(n_311),
.C1(n_313),
.C2(n_314),
.Y(n_2702)
);

AOI221xp5_ASAP7_75t_L g2703 ( 
.A1(n_2633),
.A2(n_309),
.B1(n_311),
.B2(n_313),
.C(n_314),
.Y(n_2703)
);

AOI22xp5_ASAP7_75t_L g2704 ( 
.A1(n_2602),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_2704)
);

OAI22xp33_ASAP7_75t_L g2705 ( 
.A1(n_2597),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2643),
.Y(n_2706)
);

AOI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2659),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_2707)
);

AOI211xp5_ASAP7_75t_L g2708 ( 
.A1(n_2589),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_2708)
);

OAI22xp33_ASAP7_75t_SL g2709 ( 
.A1(n_2609),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2606),
.Y(n_2710)
);

AOI22xp5_ASAP7_75t_L g2711 ( 
.A1(n_2654),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_2711)
);

NOR2xp67_ASAP7_75t_L g2712 ( 
.A(n_2629),
.B(n_325),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2636),
.Y(n_2713)
);

OAI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2630),
.A2(n_327),
.B(n_328),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2634),
.Y(n_2715)
);

XNOR2xp5_ASAP7_75t_L g2716 ( 
.A(n_2655),
.B(n_328),
.Y(n_2716)
);

OAI21xp5_ASAP7_75t_L g2717 ( 
.A1(n_2651),
.A2(n_329),
.B(n_331),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2660),
.Y(n_2718)
);

AOI211xp5_ASAP7_75t_SL g2719 ( 
.A1(n_2667),
.A2(n_2653),
.B(n_2614),
.C(n_2618),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2677),
.Y(n_2720)
);

AOI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2669),
.A2(n_2622),
.B(n_2617),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2663),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2701),
.Y(n_2723)
);

AOI221xp5_ASAP7_75t_L g2724 ( 
.A1(n_2673),
.A2(n_2628),
.B1(n_2641),
.B2(n_2642),
.C(n_2632),
.Y(n_2724)
);

O2A1O1Ixp33_ASAP7_75t_L g2725 ( 
.A1(n_2700),
.A2(n_2709),
.B(n_2586),
.C(n_2705),
.Y(n_2725)
);

HB1xp67_ASAP7_75t_L g2726 ( 
.A(n_2676),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2683),
.Y(n_2727)
);

OAI31xp33_ASAP7_75t_L g2728 ( 
.A1(n_2661),
.A2(n_2645),
.A3(n_2599),
.B(n_2607),
.Y(n_2728)
);

NOR3xp33_ASAP7_75t_L g2729 ( 
.A(n_2671),
.B(n_2670),
.C(n_2687),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2674),
.B(n_2582),
.Y(n_2730)
);

XNOR2xp5_ASAP7_75t_L g2731 ( 
.A(n_2689),
.B(n_329),
.Y(n_2731)
);

AOI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2688),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_2732)
);

XOR2xp5_ASAP7_75t_L g2733 ( 
.A(n_2675),
.B(n_334),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2684),
.Y(n_2734)
);

AOI22xp5_ASAP7_75t_L g2735 ( 
.A1(n_2665),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_2735)
);

AOI31xp33_ASAP7_75t_L g2736 ( 
.A1(n_2682),
.A2(n_339),
.A3(n_336),
.B(n_338),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2716),
.Y(n_2737)
);

OAI211xp5_ASAP7_75t_L g2738 ( 
.A1(n_2664),
.A2(n_342),
.B(n_338),
.C(n_340),
.Y(n_2738)
);

OAI22xp33_ASAP7_75t_SL g2739 ( 
.A1(n_2694),
.A2(n_346),
.B1(n_343),
.B2(n_344),
.Y(n_2739)
);

AOI322xp5_ASAP7_75t_L g2740 ( 
.A1(n_2662),
.A2(n_343),
.A3(n_344),
.B1(n_346),
.B2(n_347),
.C1(n_348),
.C2(n_349),
.Y(n_2740)
);

AOI31xp33_ASAP7_75t_L g2741 ( 
.A1(n_2682),
.A2(n_350),
.A3(n_347),
.B(n_348),
.Y(n_2741)
);

OAI211xp5_ASAP7_75t_L g2742 ( 
.A1(n_2668),
.A2(n_352),
.B(n_350),
.C(n_351),
.Y(n_2742)
);

OAI211xp5_ASAP7_75t_SL g2743 ( 
.A1(n_2666),
.A2(n_354),
.B(n_351),
.C(n_352),
.Y(n_2743)
);

NOR3x1_ASAP7_75t_L g2744 ( 
.A(n_2714),
.B(n_2717),
.C(n_2697),
.Y(n_2744)
);

AO21x1_ASAP7_75t_L g2745 ( 
.A1(n_2699),
.A2(n_356),
.B(n_357),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2698),
.B(n_356),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2712),
.Y(n_2747)
);

AOI221xp5_ASAP7_75t_L g2748 ( 
.A1(n_2672),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.C(n_361),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2713),
.B(n_358),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2707),
.B(n_362),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2702),
.B(n_364),
.Y(n_2751)
);

AOI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2715),
.A2(n_2710),
.B1(n_2692),
.B2(n_2690),
.Y(n_2752)
);

AOI221xp5_ASAP7_75t_L g2753 ( 
.A1(n_2678),
.A2(n_364),
.B1(n_366),
.B2(n_369),
.C(n_370),
.Y(n_2753)
);

OA22x2_ASAP7_75t_L g2754 ( 
.A1(n_2732),
.A2(n_2706),
.B1(n_2704),
.B2(n_2711),
.Y(n_2754)
);

OAI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2734),
.A2(n_2681),
.B1(n_2708),
.B2(n_2703),
.Y(n_2755)
);

AOI22xp33_ASAP7_75t_SL g2756 ( 
.A1(n_2726),
.A2(n_2685),
.B1(n_2693),
.B2(n_2679),
.Y(n_2756)
);

AOI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2720),
.A2(n_2691),
.B1(n_2695),
.B2(n_2680),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2731),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2733),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2749),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2740),
.B(n_2696),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2736),
.B(n_2741),
.Y(n_2762)
);

AOI22xp5_ASAP7_75t_L g2763 ( 
.A1(n_2723),
.A2(n_2686),
.B1(n_371),
.B2(n_366),
.Y(n_2763)
);

INVxp33_ASAP7_75t_SL g2764 ( 
.A(n_2752),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2729),
.A2(n_373),
.B1(n_370),
.B2(n_372),
.Y(n_2765)
);

NOR2x1_ASAP7_75t_L g2766 ( 
.A(n_2742),
.B(n_372),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2745),
.Y(n_2767)
);

NOR2xp67_ASAP7_75t_L g2768 ( 
.A(n_2738),
.B(n_374),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2739),
.Y(n_2769)
);

NOR2x1_ASAP7_75t_L g2770 ( 
.A(n_2747),
.B(n_374),
.Y(n_2770)
);

INVx3_ASAP7_75t_L g2771 ( 
.A(n_2722),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2743),
.B(n_2739),
.Y(n_2772)
);

AOI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2730),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2770),
.Y(n_2774)
);

NOR2x1p5_ASAP7_75t_L g2775 ( 
.A(n_2771),
.B(n_2751),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2766),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2769),
.Y(n_2777)
);

INVxp67_ASAP7_75t_SL g2778 ( 
.A(n_2767),
.Y(n_2778)
);

NOR2xp67_ASAP7_75t_L g2779 ( 
.A(n_2762),
.B(n_2721),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2772),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2761),
.Y(n_2781)
);

XNOR2xp5_ASAP7_75t_L g2782 ( 
.A(n_2764),
.B(n_2724),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2760),
.B(n_2727),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2754),
.Y(n_2784)
);

NOR2x1_ASAP7_75t_L g2785 ( 
.A(n_2768),
.B(n_2718),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2765),
.Y(n_2786)
);

CKINVDCx5p33_ASAP7_75t_R g2787 ( 
.A(n_2756),
.Y(n_2787)
);

XNOR2xp5_ASAP7_75t_L g2788 ( 
.A(n_2757),
.B(n_2735),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2758),
.Y(n_2789)
);

NAND4xp75_ASAP7_75t_L g2790 ( 
.A(n_2763),
.B(n_2744),
.C(n_2748),
.D(n_2737),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2787),
.A2(n_2755),
.B1(n_2759),
.B2(n_2746),
.Y(n_2791)
);

OAI221xp5_ASAP7_75t_L g2792 ( 
.A1(n_2778),
.A2(n_2728),
.B1(n_2725),
.B2(n_2719),
.C(n_2773),
.Y(n_2792)
);

OAI211xp5_ASAP7_75t_L g2793 ( 
.A1(n_2778),
.A2(n_2784),
.B(n_2779),
.C(n_2774),
.Y(n_2793)
);

OAI211xp5_ASAP7_75t_SL g2794 ( 
.A1(n_2785),
.A2(n_2750),
.B(n_2753),
.C(n_378),
.Y(n_2794)
);

OAI221xp5_ASAP7_75t_SL g2795 ( 
.A1(n_2782),
.A2(n_376),
.B1(n_377),
.B2(n_378),
.C(n_379),
.Y(n_2795)
);

NAND4xp25_ASAP7_75t_L g2796 ( 
.A(n_2779),
.B(n_382),
.C(n_380),
.D(n_381),
.Y(n_2796)
);

INVx1_ASAP7_75t_SL g2797 ( 
.A(n_2776),
.Y(n_2797)
);

OAI211xp5_ASAP7_75t_L g2798 ( 
.A1(n_2780),
.A2(n_383),
.B(n_380),
.C(n_382),
.Y(n_2798)
);

AND2x4_ASAP7_75t_L g2799 ( 
.A(n_2783),
.B(n_384),
.Y(n_2799)
);

OAI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2788),
.A2(n_384),
.B(n_385),
.Y(n_2800)
);

OAI211xp5_ASAP7_75t_L g2801 ( 
.A1(n_2781),
.A2(n_385),
.B(n_386),
.C(n_387),
.Y(n_2801)
);

O2A1O1Ixp33_ASAP7_75t_L g2802 ( 
.A1(n_2777),
.A2(n_386),
.B(n_387),
.C(n_389),
.Y(n_2802)
);

HB1xp67_ASAP7_75t_L g2803 ( 
.A(n_2775),
.Y(n_2803)
);

INVxp67_ASAP7_75t_SL g2804 ( 
.A(n_2789),
.Y(n_2804)
);

NOR3xp33_ASAP7_75t_L g2805 ( 
.A(n_2790),
.B(n_390),
.C(n_391),
.Y(n_2805)
);

AOI221xp5_ASAP7_75t_L g2806 ( 
.A1(n_2786),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.C(n_394),
.Y(n_2806)
);

OAI21xp33_ASAP7_75t_SL g2807 ( 
.A1(n_2778),
.A2(n_392),
.B(n_394),
.Y(n_2807)
);

OAI221xp5_ASAP7_75t_L g2808 ( 
.A1(n_2778),
.A2(n_395),
.B1(n_397),
.B2(n_398),
.C(n_399),
.Y(n_2808)
);

HB1xp67_ASAP7_75t_L g2809 ( 
.A(n_2774),
.Y(n_2809)
);

AND2x4_ASAP7_75t_L g2810 ( 
.A(n_2804),
.B(n_397),
.Y(n_2810)
);

HB1xp67_ASAP7_75t_L g2811 ( 
.A(n_2799),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2799),
.Y(n_2812)
);

OAI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2797),
.A2(n_399),
.B1(n_400),
.B2(n_402),
.Y(n_2813)
);

HB1xp67_ASAP7_75t_L g2814 ( 
.A(n_2807),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2809),
.Y(n_2815)
);

AND2x2_ASAP7_75t_SL g2816 ( 
.A(n_2805),
.B(n_402),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2803),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2796),
.Y(n_2818)
);

XNOR2x1_ASAP7_75t_L g2819 ( 
.A(n_2791),
.B(n_403),
.Y(n_2819)
);

XNOR2xp5_ASAP7_75t_L g2820 ( 
.A(n_2792),
.B(n_403),
.Y(n_2820)
);

NAND3xp33_ASAP7_75t_L g2821 ( 
.A(n_2793),
.B(n_405),
.C(n_406),
.Y(n_2821)
);

OAI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2794),
.A2(n_406),
.B(n_407),
.Y(n_2822)
);

NOR2x1_ASAP7_75t_L g2823 ( 
.A(n_2801),
.B(n_407),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2798),
.Y(n_2824)
);

NOR3xp33_ASAP7_75t_L g2825 ( 
.A(n_2795),
.B(n_408),
.C(n_409),
.Y(n_2825)
);

AND2x2_ASAP7_75t_SL g2826 ( 
.A(n_2806),
.B(n_408),
.Y(n_2826)
);

INVx1_ASAP7_75t_SL g2827 ( 
.A(n_2800),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2802),
.Y(n_2828)
);

OR2x2_ASAP7_75t_L g2829 ( 
.A(n_2808),
.B(n_410),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2814),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2810),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2811),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2810),
.Y(n_2833)
);

XNOR2xp5_ASAP7_75t_L g2834 ( 
.A(n_2820),
.B(n_410),
.Y(n_2834)
);

NAND2x1_ASAP7_75t_L g2835 ( 
.A(n_2812),
.B(n_411),
.Y(n_2835)
);

OR2x2_ASAP7_75t_L g2836 ( 
.A(n_2815),
.B(n_412),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2819),
.Y(n_2837)
);

OA22x2_ASAP7_75t_L g2838 ( 
.A1(n_2822),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_R g2839 ( 
.A(n_2828),
.B(n_413),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2821),
.Y(n_2840)
);

CKINVDCx5p33_ASAP7_75t_R g2841 ( 
.A(n_2817),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2816),
.Y(n_2842)
);

NOR2xp67_ASAP7_75t_L g2843 ( 
.A(n_2813),
.B(n_414),
.Y(n_2843)
);

INVx4_ASAP7_75t_L g2844 ( 
.A(n_2824),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2835),
.Y(n_2845)
);

INVx5_ASAP7_75t_L g2846 ( 
.A(n_2844),
.Y(n_2846)
);

NAND3xp33_ASAP7_75t_SL g2847 ( 
.A(n_2839),
.B(n_2827),
.C(n_2825),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2836),
.Y(n_2848)
);

OAI22xp5_ASAP7_75t_SL g2849 ( 
.A1(n_2830),
.A2(n_2826),
.B1(n_2818),
.B2(n_2823),
.Y(n_2849)
);

INVx1_ASAP7_75t_SL g2850 ( 
.A(n_2831),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2832),
.B(n_2829),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2838),
.Y(n_2852)
);

OAI22xp5_ASAP7_75t_SL g2853 ( 
.A1(n_2841),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_2853)
);

HB1xp67_ASAP7_75t_L g2854 ( 
.A(n_2833),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2834),
.Y(n_2855)
);

AOI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2834),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_2856)
);

NAND3xp33_ASAP7_75t_L g2857 ( 
.A(n_2840),
.B(n_2843),
.C(n_2842),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2837),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2856),
.B(n_418),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2854),
.Y(n_2860)
);

NOR3xp33_ASAP7_75t_L g2861 ( 
.A(n_2847),
.B(n_418),
.C(n_420),
.Y(n_2861)
);

INVxp67_ASAP7_75t_L g2862 ( 
.A(n_2845),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2850),
.B(n_2846),
.Y(n_2863)
);

AO22x2_ASAP7_75t_L g2864 ( 
.A1(n_2852),
.A2(n_420),
.B1(n_421),
.B2(n_422),
.Y(n_2864)
);

OR2x2_ASAP7_75t_L g2865 ( 
.A(n_2858),
.B(n_422),
.Y(n_2865)
);

OAI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2846),
.A2(n_424),
.B1(n_426),
.B2(n_427),
.Y(n_2866)
);

AND2x4_ASAP7_75t_L g2867 ( 
.A(n_2851),
.B(n_424),
.Y(n_2867)
);

CKINVDCx20_ASAP7_75t_R g2868 ( 
.A(n_2849),
.Y(n_2868)
);

OAI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_2857),
.A2(n_426),
.B(n_427),
.Y(n_2869)
);

AOI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2855),
.A2(n_2848),
.B1(n_2853),
.B2(n_430),
.Y(n_2870)
);

OR2x2_ASAP7_75t_L g2871 ( 
.A(n_2850),
.B(n_428),
.Y(n_2871)
);

OAI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2850),
.A2(n_429),
.B1(n_431),
.B2(n_432),
.Y(n_2872)
);

AO22x2_ASAP7_75t_L g2873 ( 
.A1(n_2845),
.A2(n_432),
.B1(n_433),
.B2(n_434),
.Y(n_2873)
);

OAI22xp5_ASAP7_75t_L g2874 ( 
.A1(n_2860),
.A2(n_433),
.B1(n_435),
.B2(n_437),
.Y(n_2874)
);

CKINVDCx20_ASAP7_75t_R g2875 ( 
.A(n_2868),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2871),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2861),
.B(n_437),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2873),
.Y(n_2878)
);

BUFx2_ASAP7_75t_L g2879 ( 
.A(n_2864),
.Y(n_2879)
);

AOI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2863),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_2880)
);

AOI22xp5_ASAP7_75t_L g2881 ( 
.A1(n_2862),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_2881)
);

OAI22x1_ASAP7_75t_L g2882 ( 
.A1(n_2870),
.A2(n_441),
.B1(n_443),
.B2(n_444),
.Y(n_2882)
);

CKINVDCx20_ASAP7_75t_R g2883 ( 
.A(n_2859),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2873),
.Y(n_2884)
);

HB1xp67_ASAP7_75t_L g2885 ( 
.A(n_2864),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2885),
.Y(n_2886)
);

OAI21xp33_ASAP7_75t_L g2887 ( 
.A1(n_2875),
.A2(n_2869),
.B(n_2872),
.Y(n_2887)
);

AOI22xp5_ASAP7_75t_L g2888 ( 
.A1(n_2883),
.A2(n_2866),
.B1(n_2867),
.B2(n_2865),
.Y(n_2888)
);

OAI22xp5_ASAP7_75t_L g2889 ( 
.A1(n_2877),
.A2(n_444),
.B1(n_445),
.B2(n_447),
.Y(n_2889)
);

CKINVDCx20_ASAP7_75t_R g2890 ( 
.A(n_2879),
.Y(n_2890)
);

OAI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2876),
.A2(n_448),
.B1(n_451),
.B2(n_452),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2882),
.Y(n_2892)
);

OAI21xp33_ASAP7_75t_L g2893 ( 
.A1(n_2878),
.A2(n_448),
.B(n_451),
.Y(n_2893)
);

OAI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2884),
.A2(n_453),
.B(n_454),
.Y(n_2894)
);

AO22x2_ASAP7_75t_L g2895 ( 
.A1(n_2874),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_2895)
);

AO21x2_ASAP7_75t_L g2896 ( 
.A1(n_2880),
.A2(n_456),
.B(n_457),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2893),
.B(n_2881),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2896),
.B(n_457),
.Y(n_2898)
);

AOI22xp5_ASAP7_75t_L g2899 ( 
.A1(n_2890),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2886),
.B(n_2895),
.Y(n_2900)
);

AOI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2887),
.A2(n_459),
.B(n_461),
.Y(n_2901)
);

AOI21xp33_ASAP7_75t_L g2902 ( 
.A1(n_2892),
.A2(n_462),
.B(n_463),
.Y(n_2902)
);

AOI21x1_ASAP7_75t_L g2903 ( 
.A1(n_2889),
.A2(n_463),
.B(n_464),
.Y(n_2903)
);

AOI222xp33_ASAP7_75t_L g2904 ( 
.A1(n_2894),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.C1(n_468),
.C2(n_472),
.Y(n_2904)
);

OAI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2888),
.A2(n_465),
.B(n_466),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2891),
.A2(n_467),
.B(n_472),
.Y(n_2906)
);

AOI22xp5_ASAP7_75t_L g2907 ( 
.A1(n_2900),
.A2(n_474),
.B1(n_475),
.B2(n_476),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2898),
.Y(n_2908)
);

AOI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2906),
.A2(n_474),
.B1(n_478),
.B2(n_479),
.Y(n_2909)
);

AOI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2904),
.A2(n_479),
.B1(n_480),
.B2(n_481),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2903),
.Y(n_2911)
);

AOI22xp5_ASAP7_75t_L g2912 ( 
.A1(n_2910),
.A2(n_2909),
.B1(n_2897),
.B2(n_2908),
.Y(n_2912)
);

AOI22xp33_ASAP7_75t_L g2913 ( 
.A1(n_2911),
.A2(n_2901),
.B1(n_2905),
.B2(n_2902),
.Y(n_2913)
);

AOI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2907),
.A2(n_2899),
.B1(n_481),
.B2(n_482),
.Y(n_2914)
);

OR2x2_ASAP7_75t_L g2915 ( 
.A(n_2914),
.B(n_480),
.Y(n_2915)
);

AOI221xp5_ASAP7_75t_L g2916 ( 
.A1(n_2915),
.A2(n_2913),
.B1(n_2912),
.B2(n_485),
.C(n_486),
.Y(n_2916)
);

AOI211xp5_ASAP7_75t_L g2917 ( 
.A1(n_2916),
.A2(n_483),
.B(n_484),
.C(n_488),
.Y(n_2917)
);


endmodule