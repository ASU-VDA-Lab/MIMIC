module fake_jpeg_25446_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_34),
.B1(n_61),
.B2(n_63),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

BUFx2_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_29),
.B1(n_28),
.B2(n_42),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_37),
.B1(n_28),
.B2(n_29),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_33),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_63),
.C(n_43),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_32),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_34),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_68),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_83),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_61),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_76),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_30),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_29),
.B1(n_17),
.B2(n_18),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_39),
.Y(n_107)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_96),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_108),
.B(n_110),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_53),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_55),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_63),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_66),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_16),
.B(n_23),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_111),
.B(n_93),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_72),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_82),
.B1(n_30),
.B2(n_23),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_68),
.C(n_66),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_79),
.C(n_83),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_121),
.A2(n_132),
.B(n_114),
.Y(n_166)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_80),
.B1(n_64),
.B2(n_87),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_140),
.B1(n_144),
.B2(n_101),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_133),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_37),
.B1(n_76),
.B2(n_64),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_135),
.B1(n_146),
.B2(n_101),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_25),
.B1(n_106),
.B2(n_89),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_100),
.B1(n_97),
.B2(n_104),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_136),
.B1(n_42),
.B2(n_38),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_66),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_78),
.B1(n_77),
.B2(n_46),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_97),
.B1(n_104),
.B2(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_138),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_98),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_9),
.C(n_11),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

AO21x2_ASAP7_75t_SL g145 ( 
.A1(n_94),
.A2(n_89),
.B(n_77),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_106),
.B(n_108),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_78),
.B1(n_44),
.B2(n_69),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_108),
.A3(n_92),
.B1(n_71),
.B2(n_75),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_148),
.A2(n_172),
.B(n_32),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_150),
.B1(n_160),
.B2(n_175),
.Y(n_186)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_155),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_120),
.B(n_121),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_141),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_158),
.C(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_122),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_114),
.C(n_91),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_99),
.B1(n_83),
.B2(n_87),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_122),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_165),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_41),
.B(n_32),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_95),
.Y(n_167)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_95),
.B1(n_44),
.B2(n_38),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_171),
.A2(n_127),
.B1(n_125),
.B2(n_73),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_87),
.B(n_1),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_62),
.B1(n_20),
.B2(n_39),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_132),
.B1(n_73),
.B2(n_67),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_20),
.B1(n_24),
.B2(n_27),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_125),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_178),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_194),
.B1(n_172),
.B2(n_152),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_192),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_201),
.C(n_154),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_204),
.B1(n_161),
.B2(n_171),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_142),
.B1(n_20),
.B2(n_67),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_191),
.A2(n_159),
.B1(n_151),
.B2(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_41),
.Y(n_195)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_196),
.A2(n_197),
.B(n_170),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_200),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_52),
.C(n_19),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_169),
.A2(n_19),
.B1(n_27),
.B2(n_24),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_173),
.B1(n_22),
.B2(n_31),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_19),
.B1(n_27),
.B2(n_24),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_31),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_201),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_0),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_178),
.C(n_181),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_153),
.B1(n_174),
.B2(n_170),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_216),
.B(n_218),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_186),
.B1(n_179),
.B2(n_202),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_220),
.B1(n_189),
.B2(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_219),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_152),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_167),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_222),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_199),
.A2(n_168),
.B1(n_8),
.B2(n_10),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_231),
.B(n_180),
.Y(n_247)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_229),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_226),
.A2(n_215),
.B1(n_230),
.B2(n_220),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_22),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_178),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_198),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_0),
.B(n_1),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_8),
.C(n_13),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_248),
.C(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_246),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_223),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_181),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_10),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_179),
.B(n_182),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_253),
.B(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_247),
.A2(n_207),
.B(n_226),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_188),
.C(n_182),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_190),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_221),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_262),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_214),
.CI(n_227),
.CON(n_260),
.SN(n_260)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_237),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_188),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_207),
.C(n_209),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_268),
.C(n_247),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_237),
.B(n_239),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_252),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_6),
.C(n_13),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_265),
.A2(n_240),
.B1(n_251),
.B2(n_245),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_272),
.A2(n_280),
.B1(n_11),
.B2(n_13),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_4),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_4),
.B(n_5),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_242),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_281),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_279),
.A2(n_11),
.B(n_12),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_238),
.C(n_249),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_284),
.C(n_259),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_238),
.C(n_235),
.Y(n_284)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_288),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_271),
.B(n_270),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_289),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_255),
.C(n_256),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_267),
.C(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_273),
.B(n_260),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_6),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_293),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_295),
.B(n_280),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_5),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_277),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_305),
.C(n_290),
.Y(n_308)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_283),
.B(n_277),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_12),
.B1(n_14),
.B2(n_2),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_3),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_312),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_14),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_310),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_304),
.A2(n_14),
.B(n_3),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_313),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_307),
.B(n_299),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_303),
.C(n_300),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_303),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_319),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_315),
.B(n_317),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_314),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_311),
.Y(n_323)
);


endmodule