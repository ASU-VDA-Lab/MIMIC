module fake_netlist_6_3582_n_29 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_8, n_29);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_8;

output n_29;

wire n_16;
wire n_18;
wire n_21;
wire n_10;
wire n_24;
wire n_15;
wire n_27;
wire n_14;
wire n_22;
wire n_26;
wire n_13;
wire n_11;
wire n_28;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_19;
wire n_25;

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_SL g12 ( 
.A(n_8),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NAND3xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_1),
.C(n_2),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

AND2x4_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_11),
.Y(n_19)
);

OAI31xp33_ASAP7_75t_SL g20 ( 
.A1(n_18),
.A2(n_15),
.A3(n_12),
.B(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_11),
.B(n_13),
.C(n_16),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

OAI221xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.C(n_4),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_16),
.B1(n_6),
.B2(n_9),
.Y(n_25)
);

OAI221xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_3),
.B1(n_4),
.B2(n_21),
.C(n_23),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_R g29 ( 
.A1(n_28),
.A2(n_24),
.B1(n_27),
.B2(n_3),
.Y(n_29)
);


endmodule