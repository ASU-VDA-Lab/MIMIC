module real_jpeg_25049_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_1),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_88),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_88),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_1),
.A2(n_66),
.B1(n_69),
.B2(n_88),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_47),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_2),
.A2(n_47),
.B1(n_66),
.B2(n_69),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_6),
.A2(n_45),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_6),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_119),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_119),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_6),
.A2(n_66),
.B1(n_69),
.B2(n_119),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_7),
.A2(n_46),
.B1(n_79),
.B2(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_7),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_172),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_172),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_7),
.A2(n_66),
.B1(n_69),
.B2(n_172),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_8),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_56),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_56),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_8),
.A2(n_56),
.B1(n_66),
.B2(n_69),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_11),
.B(n_58),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_11),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_54),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_11),
.B(n_28),
.C(n_30),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_225),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_11),
.B(n_37),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_225),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_11),
.B(n_66),
.C(n_68),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_11),
.A2(n_101),
.B(n_286),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_13),
.A2(n_46),
.B1(n_52),
.B2(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_13),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_143),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_143),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_13),
.A2(n_66),
.B1(n_69),
.B2(n_143),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_14),
.A2(n_46),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_14),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_80),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_80),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_14),
.A2(n_66),
.B1(n_69),
.B2(n_80),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_15),
.A2(n_40),
.B1(n_66),
.B2(n_69),
.Y(n_106)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_16),
.Y(n_105)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_16),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_16),
.A2(n_194),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_95),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_94),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_21),
.B(n_81),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_62),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_41),
.B1(n_60),
.B2(n_61),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_37),
.B(n_38),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_24),
.A2(n_37),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_24),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_24),
.A2(n_37),
.B1(n_190),
.B2(n_218),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_25),
.A2(n_26),
.B1(n_39),
.B2(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_25),
.A2(n_26),
.B1(n_92),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_25),
.A2(n_26),
.B1(n_123),
.B2(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_25),
.A2(n_189),
.B(n_191),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_25),
.A2(n_191),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_26),
.A2(n_139),
.B(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_26),
.A2(n_175),
.B(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_27),
.A2(n_28),
.B1(n_67),
.B2(n_68),
.Y(n_71)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_28),
.B(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_34),
.B1(n_50),
.B2(n_51),
.Y(n_54)
);

AOI32xp33_ASAP7_75t_L g200 ( 
.A1(n_33),
.A2(n_51),
.A3(n_52),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_34),
.B(n_50),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_34),
.B(n_249),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_37),
.B(n_176),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_54),
.B2(n_55),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_53),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_45),
.A2(n_225),
.B(n_226),
.Y(n_224)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_48),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_48),
.A2(n_54),
.B1(n_142),
.B2(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_48),
.A2(n_145),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_77),
.B1(n_78),
.B2(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_53),
.A2(n_87),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_53),
.B(n_117),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_53),
.A2(n_115),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_74),
.C(n_76),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_74),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_86),
.C(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_63),
.A2(n_85),
.B1(n_90),
.B2(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_70),
.B(n_72),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_70),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_64),
.A2(n_70),
.B1(n_109),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_64),
.A2(n_70),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_64),
.B(n_222),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_65),
.A2(n_73),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_65),
.A2(n_125),
.B1(n_137),
.B2(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_65),
.A2(n_182),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_65),
.A2(n_221),
.B(n_259),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_65),
.B(n_225),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_69),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_70),
.B(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_77),
.A2(n_141),
.B(n_144),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_89),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_82),
.A2(n_86),
.B1(n_155),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_86),
.A2(n_152),
.B1(n_153),
.B2(n_155),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_86),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_89),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI31xp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_156),
.A3(n_162),
.B(n_342),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_146),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_97),
.B(n_146),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_120),
.C(n_128),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_98),
.A2(n_120),
.B1(n_121),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_98),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_111),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_99),
.A2(n_100),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_107),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_100),
.A2(n_107),
.B1(n_108),
.B2(n_112),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B(n_106),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_103),
.B1(n_106),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_101),
.A2(n_103),
.B1(n_133),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_101),
.A2(n_196),
.B1(n_198),
.B2(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_101),
.B(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_101),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_102),
.Y(n_254)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_105),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_105),
.B(n_225),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_124),
.B(n_127),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_124),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_125),
.A2(n_273),
.B(n_274),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_125),
.A2(n_274),
.B(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_128),
.A2(n_129),
.B1(n_337),
.B2(n_339),
.Y(n_336)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_138),
.C(n_140),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_130),
.A2(n_131),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_138),
.B(n_140),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_149),
.C(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_157),
.A2(n_343),
.B(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_158),
.B(n_161),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_335),
.B(n_341),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_210),
.B(n_334),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_203),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_165),
.B(n_203),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_183),
.C(n_185),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_166),
.A2(n_167),
.B1(n_183),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_177),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_173),
.C(n_177),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_178),
.B(n_181),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_183),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_185),
.B(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_192),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_188),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_200),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_200),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_198),
.A2(n_299),
.B(n_307),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_205),
.B(n_206),
.C(n_209),
.Y(n_340)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_241),
.B(n_328),
.C(n_333),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_235),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_227),
.C(n_228),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_213),
.A2(n_214),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_219),
.C(n_223),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_227),
.B(n_228),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.C(n_233),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_268),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_322),
.B(n_327),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_275),
.B(n_321),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_264),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_246),
.B(n_264),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_257),
.C(n_261),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_247),
.B(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_250),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B(n_255),
.Y(n_250)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_257),
.A2(n_261),
.B1(n_262),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_269),
.B2(n_270),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_271),
.C(n_272),
.Y(n_326)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_315),
.B(n_320),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_295),
.B(n_314),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_289),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_289),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_284),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_283),
.C(n_284),
.Y(n_319)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_285),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_291),
.B1(n_293),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_293),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_303),
.B(n_313),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_301),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_301),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_308),
.B(n_312),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_306),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_326),
.Y(n_327)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_340),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_340),
.Y(n_341)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_337),
.Y(n_339)
);


endmodule