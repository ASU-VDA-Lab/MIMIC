module fake_netlist_6_40_n_4803 (n_992, n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_1030, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_1008, n_1027, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_1033, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_933, n_740, n_1038, n_578, n_703, n_1003, n_144, n_365, n_978, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_1044, n_951, n_783, n_106, n_725, n_952, n_999, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_994, n_677, n_969, n_988, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_974, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_1020, n_180, n_1009, n_1042, n_62, n_628, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_1032, n_845, n_255, n_807, n_1036, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_893, n_214, n_925, n_485, n_67, n_15, n_1026, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_1024, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_1018, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_1037, n_72, n_721, n_996, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_1015, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_56, n_763, n_1057, n_360, n_945, n_977, n_603, n_1005, n_119, n_991, n_957, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_987, n_641, n_822, n_693, n_1056, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_989, n_797, n_666, n_1016, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_1035, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_1004, n_1017, n_494, n_539, n_493, n_397, n_155, n_1022, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_1049, n_576, n_1028, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_976, n_490, n_803, n_290, n_220, n_809, n_1043, n_1011, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_986, n_80, n_734, n_708, n_196, n_919, n_402, n_352, n_917, n_668, n_478, n_626, n_990, n_574, n_779, n_9, n_800, n_929, n_460, n_107, n_907, n_854, n_6, n_1058, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_293, n_1054, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_998, n_16, n_1046, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_924, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_962, n_1000, n_279, n_686, n_796, n_1041, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_984, n_411, n_503, n_716, n_152, n_623, n_1048, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_1021, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_981, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_985, n_589, n_860, n_481, n_788, n_819, n_939, n_997, n_821, n_325, n_938, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_982, n_561, n_33, n_477, n_549, n_980, n_533, n_954, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_979, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_993, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_1051, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_249, n_201, n_386, n_764, n_1039, n_556, n_159, n_1034, n_157, n_162, n_692, n_733, n_754, n_941, n_975, n_1031, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_560, n_1014, n_753, n_642, n_995, n_276, n_569, n_441, n_221, n_811, n_882, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_1053, n_530, n_277, n_520, n_1029, n_418, n_113, n_618, n_1055, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_1047, n_1010, n_355, n_426, n_317, n_149, n_1040, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_1052, n_502, n_328, n_672, n_534, n_488, n_429, n_1006, n_373, n_1012, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_1045, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_1002, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_1019, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_983, n_64, n_288, n_427, n_1059, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_1001, n_60, n_361, n_508, n_663, n_856, n_1050, n_379, n_170, n_778, n_1025, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_1013, n_1023, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_1007, n_51, n_649, n_283, n_4803);

input n_992;
input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_1030;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_1008;
input n_1027;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_1033;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_933;
input n_740;
input n_1038;
input n_578;
input n_703;
input n_1003;
input n_144;
input n_365;
input n_978;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_1044;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_994;
input n_677;
input n_969;
input n_988;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_974;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_1020;
input n_180;
input n_1009;
input n_1042;
input n_62;
input n_628;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_1032;
input n_845;
input n_255;
input n_807;
input n_1036;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_893;
input n_214;
input n_925;
input n_485;
input n_67;
input n_15;
input n_1026;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_1024;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_1018;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_1037;
input n_72;
input n_721;
input n_996;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_1015;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_56;
input n_763;
input n_1057;
input n_360;
input n_945;
input n_977;
input n_603;
input n_1005;
input n_119;
input n_991;
input n_957;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_987;
input n_641;
input n_822;
input n_693;
input n_1056;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_989;
input n_797;
input n_666;
input n_1016;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_1035;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_1004;
input n_1017;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_1022;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_1049;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_976;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_1043;
input n_1011;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_986;
input n_80;
input n_734;
input n_708;
input n_196;
input n_919;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_990;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_1058;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_293;
input n_1054;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_998;
input n_16;
input n_1046;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_962;
input n_1000;
input n_279;
input n_686;
input n_796;
input n_1041;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_984;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_1048;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_981;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_985;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_997;
input n_821;
input n_325;
input n_938;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_982;
input n_561;
input n_33;
input n_477;
input n_549;
input n_980;
input n_533;
input n_954;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_979;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_993;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_1051;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_1039;
input n_556;
input n_159;
input n_1034;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_560;
input n_1014;
input n_753;
input n_642;
input n_995;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_1053;
input n_530;
input n_277;
input n_520;
input n_1029;
input n_418;
input n_113;
input n_618;
input n_1055;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_1047;
input n_1010;
input n_355;
input n_426;
input n_317;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_1052;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_1006;
input n_373;
input n_1012;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_1045;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_1002;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_1019;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_983;
input n_64;
input n_288;
input n_427;
input n_1059;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_1001;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_1050;
input n_379;
input n_170;
input n_778;
input n_1025;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_1013;
input n_1023;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_1007;
input n_51;
input n_649;
input n_283;

output n_4803;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_4730;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_4598;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_4649;
wire n_1674;
wire n_1199;
wire n_3392;
wire n_4670;
wire n_3266;
wire n_1351;
wire n_3574;
wire n_4620;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_4738;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_4177;
wire n_3178;
wire n_1307;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1581;
wire n_4504;
wire n_3844;
wire n_4395;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4388;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_2451;
wire n_1620;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_2324;
wire n_1854;
wire n_1575;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_2260;
wire n_3222;
wire n_1387;
wire n_1708;
wire n_1151;
wire n_4686;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_4699;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_2557;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2405;
wire n_4050;
wire n_1743;
wire n_1160;
wire n_2647;
wire n_2997;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1238;
wire n_4092;
wire n_4645;
wire n_1724;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_4755;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_4578;
wire n_2211;
wire n_1415;
wire n_1555;
wire n_4777;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4591;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_4702;
wire n_2291;
wire n_4754;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_1285;
wire n_3946;
wire n_4213;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_4531;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_3626;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1532;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_2247;
wire n_1711;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_4666;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_4617;
wire n_4733;
wire n_2129;
wire n_2340;
wire n_4764;
wire n_1261;
wire n_4724;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_4555;
wire n_4743;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_2356;
wire n_1143;
wire n_1511;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_4696;
wire n_4692;
wire n_1572;
wire n_3979;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_2739;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_3023;
wire n_3890;
wire n_3232;
wire n_2791;
wire n_1313;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_4602;
wire n_2212;
wire n_3929;
wire n_3063;
wire n_3048;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1455;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_4767;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_4722;
wire n_4606;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_4187;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_2873;
wire n_1820;
wire n_1345;
wire n_3452;
wire n_3655;
wire n_4556;
wire n_3107;
wire n_4563;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_4687;
wire n_3948;
wire n_2836;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_4619;
wire n_2378;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_4600;
wire n_4125;
wire n_2625;
wire n_3296;
wire n_1400;
wire n_4646;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_4255;
wire n_4071;
wire n_4403;
wire n_4729;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1967;
wire n_1193;
wire n_3999;
wire n_3928;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_4751;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_4605;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_4549;
wire n_4575;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_1986;
wire n_4320;
wire n_4305;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_4102;
wire n_4297;
wire n_2113;
wire n_1641;
wire n_2190;
wire n_1918;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_4662;
wire n_1843;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_4314;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_3910;
wire n_1699;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_2633;
wire n_3883;
wire n_1848;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2059;
wire n_4507;
wire n_2198;
wire n_3319;
wire n_3728;
wire n_2669;
wire n_2925;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_4677;
wire n_3272;
wire n_4765;
wire n_3193;
wire n_2522;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_4732;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_1530;
wire n_3798;
wire n_3488;
wire n_2811;
wire n_1543;
wire n_3732;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_4372;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4581;
wire n_4226;
wire n_1762;
wire n_4641;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_4795;
wire n_3630;
wire n_4698;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_4792;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_2692;
wire n_3842;
wire n_1680;
wire n_3248;
wire n_2031;
wire n_4544;
wire n_2130;
wire n_1413;
wire n_1605;
wire n_1330;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_3092;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_1233;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_4742;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_2459;
wire n_1701;
wire n_1865;
wire n_3746;
wire n_1111;
wire n_2971;
wire n_1713;
wire n_4375;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_4526;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1950;
wire n_1726;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_4613;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_3012;
wire n_3772;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_4717;
wire n_3794;
wire n_3247;
wire n_3069;
wire n_3921;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1664;
wire n_1722;
wire n_4585;
wire n_4731;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_4773;
wire n_3933;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_2254;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_1747;
wire n_3691;
wire n_4427;
wire n_3861;
wire n_2624;
wire n_4066;
wire n_4386;
wire n_4485;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_4681;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_4523;
wire n_4752;
wire n_2347;
wire n_1214;
wire n_1886;
wire n_3917;
wire n_2092;
wire n_1654;
wire n_4371;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_4552;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_4673;
wire n_4313;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_4607;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_3873;
wire n_1624;
wire n_3983;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_4510;
wire n_1515;
wire n_4473;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_4169;
wire n_4055;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_3009;
wire n_1709;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_4589;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_2271;
wire n_3192;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4560;
wire n_4737;
wire n_4685;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_4675;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_2943;
wire n_1294;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_3253;
wire n_3337;
wire n_1779;
wire n_1465;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4002;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_3021;
wire n_1712;
wire n_4603;
wire n_1391;
wire n_4663;
wire n_2750;
wire n_2558;
wire n_1523;
wire n_2775;
wire n_2893;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_4697;
wire n_2954;
wire n_3477;
wire n_4289;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4288;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_3953;
wire n_1100;
wire n_4588;
wire n_4653;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_4802;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_4728;
wire n_4385;
wire n_1952;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_1932;
wire n_1101;
wire n_2535;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_4636;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_4701;
wire n_4651;
wire n_1451;
wire n_3941;
wire n_2767;
wire n_3793;
wire n_1839;
wire n_2341;
wire n_4576;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_4615;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_3293;
wire n_1646;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_4389;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_4661;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_2747;
wire n_1513;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_4621;
wire n_4216;
wire n_3608;
wire n_4540;
wire n_4315;
wire n_4664;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4240;
wire n_3491;
wire n_4156;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_2339;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3426;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_4785;
wire n_3470;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_4713;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_3700;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_4688;
wire n_3166;
wire n_4753;
wire n_2316;
wire n_1771;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_2239;
wire n_1707;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_4775;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_4674;
wire n_2717;
wire n_1723;
wire n_2191;
wire n_4481;
wire n_1246;
wire n_4528;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_4634;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_4123;
wire n_1431;
wire n_1615;
wire n_4114;
wire n_3312;
wire n_1474;
wire n_1571;
wire n_3835;
wire n_4587;
wire n_4286;
wire n_3119;
wire n_1809;
wire n_4280;
wire n_2958;
wire n_2948;
wire n_3735;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_4718;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_4525;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_2848;
wire n_1849;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4541;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4551;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_4459;
wire n_1299;
wire n_4545;
wire n_4708;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_4627;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_4624;
wire n_2837;
wire n_4175;
wire n_4700;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_4659;
wire n_4771;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_2127;
wire n_2338;
wire n_1178;
wire n_3324;
wire n_3593;
wire n_1424;
wire n_3341;
wire n_3867;
wire n_4455;
wire n_4453;
wire n_1073;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_4514;
wire n_3191;
wire n_1626;
wire n_4005;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_3546;
wire n_4798;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4564;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_2424;
wire n_2296;
wire n_1604;
wire n_3201;
wire n_1284;
wire n_3633;
wire n_3447;
wire n_4487;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1774;
wire n_3103;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_1201;
wire n_1398;
wire n_3638;
wire n_4592;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_3393;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_3451;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_1418;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_4695;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_4401;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_4796;
wire n_3606;
wire n_3142;
wire n_1310;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_3641;
wire n_1314;
wire n_2788;
wire n_2218;
wire n_1837;
wire n_4533;
wire n_4756;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_4419;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_1410;
wire n_4746;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1736;
wire n_1564;
wire n_4069;
wire n_4053;
wire n_2748;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_4658;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_2416;
wire n_1427;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_3909;
wire n_3944;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_4665;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_4633;
wire n_4654;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_4584;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3724;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_2990;
wire n_3847;
wire n_1775;
wire n_1286;
wire n_2115;
wire n_1773;
wire n_4430;
wire n_2410;
wire n_2552;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_1093;
wire n_4428;
wire n_4597;
wire n_1783;
wire n_3364;
wire n_2929;
wire n_3226;
wire n_2780;
wire n_3323;
wire n_1533;
wire n_1597;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_4404;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_4618;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4261;
wire n_4204;
wire n_1745;
wire n_4679;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_4015;
wire n_3547;
wire n_3869;
wire n_1901;
wire n_1374;
wire n_2556;
wire n_4706;
wire n_2648;
wire n_4747;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_4570;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_3188;
wire n_1459;
wire n_1614;
wire n_3742;
wire n_1892;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_2889;
wire n_1179;
wire n_3243;
wire n_3683;
wire n_4056;
wire n_1617;
wire n_4034;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_4622;
wire n_4721;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_2732;
wire n_4693;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_3284;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_2720;
wire n_1520;
wire n_3126;
wire n_2159;
wire n_2289;
wire n_2315;
wire n_1077;
wire n_1390;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_1419;
wire n_1733;
wire n_4132;
wire n_2995;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_3051;
wire n_1636;
wire n_1437;
wire n_4614;
wire n_4609;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_4707;
wire n_3367;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_4001;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_2627;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_4647;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4126;
wire n_2829;
wire n_3845;
wire n_1995;
wire n_2181;
wire n_3751;
wire n_1594;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_4632;
wire n_1429;
wire n_4655;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_4470;
wire n_3466;
wire n_4801;
wire n_3554;
wire n_1593;
wire n_4546;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_4583;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_2942;
wire n_1635;
wire n_4014;
wire n_1079;
wire n_4704;
wire n_4714;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_4509;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_4374;
wire n_2201;
wire n_3919;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_4668;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4635;
wire n_2984;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_3276;
wire n_2597;
wire n_2375;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_4582;
wire n_1728;
wire n_3973;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_3886;
wire n_2924;
wire n_4761;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_4420;
wire n_4710;
wire n_1510;
wire n_3637;
wire n_4574;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_2598;
wire n_1916;
wire n_1270;
wire n_2549;
wire n_4690;
wire n_1187;
wire n_4405;
wire n_4234;
wire n_4304;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_4558;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_4759;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_3634;
wire n_1847;
wire n_2302;
wire n_4211;
wire n_4667;
wire n_4182;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_4230;
wire n_4656;
wire n_1841;
wire n_4660;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4637;
wire n_4274;
wire n_2423;
wire n_3277;
wire n_4797;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_4270;
wire n_4189;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_2439;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_4155;
wire n_2740;
wire n_4238;
wire n_3011;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_4611;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_3042;
wire n_3213;
wire n_1589;
wire n_4333;
wire n_3820;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_4610;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1943;
wire n_1216;
wire n_3228;
wire n_3249;
wire n_2716;
wire n_1320;
wire n_3657;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_4725;
wire n_4590;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_3238;
wire n_3529;
wire n_2171;
wire n_1213;
wire n_1891;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_2392;
wire n_1272;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_4565;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_4567;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_4554;
wire n_3594;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_4586;
wire n_4778;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_2373;
wire n_1472;
wire n_2050;
wire n_4626;
wire n_4595;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_4734;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_3475;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_4680;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_3692;
wire n_4515;
wire n_4689;
wire n_4616;
wire n_2017;
wire n_1682;
wire n_4516;
wire n_2699;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_3029;
wire n_2200;
wire n_1828;
wire n_4258;
wire n_4547;
wire n_3597;
wire n_2760;
wire n_1940;
wire n_1979;
wire n_2560;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_4548;
wire n_4643;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_2376;
wire n_1405;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_4601;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_3681;
wire n_1569;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_4623;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_4553;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_4135;
wire n_4279;
wire n_2871;
wire n_4209;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_3858;
wire n_1845;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_3292;
wire n_1271;
wire n_1496;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_4644;
wire n_4790;
wire n_2258;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_4040;
wire n_4561;
wire n_4461;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_2390;
wire n_4007;
wire n_3712;
wire n_2310;
wire n_4608;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_4716;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_3381;
wire n_3562;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_4757;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_2195;
wire n_1633;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_3528;
wire n_2172;
wire n_4682;
wire n_3489;
wire n_4571;
wire n_4343;
wire n_2835;
wire n_4715;
wire n_4530;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_4694;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_4672;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_4604;
wire n_2939;
wire n_4782;
wire n_3305;
wire n_1906;
wire n_2992;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1672;
wire n_4185;
wire n_3221;
wire n_1758;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4407;
wire n_4378;
wire n_1914;
wire n_1318;
wire n_1475;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_4774;
wire n_2056;
wire n_4205;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_4524;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_4469;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_2083;
wire n_1931;
wire n_1269;
wire n_2834;
wire n_4572;
wire n_3207;
wire n_2668;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_4776;
wire n_1941;
wire n_3483;
wire n_1375;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_4726;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_1236;
wire n_1794;
wire n_2398;
wire n_1559;
wire n_1928;
wire n_1725;
wire n_3743;
wire n_1872;
wire n_3091;
wire n_4736;
wire n_4317;
wire n_4493;
wire n_4723;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_3124;
wire n_1741;
wire n_1325;
wire n_1746;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2923;
wire n_2793;
wire n_2715;
wire n_2885;
wire n_3711;
wire n_3776;
wire n_1804;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_4650;
wire n_4788;
wire n_2062;
wire n_4539;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_4421;
wire n_4719;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_4793;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1113;
wire n_2833;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_4799;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_4789;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_3621;
wire n_1476;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1800;
wire n_2241;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_4203;
wire n_3515;
wire n_1150;
wire n_3808;
wire n_3190;
wire n_1742;
wire n_4505;
wire n_4657;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1929;
wire n_1807;
wire n_2369;
wire n_1378;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_4542;
wire n_3199;
wire n_2931;
wire n_4462;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_4536;
wire n_4741;
wire n_4543;
wire n_3343;
wire n_3303;
wire n_4173;
wire n_2752;
wire n_4157;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4630;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_4550;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_2140;
wire n_4652;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_2358;
wire n_1401;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_4534;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_1132;
wire n_4748;
wire n_1074;
wire n_4439;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_4783;
wire n_3874;
wire n_2814;
wire n_2528;
wire n_1379;
wire n_4639;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_3027;
wire n_3231;
wire n_1554;
wire n_4083;
wire n_4494;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_4786;
wire n_4295;
wire n_1120;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_4579;
wire n_2020;
wire n_1643;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_4023;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_3583;
wire n_2883;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_2385;
wire n_1283;
wire n_4112;
wire n_4009;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_3268;
wire n_4027;
wire n_2149;
wire n_3057;
wire n_1754;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_2584;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_1994;
wire n_1812;
wire n_4557;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_4432;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_4593;
wire n_2906;
wire n_2769;
wire n_1303;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_4568;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1721;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_4569;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_4559;
wire n_1347;
wire n_4106;
wire n_3604;
wire n_1501;
wire n_1221;
wire n_3334;
wire n_4373;
wire n_1245;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_4711;
wire n_2952;
wire n_3068;
wire n_3853;
wire n_4740;
wire n_2117;
wire n_2234;
wire n_4631;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_3811;
wire n_4720;
wire n_3494;
wire n_1656;
wire n_1460;
wire n_2112;
wire n_2255;
wire n_2430;
wire n_3584;
wire n_1464;
wire n_1737;
wire n_3486;
wire n_1414;
wire n_4678;
wire n_4086;
wire n_2721;
wire n_2649;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_4068;
wire n_2032;
wire n_4625;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_4521;
wire n_2444;
wire n_2437;
wire n_1215;
wire n_2743;
wire n_3962;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_4766;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_4166;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_1253;
wire n_2242;
wire n_1266;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4744;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_3802;
wire n_1276;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1696;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_2609;
wire n_1161;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_4115;
wire n_2999;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_4265;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_4532;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4105;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_4244;
wire n_4486;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_4612;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_4353;
wire n_4104;
wire n_2531;
wire n_1789;
wire n_1770;
wire n_4787;
wire n_3285;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_4529;
wire n_3361;
wire n_3596;
wire n_3478;
wire n_4537;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4351;
wire n_4346;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_4316;
wire n_2723;
wire n_2440;
wire n_2233;
wire n_4779;
wire n_4640;
wire n_3521;
wire n_3233;
wire n_4599;
wire n_2800;
wire n_1710;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_2805;
wire n_1301;
wire n_4769;
wire n_3310;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_4628;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_4784;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_4508;
wire n_1763;
wire n_4594;
wire n_1998;
wire n_3066;
wire n_4727;
wire n_3101;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_1574;
wire n_3989;
wire n_2478;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_4108;
wire n_1133;
wire n_4460;
wire n_1194;
wire n_3374;
wire n_4538;
wire n_4506;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_4429;
wire n_2640;
wire n_3695;
wire n_4642;
wire n_4051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_4293;
wire n_3552;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_4684;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_4580;
wire n_3330;
wire n_1479;
wire n_4768;
wire n_2217;
wire n_2197;
wire n_1675;
wire n_4758;
wire n_4781;
wire n_2065;
wire n_2879;
wire n_3717;
wire n_4522;
wire n_4148;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_1629;
wire n_1170;
wire n_2221;
wire n_4263;
wire n_2055;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1861;
wire n_3110;
wire n_3017;
wire n_1632;
wire n_1890;
wire n_3955;
wire n_2477;
wire n_1805;
wire n_2280;
wire n_1888;
wire n_1557;
wire n_1833;
wire n_3903;
wire n_1311;
wire n_3945;
wire n_4780;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_1612;
wire n_2162;
wire n_3908;
wire n_2333;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_4750;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_4648;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_4129;
wire n_4457;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_4794;
wire n_4500;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1423;
wire n_1935;
wire n_4039;
wire n_4745;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4566;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_4275;
wire n_4482;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_1801;
wire n_4426;
wire n_2912;
wire n_4703;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_4762;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_4030;
wire n_3113;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_783),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_925),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_824),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_878),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_909),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_866),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_699),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_583),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_529),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_785),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_284),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_399),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_606),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_41),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_688),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_383),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_515),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_617),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_77),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_484),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_177),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_499),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_895),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_635),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_742),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_180),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_462),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_690),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_76),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_511),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_364),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_790),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_899),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_187),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_219),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_691),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1004),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_66),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_437),
.Y(n_1098)
);

CKINVDCx12_ASAP7_75t_R g1099 ( 
.A(n_269),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_210),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_63),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_790),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_890),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_627),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1032),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_488),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_539),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_351),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_884),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_604),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_529),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_631),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1027),
.Y(n_1113)
);

CKINVDCx14_ASAP7_75t_R g1114 ( 
.A(n_982),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_109),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1024),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_921),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_293),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_905),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_426),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_13),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_772),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_214),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_916),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_197),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_586),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_187),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_85),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_346),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_843),
.Y(n_1130)
);

CKINVDCx16_ASAP7_75t_R g1131 ( 
.A(n_266),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_523),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_310),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_858),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_874),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_587),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_357),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_50),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_92),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1044),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_377),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_936),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_921),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_908),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_877),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_197),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_959),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_693),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_167),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_823),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_945),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_5),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_545),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_501),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_920),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_818),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_199),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_704),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_784),
.Y(n_1159)
);

BUFx10_ASAP7_75t_L g1160 ( 
.A(n_203),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_328),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_507),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_164),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_387),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_40),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_542),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_615),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_847),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_10),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_825),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_867),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_468),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_287),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_566),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_665),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_39),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_650),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_803),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_884),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_802),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_56),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_208),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_815),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_806),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_54),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_560),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_137),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_844),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_938),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_235),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_466),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_432),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_413),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_396),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_112),
.Y(n_1195)
);

BUFx5_ASAP7_75t_L g1196 ( 
.A(n_484),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_176),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_928),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_602),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_172),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_542),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_337),
.Y(n_1202)
);

BUFx8_ASAP7_75t_SL g1203 ( 
.A(n_758),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_212),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_882),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_25),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_631),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_863),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_878),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_663),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_837),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_695),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_860),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_919),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_352),
.Y(n_1215)
);

BUFx10_ASAP7_75t_L g1216 ( 
.A(n_446),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_56),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_261),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_567),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_52),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_935),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_956),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_892),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_490),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_639),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_970),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_148),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_204),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1046),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_993),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_905),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_617),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_155),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_1007),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_527),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_21),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_12),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_877),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_85),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_663),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_855),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_499),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_694),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_120),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_21),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_452),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_119),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_557),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_781),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_565),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_959),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_789),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_568),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_386),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_417),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_729),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_704),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_118),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_132),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_188),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_830),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_392),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_705),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_270),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_979),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_931),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_132),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_561),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_629),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_870),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_324),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_690),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_960),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_290),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_310),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_772),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_164),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_459),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_44),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_403),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_943),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_573),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_983),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_148),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_448),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_909),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_28),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_699),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_630),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_823),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_309),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_879),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1033),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_123),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_578),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_429),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_998),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_953),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_837),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_177),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_514),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_710),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_702),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_390),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_3),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_376),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_983),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_646),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_721),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_228),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_354),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_974),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_586),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_730),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_376),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_652),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_8),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_639),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_479),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_182),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_788),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_913),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_693),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_970),
.Y(n_1324)
);

CKINVDCx16_ASAP7_75t_R g1325 ( 
.A(n_454),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_933),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_193),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_896),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_606),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_745),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_317),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_912),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_992),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_875),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_769),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_434),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_950),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_767),
.Y(n_1338)
);

INVxp33_ASAP7_75t_L g1339 ( 
.A(n_709),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_664),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_791),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_408),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_603),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_926),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_137),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_865),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_79),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1031),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_189),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_175),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_458),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_826),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_872),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_449),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_396),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_697),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_603),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_660),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_920),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_838),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_910),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_835),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_165),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_789),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_868),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_716),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_974),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1056),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_950),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_634),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_810),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_622),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_410),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_757),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_435),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_855),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_953),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_500),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_350),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_295),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_493),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_297),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_664),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_82),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_282),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_67),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_913),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_907),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_806),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_829),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_79),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_613),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_541),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_57),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_71),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_633),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_408),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_182),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_340),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_888),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_911),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_149),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_387),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_13),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_641),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_519),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_981),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_346),
.Y(n_1408)
);

BUFx10_ASAP7_75t_L g1409 ( 
.A(n_466),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_661),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_541),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_153),
.Y(n_1412)
);

CKINVDCx16_ASAP7_75t_R g1413 ( 
.A(n_963),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_412),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_486),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_42),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_166),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1015),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_258),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_715),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_18),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_115),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_70),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_733),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_733),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1040),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_917),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_436),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_260),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_567),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_29),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_731),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_843),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_881),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_500),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_903),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_948),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_384),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_507),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_849),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_129),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_276),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_766),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_834),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_734),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_816),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_879),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_373),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1017),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_779),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_230),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_568),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_939),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_398),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_381),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_956),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_326),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_780),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_334),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_781),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_342),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1058),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1043),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_420),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_778),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_398),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_694),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_154),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_846),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_454),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_23),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_900),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_273),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_521),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_771),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_701),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_95),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_391),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_707),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_805),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_120),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_426),
.Y(n_1482)
);

BUFx10_ASAP7_75t_L g1483 ( 
.A(n_477),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_181),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_611),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_151),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_278),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_626),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_873),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_436),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_751),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_531),
.Y(n_1492)
);

CKINVDCx16_ASAP7_75t_R g1493 ( 
.A(n_520),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_180),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_940),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_598),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_902),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_649),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_863),
.Y(n_1499)
);

CKINVDCx16_ASAP7_75t_R g1500 ( 
.A(n_677),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_944),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_54),
.Y(n_1502)
);

BUFx10_ASAP7_75t_L g1503 ( 
.A(n_36),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_692),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_749),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_922),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_758),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_797),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_688),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_288),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_839),
.Y(n_1511)
);

CKINVDCx16_ASAP7_75t_R g1512 ( 
.A(n_810),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_304),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_591),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_417),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_535),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_418),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_535),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_850),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_493),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_862),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_864),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_818),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_547),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_202),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_167),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_701),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1010),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_501),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_765),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_275),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_645),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_685),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1036),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_986),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_248),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_420),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_825),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_816),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_548),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_522),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_949),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_661),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_101),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_409),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_773),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_388),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_760),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1022),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_935),
.Y(n_1551)
);

BUFx10_ASAP7_75t_L g1552 ( 
.A(n_80),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_370),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_430),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_402),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_286),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_760),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_433),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_336),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_393),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_479),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_629),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_441),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_622),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_946),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_602),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_927),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_442),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_644),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_869),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_928),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1038),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_557),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_649),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_147),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_357),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_354),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_583),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_918),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1034),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_932),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_130),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_57),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_423),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_839),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_652),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1059),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_343),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_162),
.Y(n_1589)
);

BUFx10_ASAP7_75t_L g1590 ( 
.A(n_930),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_106),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_579),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_61),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_179),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_900),
.Y(n_1595)
);

CKINVDCx16_ASAP7_75t_R g1596 ( 
.A(n_250),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_695),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_856),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1009),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_889),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_817),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_522),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_979),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_41),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1003),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_285),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_351),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_675),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_898),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_467),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_569),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_822),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_697),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_290),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_582),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_227),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_457),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_198),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_978),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_238),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_121),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_859),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_957),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_34),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_116),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_40),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_747),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_319),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_166),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_740),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_952),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_419),
.Y(n_1632)
);

BUFx10_ASAP7_75t_L g1633 ( 
.A(n_718),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_997),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_907),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_526),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_709),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_885),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_914),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_212),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_836),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_35),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_591),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_289),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_419),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_764),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_513),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_100),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_63),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_580),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_359),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_876),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_506),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_518),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_641),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_604),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_538),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_273),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_315),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_394),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_195),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_300),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_613),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_343),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_761),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_725),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_223),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_457),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_819),
.Y(n_1669)
);

CKINVDCx16_ASAP7_75t_R g1670 ( 
.A(n_941),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_947),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_464),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_313),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_937),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_66),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_152),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_908),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_817),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_657),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_869),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_276),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_217),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_828),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_813),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_452),
.Y(n_1685)
);

CKINVDCx16_ASAP7_75t_R g1686 ( 
.A(n_339),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1054),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_362),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_355),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_852),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_453),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_241),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_576),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_881),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_686),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_280),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_293),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_209),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_456),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_918),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_851),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_753),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_483),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_646),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_880),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_811),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_845),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_708),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_584),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_893),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_608),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_477),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_307),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_845),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_515),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_476),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_20),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_546),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_264),
.Y(n_1719)
);

BUFx10_ASAP7_75t_L g1720 ( 
.A(n_889),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_931),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_906),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_307),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1014),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_317),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_942),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_562),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_871),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_894),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_73),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_848),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_723),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_392),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_136),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_98),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_680),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_914),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_20),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_37),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_463),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_934),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_549),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_842),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_304),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_104),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_800),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_219),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_692),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_55),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_556),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_486),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_388),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_990),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_430),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_947),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_460),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1008),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_734),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_51),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_871),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_851),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_17),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_517),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_924),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_558),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_98),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_632),
.Y(n_1767)
);

CKINVDCx20_ASAP7_75t_R g1768 ( 
.A(n_397),
.Y(n_1768)
);

BUFx10_ASAP7_75t_L g1769 ( 
.A(n_572),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_800),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_849),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_509),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_175),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_249),
.Y(n_1774)
);

BUFx3_ASAP7_75t_L g1775 ( 
.A(n_739),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_0),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1005),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_966),
.Y(n_1778)
);

CKINVDCx16_ASAP7_75t_R g1779 ( 
.A(n_87),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_550),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_445),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_833),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_333),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_861),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_774),
.Y(n_1785)
);

INVxp33_ASAP7_75t_SL g1786 ( 
.A(n_547),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_916),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1057),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_580),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_929),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_999),
.Y(n_1791)
);

CKINVDCx20_ASAP7_75t_R g1792 ( 
.A(n_227),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_283),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_517),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_300),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1039),
.Y(n_1796)
);

CKINVDCx16_ASAP7_75t_R g1797 ( 
.A(n_257),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_936),
.Y(n_1798)
);

CKINVDCx20_ASAP7_75t_R g1799 ( 
.A(n_798),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_298),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_147),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_369),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_157),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_892),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_127),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_961),
.Y(n_1807)
);

BUFx8_ASAP7_75t_SL g1808 ( 
.A(n_840),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_915),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_244),
.Y(n_1810)
);

CKINVDCx16_ASAP7_75t_R g1811 ( 
.A(n_316),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_904),
.Y(n_1812)
);

BUFx10_ASAP7_75t_L g1813 ( 
.A(n_505),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_901),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_404),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_654),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_162),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_886),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_558),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_207),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_819),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_490),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_794),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_84),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_841),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_78),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_360),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_755),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_844),
.Y(n_1829)
);

CKINVDCx16_ASAP7_75t_R g1830 ( 
.A(n_891),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_241),
.Y(n_1831)
);

INVxp33_ASAP7_75t_SL g1832 ( 
.A(n_721),
.Y(n_1832)
);

CKINVDCx20_ASAP7_75t_R g1833 ( 
.A(n_506),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_471),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_711),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_873),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_954),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_2),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_548),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_367),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1001),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_11),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_220),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_342),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_955),
.Y(n_1845)
);

BUFx10_ASAP7_75t_L g1846 ( 
.A(n_850),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_521),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_168),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_223),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_131),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_306),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_972),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_399),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_5),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_977),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_750),
.Y(n_1856)
);

CKINVDCx20_ASAP7_75t_R g1857 ( 
.A(n_689),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_279),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_221),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_23),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1053),
.Y(n_1861)
);

CKINVDCx20_ASAP7_75t_R g1862 ( 
.A(n_834),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_961),
.Y(n_1863)
);

CKINVDCx16_ASAP7_75t_R g1864 ( 
.A(n_411),
.Y(n_1864)
);

BUFx10_ASAP7_75t_L g1865 ( 
.A(n_226),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_47),
.Y(n_1866)
);

CKINVDCx20_ASAP7_75t_R g1867 ( 
.A(n_11),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_627),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_805),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_755),
.Y(n_1870)
);

CKINVDCx20_ASAP7_75t_R g1871 ( 
.A(n_857),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_943),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_666),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_468),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1025),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_45),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_962),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_880),
.Y(n_1878)
);

CKINVDCx20_ASAP7_75t_R g1879 ( 
.A(n_502),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_198),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1011),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_932),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_923),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_824),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_464),
.Y(n_1885)
);

CKINVDCx20_ASAP7_75t_R g1886 ( 
.A(n_713),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_958),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_544),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_554),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_713),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_968),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_367),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_401),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_883),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_72),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_887),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_113),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_854),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1021),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_788),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_383),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1028),
.Y(n_1902)
);

BUFx10_ASAP7_75t_L g1903 ( 
.A(n_205),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_298),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_600),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_971),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_67),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_853),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_365),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_897),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_658),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_972),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_199),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_554),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_951),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_827),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_352),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_43),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_596),
.Y(n_1919)
);

BUFx10_ASAP7_75t_L g1920 ( 
.A(n_667),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1196),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1196),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1116),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1203),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1099),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1196),
.Y(n_1926)
);

CKINVDCx14_ASAP7_75t_R g1927 ( 
.A(n_1114),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1196),
.Y(n_1928)
);

INVxp67_ASAP7_75t_SL g1929 ( 
.A(n_1229),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1196),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1203),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1196),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1196),
.Y(n_1933)
);

BUFx2_ASAP7_75t_SL g1934 ( 
.A(n_1116),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_1449),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1808),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1100),
.Y(n_1937)
);

CKINVDCx20_ASAP7_75t_R g1938 ( 
.A(n_1449),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1100),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1100),
.Y(n_1940)
);

INVx1_ASAP7_75t_SL g1941 ( 
.A(n_1153),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1529),
.Y(n_1942)
);

CKINVDCx16_ASAP7_75t_R g1943 ( 
.A(n_1117),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1529),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_1808),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1529),
.Y(n_1946)
);

INVxp67_ASAP7_75t_SL g1947 ( 
.A(n_1777),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1109),
.Y(n_1948)
);

INVxp33_ASAP7_75t_SL g1949 ( 
.A(n_1147),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1109),
.Y(n_1950)
);

CKINVDCx14_ASAP7_75t_R g1951 ( 
.A(n_1370),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1516),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1131),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1166),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1166),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1223),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1223),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1224),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1629),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1224),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1227),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1105),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1227),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1258),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1258),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_1230),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1259),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1259),
.Y(n_1968)
);

INVxp67_ASAP7_75t_SL g1969 ( 
.A(n_1411),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_1549),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1472),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1077),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1472),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1293),
.Y(n_1974)
);

INVxp67_ASAP7_75t_L g1975 ( 
.A(n_1734),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1333),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1348),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1481),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1481),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1491),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1491),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1525),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1525),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1535),
.Y(n_1984)
);

INVxp33_ASAP7_75t_SL g1985 ( 
.A(n_1460),
.Y(n_1985)
);

INVxp67_ASAP7_75t_SL g1986 ( 
.A(n_1603),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1535),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1568),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1568),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1077),
.Y(n_1990)
);

INVxp33_ASAP7_75t_SL g1991 ( 
.A(n_1630),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1609),
.Y(n_1992)
);

INVxp33_ASAP7_75t_L g1993 ( 
.A(n_1818),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1609),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1325),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1694),
.Y(n_1996)
);

INVxp33_ASAP7_75t_SL g1997 ( 
.A(n_1133),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1694),
.Y(n_1998)
);

CKINVDCx16_ASAP7_75t_R g1999 ( 
.A(n_1413),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1775),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1775),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1785),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1785),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1820),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1820),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1077),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1836),
.Y(n_2007)
);

CKINVDCx20_ASAP7_75t_R g2008 ( 
.A(n_1549),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1418),
.Y(n_2009)
);

INVxp67_ASAP7_75t_L g2010 ( 
.A(n_1920),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1836),
.Y(n_2011)
);

INVx1_ASAP7_75t_SL g2012 ( 
.A(n_1451),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1493),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1077),
.Y(n_2014)
);

INVxp67_ASAP7_75t_SL g2015 ( 
.A(n_1087),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1528),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1087),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1071),
.Y(n_2018)
);

CKINVDCx20_ASAP7_75t_R g2019 ( 
.A(n_1234),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1534),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1087),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1087),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1141),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1141),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1141),
.Y(n_2025)
);

INVxp67_ASAP7_75t_L g2026 ( 
.A(n_1920),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1572),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1141),
.Y(n_2028)
);

INVxp67_ASAP7_75t_SL g2029 ( 
.A(n_1144),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1144),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1144),
.Y(n_2031)
);

INVxp33_ASAP7_75t_SL g2032 ( 
.A(n_1133),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1144),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1219),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1219),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1219),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1219),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1580),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1261),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1261),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1261),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1261),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1634),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_1687),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1462),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1500),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1276),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_1753),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1276),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1757),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1276),
.Y(n_2051)
);

INVxp33_ASAP7_75t_SL g2052 ( 
.A(n_1134),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1276),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1289),
.Y(n_2054)
);

INVxp67_ASAP7_75t_SL g2055 ( 
.A(n_1289),
.Y(n_2055)
);

CKINVDCx16_ASAP7_75t_R g2056 ( 
.A(n_1512),
.Y(n_2056)
);

INVxp67_ASAP7_75t_SL g2057 ( 
.A(n_1289),
.Y(n_2057)
);

INVxp67_ASAP7_75t_SL g2058 ( 
.A(n_1289),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_1788),
.Y(n_2059)
);

INVxp33_ASAP7_75t_SL g2060 ( 
.A(n_1134),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_1861),
.Y(n_2061)
);

INVxp67_ASAP7_75t_L g2062 ( 
.A(n_1920),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1355),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1355),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1899),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1355),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1355),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1367),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1367),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1367),
.Y(n_2070)
);

CKINVDCx14_ASAP7_75t_R g2071 ( 
.A(n_1128),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1367),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1480),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1480),
.Y(n_2074)
);

INVxp33_ASAP7_75t_L g2075 ( 
.A(n_1339),
.Y(n_2075)
);

INVxp67_ASAP7_75t_L g2076 ( 
.A(n_1128),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1480),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_1902),
.Y(n_2078)
);

CKINVDCx20_ASAP7_75t_R g2079 ( 
.A(n_1587),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_1596),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1480),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1514),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_1587),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1514),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1670),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1514),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1514),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1518),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1518),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1518),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1518),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1686),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1540),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1540),
.Y(n_2094)
);

INVxp67_ASAP7_75t_SL g2095 ( 
.A(n_1540),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1540),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_1128),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1622),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1622),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1622),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1622),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1657),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1779),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1657),
.Y(n_2104)
);

CKINVDCx16_ASAP7_75t_R g2105 ( 
.A(n_1797),
.Y(n_2105)
);

INVxp67_ASAP7_75t_SL g2106 ( 
.A(n_1657),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1657),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1676),
.Y(n_2108)
);

INVxp67_ASAP7_75t_SL g2109 ( 
.A(n_1676),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1676),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1676),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1677),
.Y(n_2112)
);

INVxp33_ASAP7_75t_L g2113 ( 
.A(n_1073),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1677),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1677),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1677),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1462),
.Y(n_2117)
);

INVxp33_ASAP7_75t_SL g2118 ( 
.A(n_1136),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1972),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2015),
.Y(n_2120)
);

BUFx8_ASAP7_75t_L g2121 ( 
.A(n_1948),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2029),
.Y(n_2122)
);

OAI22xp5_ASAP7_75t_SL g2123 ( 
.A1(n_2019),
.A2(n_1081),
.B1(n_1093),
.B2(n_1072),
.Y(n_2123)
);

INVx6_ASAP7_75t_L g2124 ( 
.A(n_1943),
.Y(n_2124)
);

NAND2xp33_ASAP7_75t_L g2125 ( 
.A(n_2080),
.B(n_1136),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_SL g2126 ( 
.A1(n_1951),
.A2(n_1081),
.B1(n_1093),
.B2(n_1072),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1962),
.B(n_1841),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1990),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2055),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2006),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1966),
.B(n_1974),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_2061),
.B(n_1368),
.Y(n_2132)
);

AND2x6_ASAP7_75t_L g2133 ( 
.A(n_1921),
.B(n_1841),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2034),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2057),
.Y(n_2135)
);

OA21x2_ASAP7_75t_L g2136 ( 
.A1(n_1937),
.A2(n_1940),
.B(n_1939),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2035),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2037),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2053),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_2045),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_2045),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2058),
.Y(n_2142)
);

OAI21x1_ASAP7_75t_L g2143 ( 
.A1(n_1922),
.A2(n_1113),
.B(n_1096),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2095),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1950),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1927),
.B(n_1811),
.Y(n_2146)
);

OA21x2_ASAP7_75t_L g2147 ( 
.A1(n_1942),
.A2(n_1297),
.B(n_1140),
.Y(n_2147)
);

INVx4_ASAP7_75t_L g2148 ( 
.A(n_1976),
.Y(n_2148)
);

INVx3_ASAP7_75t_L g2149 ( 
.A(n_2102),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_2045),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2075),
.B(n_1830),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2106),
.Y(n_2152)
);

INVx5_ASAP7_75t_L g2153 ( 
.A(n_2117),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_1977),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2014),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_2117),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_2117),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_L g2158 ( 
.A(n_2085),
.Y(n_2158)
);

OA21x2_ASAP7_75t_L g2159 ( 
.A1(n_1944),
.A2(n_1946),
.B(n_1928),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2017),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_1947),
.B(n_1796),
.Y(n_2161)
);

OAI21x1_ASAP7_75t_L g2162 ( 
.A1(n_1926),
.A2(n_1463),
.B(n_1426),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2009),
.B(n_1599),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_2021),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2109),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2022),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2023),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2016),
.B(n_1605),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2024),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2025),
.Y(n_2170)
);

OAI21x1_ASAP7_75t_L g2171 ( 
.A1(n_1930),
.A2(n_1933),
.B(n_1932),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2028),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2030),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_2031),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_L g2175 ( 
.A(n_2033),
.Y(n_2175)
);

BUFx8_ASAP7_75t_L g2176 ( 
.A(n_1954),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2036),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2039),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_SL g2179 ( 
.A1(n_2079),
.A2(n_1121),
.B1(n_1124),
.B2(n_1118),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_2040),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2041),
.Y(n_2181)
);

AND2x6_ASAP7_75t_L g2182 ( 
.A(n_2042),
.B(n_1462),
.Y(n_2182)
);

INVxp67_ASAP7_75t_L g2183 ( 
.A(n_1953),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2047),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2049),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2051),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2054),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1929),
.B(n_1864),
.Y(n_2188)
);

INVx5_ASAP7_75t_L g2189 ( 
.A(n_1999),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2063),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2064),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_1949),
.A2(n_1832),
.B1(n_1786),
.B2(n_1061),
.Y(n_2192)
);

BUFx2_ASAP7_75t_L g2193 ( 
.A(n_2083),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_1969),
.B(n_1791),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2066),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_2067),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2068),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2069),
.Y(n_2198)
);

AOI22x1_ASAP7_75t_SL g2199 ( 
.A1(n_1923),
.A2(n_1121),
.B1(n_1124),
.B2(n_1118),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2070),
.Y(n_2200)
);

INVxp67_ASAP7_75t_L g2201 ( 
.A(n_1995),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2072),
.Y(n_2202)
);

BUFx3_ASAP7_75t_L g2203 ( 
.A(n_1955),
.Y(n_2203)
);

BUFx2_ASAP7_75t_L g2204 ( 
.A(n_2092),
.Y(n_2204)
);

OAI21x1_ASAP7_75t_L g2205 ( 
.A1(n_2073),
.A2(n_1127),
.B(n_1091),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2074),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2077),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2020),
.B(n_1881),
.Y(n_2208)
);

BUFx6f_ASAP7_75t_L g2209 ( 
.A(n_2081),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1985),
.A2(n_1832),
.B1(n_1786),
.B2(n_1062),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2082),
.Y(n_2211)
);

CKINVDCx20_ASAP7_75t_R g2212 ( 
.A(n_1935),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2084),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2071),
.B(n_1160),
.Y(n_2214)
);

INVxp67_ASAP7_75t_L g2215 ( 
.A(n_2013),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2018),
.B(n_1160),
.Y(n_2216)
);

INVx4_ASAP7_75t_L g2217 ( 
.A(n_2027),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2086),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_2087),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2038),
.B(n_1881),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2088),
.Y(n_2221)
);

BUFx6f_ASAP7_75t_L g2222 ( 
.A(n_2089),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2043),
.B(n_1462),
.Y(n_2223)
);

BUFx6f_ASAP7_75t_L g2224 ( 
.A(n_2090),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_1986),
.B(n_1185),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2091),
.Y(n_2226)
);

BUFx8_ASAP7_75t_L g2227 ( 
.A(n_1956),
.Y(n_2227)
);

BUFx2_ASAP7_75t_L g2228 ( 
.A(n_2103),
.Y(n_2228)
);

NAND2x1p5_ASAP7_75t_L g2229 ( 
.A(n_2018),
.B(n_1724),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2044),
.B(n_1160),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_2048),
.B(n_1185),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_2050),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2093),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2094),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2096),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2098),
.Y(n_2236)
);

INVx3_ASAP7_75t_L g2237 ( 
.A(n_2099),
.Y(n_2237)
);

INVx5_ASAP7_75t_L g2238 ( 
.A(n_2056),
.Y(n_2238)
);

BUFx6f_ASAP7_75t_L g2239 ( 
.A(n_2100),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2101),
.Y(n_2240)
);

BUFx12f_ASAP7_75t_L g2241 ( 
.A(n_1924),
.Y(n_2241)
);

INVx4_ASAP7_75t_L g2242 ( 
.A(n_2059),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2104),
.Y(n_2243)
);

BUFx3_ASAP7_75t_L g2244 ( 
.A(n_1957),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2107),
.Y(n_2245)
);

BUFx3_ASAP7_75t_L g2246 ( 
.A(n_1958),
.Y(n_2246)
);

NAND2x1p5_ASAP7_75t_L g2247 ( 
.A(n_2012),
.B(n_1724),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_2108),
.Y(n_2248)
);

BUFx8_ASAP7_75t_SL g2249 ( 
.A(n_1931),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_2065),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_1959),
.B(n_1189),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2110),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_SL g2253 ( 
.A(n_1952),
.B(n_1195),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2111),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_2078),
.B(n_1189),
.Y(n_2255)
);

BUFx12f_ASAP7_75t_L g2256 ( 
.A(n_1936),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_1975),
.B(n_1225),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2112),
.Y(n_2258)
);

INVxp67_ASAP7_75t_L g2259 ( 
.A(n_2046),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1960),
.B(n_1961),
.Y(n_2260)
);

BUFx8_ASAP7_75t_L g2261 ( 
.A(n_1963),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2114),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2115),
.Y(n_2263)
);

OAI22x1_ASAP7_75t_SL g2264 ( 
.A1(n_1991),
.A2(n_1200),
.B1(n_1210),
.B2(n_1195),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_1934),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2116),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_1945),
.Y(n_2267)
);

AOI22x1_ASAP7_75t_SL g2268 ( 
.A1(n_1938),
.A2(n_1210),
.B1(n_1255),
.B2(n_1200),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1964),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_1965),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2105),
.B(n_1163),
.Y(n_2271)
);

INVx3_ASAP7_75t_L g2272 ( 
.A(n_1967),
.Y(n_2272)
);

INVx3_ASAP7_75t_L g2273 ( 
.A(n_1968),
.Y(n_2273)
);

AND2x6_ASAP7_75t_L g2274 ( 
.A(n_1971),
.B(n_1724),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1973),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_1970),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1978),
.B(n_1724),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1979),
.B(n_1875),
.Y(n_2278)
);

OAI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_1941),
.A2(n_1296),
.B1(n_1538),
.B2(n_1292),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_1925),
.B(n_1225),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1980),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_1952),
.A2(n_1139),
.B1(n_1142),
.B2(n_1138),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1981),
.Y(n_2283)
);

INVx2_ASAP7_75t_SL g2284 ( 
.A(n_1982),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_1983),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1984),
.B(n_1875),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1987),
.B(n_1875),
.Y(n_2287)
);

INVx5_ASAP7_75t_L g2288 ( 
.A(n_1997),
.Y(n_2288)
);

INVx5_ASAP7_75t_L g2289 ( 
.A(n_2032),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1988),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_2010),
.Y(n_2291)
);

OA21x2_ASAP7_75t_L g2292 ( 
.A1(n_1989),
.A2(n_1127),
.B(n_1091),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_1992),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2026),
.B(n_1327),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1994),
.Y(n_2295)
);

OA21x2_ASAP7_75t_L g2296 ( 
.A1(n_1996),
.A2(n_1205),
.B(n_1162),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_2052),
.B(n_2060),
.Y(n_2297)
);

BUFx2_ASAP7_75t_L g2298 ( 
.A(n_2062),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_1998),
.B(n_1875),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2000),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2001),
.Y(n_2301)
);

INVx4_ASAP7_75t_L g2302 ( 
.A(n_2002),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2003),
.B(n_1327),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_2008),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2004),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2005),
.B(n_1357),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2007),
.B(n_2011),
.Y(n_2307)
);

INVx4_ASAP7_75t_L g2308 ( 
.A(n_2118),
.Y(n_2308)
);

OAI22xp5_ASAP7_75t_SL g2309 ( 
.A1(n_1993),
.A2(n_1262),
.B1(n_1290),
.B2(n_1255),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2113),
.Y(n_2310)
);

BUFx3_ASAP7_75t_L g2311 ( 
.A(n_2076),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2097),
.Y(n_2312)
);

AND2x4_ASAP7_75t_L g2313 ( 
.A(n_2061),
.B(n_1357),
.Y(n_2313)
);

AOI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_1949),
.A2(n_1063),
.B1(n_1064),
.B2(n_1060),
.Y(n_2314)
);

OA21x2_ASAP7_75t_L g2315 ( 
.A1(n_1937),
.A2(n_1205),
.B(n_1162),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_1972),
.Y(n_2316)
);

INVx3_ASAP7_75t_L g2317 ( 
.A(n_1972),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_1927),
.B(n_1163),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2015),
.Y(n_2319)
);

INVx5_ASAP7_75t_L g2320 ( 
.A(n_2045),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1962),
.B(n_1363),
.Y(n_2321)
);

AND2x4_ASAP7_75t_L g2322 ( 
.A(n_2061),
.B(n_1363),
.Y(n_2322)
);

BUFx6f_ASAP7_75t_L g2323 ( 
.A(n_2045),
.Y(n_2323)
);

OA21x2_ASAP7_75t_L g2324 ( 
.A1(n_1937),
.A2(n_1243),
.B(n_1231),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1972),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_L g2326 ( 
.A(n_2045),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1972),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2015),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2015),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1972),
.Y(n_2330)
);

AND2x4_ASAP7_75t_L g2331 ( 
.A(n_2061),
.B(n_1494),
.Y(n_2331)
);

OA21x2_ASAP7_75t_L g2332 ( 
.A1(n_1937),
.A2(n_1243),
.B(n_1231),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_1972),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1972),
.Y(n_2334)
);

OA21x2_ASAP7_75t_L g2335 ( 
.A1(n_1937),
.A2(n_1282),
.B(n_1280),
.Y(n_2335)
);

OAI21x1_ASAP7_75t_L g2336 ( 
.A1(n_1921),
.A2(n_1282),
.B(n_1280),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_1972),
.Y(n_2337)
);

OAI22x1_ASAP7_75t_R g2338 ( 
.A1(n_1923),
.A2(n_1290),
.B1(n_1322),
.B2(n_1262),
.Y(n_2338)
);

INVx3_ASAP7_75t_L g2339 ( 
.A(n_1972),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2015),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_1962),
.B(n_1494),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2015),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1972),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_1972),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_1972),
.Y(n_2345)
);

BUFx3_ASAP7_75t_L g2346 ( 
.A(n_2061),
.Y(n_2346)
);

BUFx12f_ASAP7_75t_L g2347 ( 
.A(n_1924),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2015),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2061),
.B(n_1595),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2015),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1962),
.B(n_1595),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_1972),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_2061),
.B(n_1666),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2015),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2015),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_2045),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2015),
.Y(n_2357)
);

AND2x4_ASAP7_75t_L g2358 ( 
.A(n_2061),
.B(n_1666),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_L g2359 ( 
.A(n_2045),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_2045),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2015),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1972),
.Y(n_2362)
);

BUFx6f_ASAP7_75t_L g2363 ( 
.A(n_2045),
.Y(n_2363)
);

OAI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_1949),
.A2(n_1139),
.B1(n_1142),
.B2(n_1138),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_1962),
.B(n_1683),
.Y(n_2365)
);

BUFx6f_ASAP7_75t_L g2366 ( 
.A(n_2045),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1962),
.B(n_1683),
.Y(n_2367)
);

OA21x2_ASAP7_75t_L g2368 ( 
.A1(n_1937),
.A2(n_1295),
.B(n_1288),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1972),
.Y(n_2369)
);

OAI21x1_ASAP7_75t_L g2370 ( 
.A1(n_1921),
.A2(n_1295),
.B(n_1288),
.Y(n_2370)
);

INVx5_ASAP7_75t_L g2371 ( 
.A(n_2045),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_L g2372 ( 
.A(n_2045),
.Y(n_2372)
);

BUFx12f_ASAP7_75t_L g2373 ( 
.A(n_1924),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_1972),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2015),
.Y(n_2375)
);

BUFx6f_ASAP7_75t_L g2376 ( 
.A(n_2045),
.Y(n_2376)
);

OAI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_1949),
.A2(n_1592),
.B1(n_1869),
.B2(n_1586),
.Y(n_2377)
);

CKINVDCx6p67_ASAP7_75t_R g2378 ( 
.A(n_1943),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_1962),
.B(n_1689),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_1962),
.B(n_1689),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_1972),
.Y(n_2381)
);

BUFx2_ASAP7_75t_L g2382 ( 
.A(n_2079),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_2080),
.Y(n_2383)
);

OAI21x1_ASAP7_75t_L g2384 ( 
.A1(n_1921),
.A2(n_1332),
.B(n_1300),
.Y(n_2384)
);

BUFx8_ASAP7_75t_SL g2385 ( 
.A(n_1924),
.Y(n_2385)
);

AOI22xp5_ASAP7_75t_L g2386 ( 
.A1(n_1949),
.A2(n_1066),
.B1(n_1067),
.B2(n_1065),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2061),
.B(n_1717),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_1972),
.Y(n_2388)
);

BUFx2_ASAP7_75t_L g2389 ( 
.A(n_2079),
.Y(n_2389)
);

INVx4_ASAP7_75t_L g2390 ( 
.A(n_1962),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2015),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_1972),
.Y(n_2392)
);

INVx6_ASAP7_75t_L g2393 ( 
.A(n_1943),
.Y(n_2393)
);

AOI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_1949),
.A2(n_1069),
.B1(n_1070),
.B2(n_1068),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_1972),
.Y(n_2395)
);

AND2x6_ASAP7_75t_L g2396 ( 
.A(n_1921),
.B(n_1300),
.Y(n_2396)
);

BUFx3_ASAP7_75t_L g2397 ( 
.A(n_2061),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_1962),
.Y(n_2398)
);

OA21x2_ASAP7_75t_L g2399 ( 
.A1(n_1937),
.A2(n_1356),
.B(n_1332),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2015),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_2045),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2015),
.Y(n_2402)
);

INVx3_ASAP7_75t_L g2403 ( 
.A(n_1972),
.Y(n_2403)
);

AND2x4_ASAP7_75t_L g2404 ( 
.A(n_2061),
.B(n_1717),
.Y(n_2404)
);

XNOR2x1_ASAP7_75t_L g2405 ( 
.A(n_1952),
.B(n_1586),
.Y(n_2405)
);

OAI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_1949),
.A2(n_1869),
.B1(n_1870),
.B2(n_1592),
.Y(n_2406)
);

OAI21x1_ASAP7_75t_L g2407 ( 
.A1(n_1921),
.A2(n_1364),
.B(n_1356),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_1972),
.Y(n_2408)
);

AND2x4_ASAP7_75t_L g2409 ( 
.A(n_2061),
.B(n_1760),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2015),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_1962),
.B(n_1760),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2015),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_1927),
.B(n_1163),
.Y(n_2413)
);

OAI22xp5_ASAP7_75t_SL g2414 ( 
.A1(n_2019),
.A2(n_1352),
.B1(n_1359),
.B2(n_1322),
.Y(n_2414)
);

INVx3_ASAP7_75t_L g2415 ( 
.A(n_1972),
.Y(n_2415)
);

INVx4_ASAP7_75t_L g2416 ( 
.A(n_1962),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2015),
.Y(n_2417)
);

HB1xp67_ASAP7_75t_L g2418 ( 
.A(n_2080),
.Y(n_2418)
);

INVx6_ASAP7_75t_L g2419 ( 
.A(n_1943),
.Y(n_2419)
);

INVx3_ASAP7_75t_L g2420 ( 
.A(n_1972),
.Y(n_2420)
);

BUFx6f_ASAP7_75t_L g2421 ( 
.A(n_2045),
.Y(n_2421)
);

INVx5_ASAP7_75t_L g2422 ( 
.A(n_2045),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_1972),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_2061),
.B(n_1793),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_1972),
.Y(n_2425)
);

AND2x4_ASAP7_75t_L g2426 ( 
.A(n_2061),
.B(n_1793),
.Y(n_2426)
);

OA21x2_ASAP7_75t_L g2427 ( 
.A1(n_1937),
.A2(n_1376),
.B(n_1364),
.Y(n_2427)
);

OAI21x1_ASAP7_75t_L g2428 ( 
.A1(n_1921),
.A2(n_1412),
.B(n_1376),
.Y(n_2428)
);

BUFx2_ASAP7_75t_L g2429 ( 
.A(n_2079),
.Y(n_2429)
);

BUFx8_ASAP7_75t_SL g2430 ( 
.A(n_1924),
.Y(n_2430)
);

CKINVDCx5p33_ASAP7_75t_R g2431 ( 
.A(n_1962),
.Y(n_2431)
);

AOI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_1949),
.A2(n_1075),
.B1(n_1076),
.B2(n_1074),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2015),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_1972),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_1972),
.Y(n_2435)
);

OA21x2_ASAP7_75t_L g2436 ( 
.A1(n_1937),
.A2(n_1422),
.B(n_1412),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_1972),
.Y(n_2437)
);

OAI22xp5_ASAP7_75t_SL g2438 ( 
.A1(n_2019),
.A2(n_1359),
.B1(n_1361),
.B2(n_1352),
.Y(n_2438)
);

CKINVDCx8_ASAP7_75t_R g2439 ( 
.A(n_1934),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2015),
.Y(n_2440)
);

OAI21x1_ASAP7_75t_L g2441 ( 
.A1(n_1921),
.A2(n_1425),
.B(n_1422),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2015),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_1949),
.A2(n_1872),
.B1(n_1873),
.B2(n_1870),
.Y(n_2443)
);

NAND2xp33_ASAP7_75t_L g2444 ( 
.A(n_2080),
.B(n_1872),
.Y(n_2444)
);

BUFx2_ASAP7_75t_L g2445 ( 
.A(n_2079),
.Y(n_2445)
);

AND2x4_ASAP7_75t_L g2446 ( 
.A(n_2061),
.B(n_1078),
.Y(n_2446)
);

OA21x2_ASAP7_75t_L g2447 ( 
.A1(n_1937),
.A2(n_1434),
.B(n_1425),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_1927),
.B(n_1216),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2015),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2015),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_1972),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_1972),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_1972),
.Y(n_2453)
);

INVx3_ASAP7_75t_L g2454 ( 
.A(n_1972),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2015),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_1962),
.B(n_1079),
.Y(n_2456)
);

INVx3_ASAP7_75t_L g2457 ( 
.A(n_1972),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_1962),
.B(n_1080),
.Y(n_2458)
);

OAI22xp5_ASAP7_75t_SL g2459 ( 
.A1(n_2019),
.A2(n_1369),
.B1(n_1386),
.B2(n_1361),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_1972),
.Y(n_2460)
);

CKINVDCx20_ASAP7_75t_R g2461 ( 
.A(n_2212),
.Y(n_2461)
);

CKINVDCx20_ASAP7_75t_R g2462 ( 
.A(n_2276),
.Y(n_2462)
);

NAND2xp33_ASAP7_75t_R g2463 ( 
.A(n_2298),
.B(n_1873),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_2216),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2164),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_2154),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_2232),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_2250),
.Y(n_2468)
);

CKINVDCx20_ASAP7_75t_R g2469 ( 
.A(n_2304),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2398),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_2140),
.Y(n_2471)
);

XNOR2xp5_ASAP7_75t_L g2472 ( 
.A(n_2126),
.B(n_1369),
.Y(n_2472)
);

CKINVDCx20_ASAP7_75t_R g2473 ( 
.A(n_2378),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2164),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2269),
.Y(n_2475)
);

NAND2xp33_ASAP7_75t_R g2476 ( 
.A(n_2204),
.B(n_2228),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2431),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_2265),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_2249),
.Y(n_2479)
);

CKINVDCx16_ASAP7_75t_R g2480 ( 
.A(n_2338),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2223),
.B(n_1434),
.Y(n_2481)
);

CKINVDCx5p33_ASAP7_75t_R g2482 ( 
.A(n_2385),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2174),
.Y(n_2483)
);

BUFx3_ASAP7_75t_L g2484 ( 
.A(n_2346),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2275),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2281),
.Y(n_2486)
);

CKINVDCx20_ASAP7_75t_R g2487 ( 
.A(n_2439),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2430),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2283),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_R g2490 ( 
.A(n_2267),
.B(n_1084),
.Y(n_2490)
);

NOR2x1p5_ASAP7_75t_L g2491 ( 
.A(n_2214),
.B(n_1874),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2290),
.Y(n_2492)
);

CKINVDCx20_ASAP7_75t_R g2493 ( 
.A(n_2193),
.Y(n_2493)
);

CKINVDCx20_ASAP7_75t_R g2494 ( 
.A(n_2382),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2241),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2127),
.B(n_1458),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_2256),
.Y(n_2497)
);

INVxp67_ASAP7_75t_L g2498 ( 
.A(n_2253),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2174),
.Y(n_2499)
);

CKINVDCx5p33_ASAP7_75t_R g2500 ( 
.A(n_2347),
.Y(n_2500)
);

BUFx2_ASAP7_75t_L g2501 ( 
.A(n_2151),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_2373),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2148),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2217),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_2242),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2175),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2140),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2300),
.Y(n_2508)
);

AND2x6_ASAP7_75t_L g2509 ( 
.A(n_2318),
.B(n_1458),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_2390),
.Y(n_2510)
);

INVxp67_ASAP7_75t_L g2511 ( 
.A(n_2310),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_2416),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2175),
.Y(n_2513)
);

OAI22xp5_ASAP7_75t_L g2514 ( 
.A1(n_2192),
.A2(n_1088),
.B1(n_1090),
.B2(n_1086),
.Y(n_2514)
);

AOI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2188),
.A2(n_1132),
.B1(n_1156),
.B2(n_1129),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2180),
.Y(n_2516)
);

OAI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_2210),
.A2(n_1181),
.B1(n_1217),
.B2(n_1169),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_R g2518 ( 
.A(n_2125),
.B(n_1092),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2305),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_2397),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_2389),
.Y(n_2521)
);

CKINVDCx20_ASAP7_75t_R g2522 ( 
.A(n_2429),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2270),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_2141),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_2445),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2131),
.Y(n_2526)
);

CKINVDCx5p33_ASAP7_75t_R g2527 ( 
.A(n_2189),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2270),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_L g2529 ( 
.A(n_2163),
.B(n_1097),
.Y(n_2529)
);

INVxp67_ASAP7_75t_SL g2530 ( 
.A(n_2141),
.Y(n_2530)
);

INVx3_ASAP7_75t_L g2531 ( 
.A(n_2150),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2189),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_2238),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2150),
.Y(n_2534)
);

OAI22xp33_ASAP7_75t_L g2535 ( 
.A1(n_2314),
.A2(n_1242),
.B1(n_1340),
.B2(n_1228),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_2238),
.Y(n_2536)
);

CKINVDCx20_ASAP7_75t_R g2537 ( 
.A(n_2124),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2285),
.Y(n_2538)
);

BUFx10_ASAP7_75t_L g2539 ( 
.A(n_2297),
.Y(n_2539)
);

CKINVDCx5p33_ASAP7_75t_R g2540 ( 
.A(n_2393),
.Y(n_2540)
);

CKINVDCx20_ASAP7_75t_R g2541 ( 
.A(n_2419),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_R g2542 ( 
.A(n_2444),
.B(n_1098),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_2288),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_2288),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_R g2545 ( 
.A(n_2120),
.B(n_1102),
.Y(n_2545)
);

CKINVDCx5p33_ASAP7_75t_R g2546 ( 
.A(n_2289),
.Y(n_2546)
);

INVx3_ASAP7_75t_L g2547 ( 
.A(n_2156),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2229),
.Y(n_2548)
);

NOR2xp67_ASAP7_75t_L g2549 ( 
.A(n_2289),
.B(n_991),
.Y(n_2549)
);

CKINVDCx20_ASAP7_75t_R g2550 ( 
.A(n_2158),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2285),
.Y(n_2551)
);

HB1xp67_ASAP7_75t_L g2552 ( 
.A(n_2247),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2293),
.Y(n_2553)
);

CKINVDCx20_ASAP7_75t_R g2554 ( 
.A(n_2383),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_2418),
.Y(n_2555)
);

CKINVDCx5p33_ASAP7_75t_R g2556 ( 
.A(n_2208),
.Y(n_2556)
);

CKINVDCx20_ASAP7_75t_R g2557 ( 
.A(n_2308),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_2220),
.Y(n_2558)
);

CKINVDCx11_ASAP7_75t_R g2559 ( 
.A(n_2311),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2180),
.Y(n_2560)
);

CKINVDCx20_ASAP7_75t_R g2561 ( 
.A(n_2456),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2146),
.B(n_1216),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2458),
.Y(n_2563)
);

BUFx10_ASAP7_75t_L g2564 ( 
.A(n_2231),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2413),
.B(n_1216),
.Y(n_2565)
);

CKINVDCx5p33_ASAP7_75t_R g2566 ( 
.A(n_2132),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2255),
.Y(n_2567)
);

AOI21x1_ASAP7_75t_L g2568 ( 
.A1(n_2168),
.A2(n_1083),
.B(n_1082),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2196),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2293),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_R g2571 ( 
.A(n_2122),
.B(n_1103),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2291),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2123),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_R g2574 ( 
.A(n_2129),
.B(n_1104),
.Y(n_2574)
);

INVx2_ASAP7_75t_SL g2575 ( 
.A(n_2230),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_2414),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2295),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2301),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2196),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_2438),
.Y(n_2580)
);

NAND2xp33_ASAP7_75t_R g2581 ( 
.A(n_2313),
.B(n_2322),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2145),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_L g2583 ( 
.A(n_2321),
.B(n_1106),
.Y(n_2583)
);

CKINVDCx20_ASAP7_75t_R g2584 ( 
.A(n_2459),
.Y(n_2584)
);

INVxp33_ASAP7_75t_L g2585 ( 
.A(n_2405),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2203),
.Y(n_2586)
);

NOR2xp33_ASAP7_75t_R g2587 ( 
.A(n_2135),
.B(n_1108),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_2179),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_R g2589 ( 
.A(n_2142),
.B(n_1110),
.Y(n_2589)
);

CKINVDCx20_ASAP7_75t_R g2590 ( 
.A(n_2183),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_2341),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2156),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2351),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_2365),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2367),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_R g2596 ( 
.A(n_2144),
.B(n_1111),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_R g2597 ( 
.A(n_2152),
.B(n_1112),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_R g2598 ( 
.A(n_2165),
.B(n_1120),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2379),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2244),
.Y(n_2600)
);

CKINVDCx20_ASAP7_75t_R g2601 ( 
.A(n_2201),
.Y(n_2601)
);

CKINVDCx5p33_ASAP7_75t_R g2602 ( 
.A(n_2380),
.Y(n_2602)
);

NAND2xp33_ASAP7_75t_R g2603 ( 
.A(n_2331),
.B(n_1874),
.Y(n_2603)
);

CKINVDCx5p33_ASAP7_75t_R g2604 ( 
.A(n_2411),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2319),
.B(n_1487),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_R g2606 ( 
.A(n_2328),
.B(n_2329),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2246),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2199),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_R g2609 ( 
.A(n_2340),
.B(n_1123),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_R g2610 ( 
.A(n_2342),
.B(n_1125),
.Y(n_2610)
);

INVx3_ASAP7_75t_L g2611 ( 
.A(n_2157),
.Y(n_2611)
);

BUFx10_ASAP7_75t_L g2612 ( 
.A(n_2251),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2348),
.Y(n_2613)
);

BUFx6f_ASAP7_75t_L g2614 ( 
.A(n_2157),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2268),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2209),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_R g2617 ( 
.A(n_2350),
.B(n_1126),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2209),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_2386),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_R g2620 ( 
.A(n_2354),
.B(n_1146),
.Y(n_2620)
);

NOR2xp67_ASAP7_75t_L g2621 ( 
.A(n_2215),
.B(n_994),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2355),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_2394),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2432),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2219),
.Y(n_2625)
);

BUFx3_ASAP7_75t_L g2626 ( 
.A(n_2136),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_2349),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_2353),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2358),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_2387),
.Y(n_2630)
);

CKINVDCx5p33_ASAP7_75t_R g2631 ( 
.A(n_2404),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_2409),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_2424),
.Y(n_2633)
);

HB1xp67_ASAP7_75t_L g2634 ( 
.A(n_2259),
.Y(n_2634)
);

CKINVDCx20_ASAP7_75t_R g2635 ( 
.A(n_2271),
.Y(n_2635)
);

CKINVDCx20_ASAP7_75t_R g2636 ( 
.A(n_2309),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2219),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2357),
.Y(n_2638)
);

INVx3_ASAP7_75t_L g2639 ( 
.A(n_2323),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2222),
.Y(n_2640)
);

CKINVDCx5p33_ASAP7_75t_R g2641 ( 
.A(n_2426),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_R g2642 ( 
.A(n_2361),
.B(n_1148),
.Y(n_2642)
);

AND3x2_ASAP7_75t_L g2643 ( 
.A(n_2448),
.B(n_1497),
.C(n_1487),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_2446),
.Y(n_2644)
);

INVx3_ASAP7_75t_L g2645 ( 
.A(n_2323),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_2312),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2326),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_2264),
.Y(n_2648)
);

HB1xp67_ASAP7_75t_L g2649 ( 
.A(n_2294),
.Y(n_2649)
);

CKINVDCx20_ASAP7_75t_R g2650 ( 
.A(n_2121),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2161),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2222),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_2364),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_2280),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_2377),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2375),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_2406),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_2443),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_2391),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2224),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2400),
.Y(n_2661)
);

CKINVDCx20_ASAP7_75t_R g2662 ( 
.A(n_2176),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2402),
.B(n_1497),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_R g2664 ( 
.A(n_2410),
.B(n_1151),
.Y(n_2664)
);

NAND2xp33_ASAP7_75t_R g2665 ( 
.A(n_2194),
.B(n_1877),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2412),
.Y(n_2666)
);

CKINVDCx5p33_ASAP7_75t_R g2667 ( 
.A(n_2417),
.Y(n_2667)
);

BUFx2_ASAP7_75t_SL g2668 ( 
.A(n_2284),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2433),
.B(n_1502),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_2440),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_2442),
.Y(n_2671)
);

INVx3_ASAP7_75t_L g2672 ( 
.A(n_2326),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_2449),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2450),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_R g2675 ( 
.A(n_2455),
.B(n_1152),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2224),
.Y(n_2676)
);

NOR2xp67_ASAP7_75t_L g2677 ( 
.A(n_2302),
.B(n_995),
.Y(n_2677)
);

CKINVDCx5p33_ASAP7_75t_R g2678 ( 
.A(n_2225),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2159),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2227),
.Y(n_2680)
);

CKINVDCx5p33_ASAP7_75t_R g2681 ( 
.A(n_2261),
.Y(n_2681)
);

BUFx2_ASAP7_75t_L g2682 ( 
.A(n_2257),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_2282),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2292),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2296),
.Y(n_2685)
);

BUFx6f_ASAP7_75t_L g2686 ( 
.A(n_2356),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2239),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2279),
.Y(n_2688)
);

CKINVDCx5p33_ASAP7_75t_R g2689 ( 
.A(n_2239),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_2263),
.Y(n_2690)
);

NAND2xp33_ASAP7_75t_R g2691 ( 
.A(n_2147),
.B(n_1877),
.Y(n_2691)
);

BUFx6f_ASAP7_75t_L g2692 ( 
.A(n_2356),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_2263),
.Y(n_2693)
);

CKINVDCx5p33_ASAP7_75t_R g2694 ( 
.A(n_2272),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_2273),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2260),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_2307),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2172),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2173),
.Y(n_2699)
);

NAND2xp33_ASAP7_75t_SL g2700 ( 
.A(n_2303),
.B(n_1386),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2119),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2306),
.Y(n_2702)
);

CKINVDCx20_ASAP7_75t_R g2703 ( 
.A(n_2277),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_2359),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2181),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2128),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_2359),
.Y(n_2707)
);

INVxp67_ASAP7_75t_SL g2708 ( 
.A(n_2360),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2187),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_2360),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_2363),
.Y(n_2711)
);

INVx1_ASAP7_75t_SL g2712 ( 
.A(n_2278),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_2363),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2130),
.Y(n_2714)
);

CKINVDCx5p33_ASAP7_75t_R g2715 ( 
.A(n_2366),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_2366),
.Y(n_2716)
);

INVx3_ASAP7_75t_L g2717 ( 
.A(n_2372),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2134),
.B(n_1502),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2137),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2149),
.B(n_2317),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2190),
.Y(n_2721)
);

HB1xp67_ASAP7_75t_L g2722 ( 
.A(n_2339),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2372),
.Y(n_2723)
);

INVx3_ASAP7_75t_L g2724 ( 
.A(n_2376),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_2376),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_2401),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2138),
.B(n_1561),
.Y(n_2727)
);

CKINVDCx20_ASAP7_75t_R g2728 ( 
.A(n_2286),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2401),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_2421),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_2421),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2139),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2352),
.B(n_1409),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2316),
.Y(n_2734)
);

INVx2_ASAP7_75t_SL g2735 ( 
.A(n_2388),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2325),
.Y(n_2736)
);

INVxp67_ASAP7_75t_L g2737 ( 
.A(n_2195),
.Y(n_2737)
);

CKINVDCx16_ASAP7_75t_R g2738 ( 
.A(n_2396),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_2327),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2330),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_2333),
.Y(n_2741)
);

HB1xp67_ASAP7_75t_L g2742 ( 
.A(n_2403),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_2334),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2197),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2206),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2337),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2226),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_2343),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2344),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2234),
.Y(n_2750)
);

CKINVDCx20_ASAP7_75t_R g2751 ( 
.A(n_2287),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2240),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_2345),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2243),
.Y(n_2754)
);

CKINVDCx20_ASAP7_75t_R g2755 ( 
.A(n_2299),
.Y(n_2755)
);

CKINVDCx5p33_ASAP7_75t_R g2756 ( 
.A(n_2362),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2369),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_2374),
.Y(n_2758)
);

INVx3_ASAP7_75t_L g2759 ( 
.A(n_2153),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_2381),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2392),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2395),
.Y(n_2762)
);

AND3x2_ASAP7_75t_L g2763 ( 
.A(n_2245),
.B(n_1571),
.C(n_1561),
.Y(n_2763)
);

BUFx3_ASAP7_75t_L g2764 ( 
.A(n_2315),
.Y(n_2764)
);

BUFx3_ASAP7_75t_L g2765 ( 
.A(n_2324),
.Y(n_2765)
);

CKINVDCx20_ASAP7_75t_R g2766 ( 
.A(n_2332),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2252),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2254),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2466),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2712),
.B(n_2396),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2701),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2706),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2475),
.Y(n_2773)
);

AO21x2_ASAP7_75t_L g2774 ( 
.A1(n_2684),
.A2(n_2143),
.B(n_2171),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2485),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2467),
.Y(n_2776)
);

BUFx6f_ASAP7_75t_L g2777 ( 
.A(n_2471),
.Y(n_2777)
);

BUFx6f_ASAP7_75t_L g2778 ( 
.A(n_2471),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2486),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2489),
.Y(n_2780)
);

AND2x6_ASAP7_75t_L g2781 ( 
.A(n_2685),
.B(n_1571),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2492),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2714),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2508),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2591),
.B(n_2153),
.Y(n_2785)
);

INVx4_ASAP7_75t_L g2786 ( 
.A(n_2689),
.Y(n_2786)
);

AO22x2_ASAP7_75t_L g2787 ( 
.A1(n_2514),
.A2(n_1362),
.B1(n_1365),
.B2(n_1343),
.Y(n_2787)
);

OR2x2_ASAP7_75t_L g2788 ( 
.A(n_2464),
.B(n_1432),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_2471),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2593),
.B(n_2320),
.Y(n_2790)
);

AOI22xp33_ASAP7_75t_L g2791 ( 
.A1(n_2626),
.A2(n_2396),
.B1(n_2133),
.B2(n_2428),
.Y(n_2791)
);

BUFx3_ASAP7_75t_L g2792 ( 
.A(n_2537),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2696),
.B(n_1409),
.Y(n_2793)
);

BUFx6f_ASAP7_75t_L g2794 ( 
.A(n_2614),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2519),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2722),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2567),
.B(n_2594),
.Y(n_2797)
);

NAND2x1p5_ASAP7_75t_L g2798 ( 
.A(n_2484),
.B(n_2428),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2563),
.B(n_2133),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2742),
.Y(n_2800)
);

INVx2_ASAP7_75t_SL g2801 ( 
.A(n_2612),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2698),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2699),
.Y(n_2803)
);

INVx5_ASAP7_75t_L g2804 ( 
.A(n_2612),
.Y(n_2804)
);

AND2x6_ASAP7_75t_L g2805 ( 
.A(n_2679),
.B(n_1604),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2705),
.Y(n_2806)
);

BUFx6f_ASAP7_75t_L g2807 ( 
.A(n_2614),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2719),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2709),
.Y(n_2809)
);

INVx8_ASAP7_75t_L g2810 ( 
.A(n_2541),
.Y(n_2810)
);

CKINVDCx20_ASAP7_75t_R g2811 ( 
.A(n_2461),
.Y(n_2811)
);

AND2x4_ASAP7_75t_L g2812 ( 
.A(n_2735),
.B(n_2266),
.Y(n_2812)
);

OR2x2_ASAP7_75t_L g2813 ( 
.A(n_2501),
.B(n_2682),
.Y(n_2813)
);

BUFx3_ASAP7_75t_L g2814 ( 
.A(n_2690),
.Y(n_2814)
);

NAND2x1p5_ASAP7_75t_L g2815 ( 
.A(n_2575),
.B(n_2335),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2697),
.B(n_1409),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2734),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2736),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2721),
.Y(n_2819)
);

INVx2_ASAP7_75t_SL g2820 ( 
.A(n_2733),
.Y(n_2820)
);

BUFx2_ASAP7_75t_L g2821 ( 
.A(n_2566),
.Y(n_2821)
);

AND2x6_ASAP7_75t_L g2822 ( 
.A(n_2565),
.B(n_1604),
.Y(n_2822)
);

BUFx3_ASAP7_75t_L g2823 ( 
.A(n_2693),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2744),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2745),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2762),
.Y(n_2826)
);

OR2x2_ASAP7_75t_L g2827 ( 
.A(n_2511),
.B(n_1707),
.Y(n_2827)
);

INVx3_ASAP7_75t_L g2828 ( 
.A(n_2614),
.Y(n_2828)
);

BUFx3_ASAP7_75t_L g2829 ( 
.A(n_2540),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2747),
.Y(n_2830)
);

INVx2_ASAP7_75t_SL g2831 ( 
.A(n_2678),
.Y(n_2831)
);

BUFx6f_ASAP7_75t_L g2832 ( 
.A(n_2686),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2750),
.Y(n_2833)
);

INVxp67_ASAP7_75t_L g2834 ( 
.A(n_2463),
.Y(n_2834)
);

BUFx4f_ASAP7_75t_L g2835 ( 
.A(n_2562),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2720),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2752),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2577),
.Y(n_2838)
);

INVxp67_ASAP7_75t_L g2839 ( 
.A(n_2603),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2754),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2767),
.Y(n_2841)
);

BUFx6f_ASAP7_75t_L g2842 ( 
.A(n_2686),
.Y(n_2842)
);

INVx6_ASAP7_75t_L g2843 ( 
.A(n_2539),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_SL g2844 ( 
.A(n_2595),
.B(n_2320),
.Y(n_2844)
);

NAND3xp33_ASAP7_75t_L g2845 ( 
.A(n_2529),
.B(n_1155),
.C(n_1154),
.Y(n_2845)
);

INVx4_ASAP7_75t_L g2846 ( 
.A(n_2704),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2768),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2578),
.Y(n_2848)
);

INVx3_ASAP7_75t_L g2849 ( 
.A(n_2686),
.Y(n_2849)
);

INVx4_ASAP7_75t_L g2850 ( 
.A(n_2707),
.Y(n_2850)
);

BUFx3_ASAP7_75t_L g2851 ( 
.A(n_2710),
.Y(n_2851)
);

BUFx6f_ASAP7_75t_L g2852 ( 
.A(n_2692),
.Y(n_2852)
);

BUFx6f_ASAP7_75t_L g2853 ( 
.A(n_2692),
.Y(n_2853)
);

INVx6_ASAP7_75t_L g2854 ( 
.A(n_2539),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2613),
.Y(n_2855)
);

NAND2x1p5_ASAP7_75t_L g2856 ( 
.A(n_2549),
.B(n_2368),
.Y(n_2856)
);

AND2x4_ASAP7_75t_L g2857 ( 
.A(n_2523),
.B(n_2423),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_SL g2858 ( 
.A(n_2599),
.B(n_2602),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2764),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2556),
.B(n_2133),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2558),
.B(n_2399),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2622),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2765),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2638),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2656),
.Y(n_2865)
);

BUFx3_ASAP7_75t_L g2866 ( 
.A(n_2711),
.Y(n_2866)
);

INVx4_ASAP7_75t_L g2867 ( 
.A(n_2713),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2661),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2666),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_SL g2870 ( 
.A(n_2604),
.B(n_2371),
.Y(n_2870)
);

AND2x2_ASAP7_75t_SL g2871 ( 
.A(n_2480),
.B(n_1610),
.Y(n_2871)
);

HB1xp67_ASAP7_75t_L g2872 ( 
.A(n_2581),
.Y(n_2872)
);

NAND3xp33_ASAP7_75t_L g2873 ( 
.A(n_2583),
.B(n_2667),
.C(n_2659),
.Y(n_2873)
);

BUFx2_ASAP7_75t_L g2874 ( 
.A(n_2590),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2526),
.B(n_2427),
.Y(n_2875)
);

NOR2xp33_ASAP7_75t_L g2876 ( 
.A(n_2702),
.B(n_1723),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2674),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2718),
.Y(n_2878)
);

NAND3xp33_ASAP7_75t_L g2879 ( 
.A(n_2670),
.B(n_1159),
.C(n_1157),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2481),
.B(n_2436),
.Y(n_2880)
);

CKINVDCx11_ASAP7_75t_R g2881 ( 
.A(n_2473),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_SL g2882 ( 
.A(n_2671),
.B(n_2371),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2673),
.B(n_1735),
.Y(n_2883)
);

BUFx2_ASAP7_75t_L g2884 ( 
.A(n_2601),
.Y(n_2884)
);

INVx4_ASAP7_75t_SL g2885 ( 
.A(n_2509),
.Y(n_2885)
);

INVxp67_ASAP7_75t_SL g2886 ( 
.A(n_2692),
.Y(n_2886)
);

AND2x6_ASAP7_75t_L g2887 ( 
.A(n_2496),
.B(n_1610),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2646),
.B(n_1736),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2766),
.A2(n_2370),
.B1(n_2384),
.B2(n_2336),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2727),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2738),
.B(n_2422),
.Y(n_2891)
);

AND2x4_ASAP7_75t_L g2892 ( 
.A(n_2528),
.B(n_2425),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_SL g2893 ( 
.A(n_2694),
.B(n_2422),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2509),
.B(n_2447),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2509),
.B(n_2434),
.Y(n_2895)
);

BUFx3_ASAP7_75t_L g2896 ( 
.A(n_2715),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2732),
.Y(n_2897)
);

AND2x2_ASAP7_75t_L g2898 ( 
.A(n_2668),
.B(n_1483),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2739),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2740),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2564),
.B(n_1762),
.Y(n_2901)
);

NOR3xp33_ASAP7_75t_L g2902 ( 
.A(n_2535),
.B(n_1780),
.C(n_1772),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2465),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2741),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_SL g2905 ( 
.A(n_2695),
.B(n_2155),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2509),
.B(n_2435),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2654),
.B(n_1483),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_L g2908 ( 
.A(n_2559),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2743),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2746),
.B(n_2437),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2748),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2749),
.Y(n_2912)
);

OAI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2651),
.A2(n_1878),
.B1(n_1883),
.B2(n_1807),
.Y(n_2913)
);

AND2x4_ASAP7_75t_L g2914 ( 
.A(n_2538),
.B(n_2451),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2753),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2474),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2756),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2564),
.B(n_2627),
.Y(n_2918)
);

BUFx3_ASAP7_75t_L g2919 ( 
.A(n_2716),
.Y(n_2919)
);

AND2x6_ASAP7_75t_L g2920 ( 
.A(n_2582),
.B(n_1727),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2483),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2634),
.B(n_1910),
.Y(n_2922)
);

AO22x1_ASAP7_75t_L g2923 ( 
.A1(n_2683),
.A2(n_1882),
.B1(n_1089),
.B2(n_1094),
.Y(n_2923)
);

INVx3_ASAP7_75t_L g2924 ( 
.A(n_2507),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2757),
.Y(n_2925)
);

BUFx6f_ASAP7_75t_L g2926 ( 
.A(n_2723),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2758),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2760),
.B(n_2452),
.Y(n_2928)
);

CKINVDCx20_ASAP7_75t_R g2929 ( 
.A(n_2462),
.Y(n_2929)
);

AND2x4_ASAP7_75t_L g2930 ( 
.A(n_2551),
.B(n_2453),
.Y(n_2930)
);

INVx3_ASAP7_75t_L g2931 ( 
.A(n_2507),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2649),
.B(n_1483),
.Y(n_2932)
);

NOR2xp33_ASAP7_75t_L g2933 ( 
.A(n_2703),
.B(n_1164),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2628),
.B(n_1503),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2629),
.B(n_1503),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2761),
.Y(n_2936)
);

AND2x6_ASAP7_75t_L g2937 ( 
.A(n_2586),
.B(n_1727),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2499),
.Y(n_2938)
);

NOR2xp33_ASAP7_75t_L g2939 ( 
.A(n_2728),
.B(n_1165),
.Y(n_2939)
);

AND2x6_ASAP7_75t_L g2940 ( 
.A(n_2600),
.B(n_1750),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2605),
.Y(n_2941)
);

INVxp67_ASAP7_75t_L g2942 ( 
.A(n_2665),
.Y(n_2942)
);

AND2x2_ASAP7_75t_L g2943 ( 
.A(n_2630),
.B(n_1503),
.Y(n_2943)
);

INVx4_ASAP7_75t_L g2944 ( 
.A(n_2725),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2663),
.Y(n_2945)
);

NAND2xp33_ASAP7_75t_L g2946 ( 
.A(n_2518),
.B(n_2274),
.Y(n_2946)
);

BUFx2_ASAP7_75t_L g2947 ( 
.A(n_2493),
.Y(n_2947)
);

BUFx6f_ASAP7_75t_L g2948 ( 
.A(n_2726),
.Y(n_2948)
);

BUFx2_ASAP7_75t_L g2949 ( 
.A(n_2494),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_SL g2950 ( 
.A(n_2631),
.B(n_2160),
.Y(n_2950)
);

BUFx3_ASAP7_75t_L g2951 ( 
.A(n_2729),
.Y(n_2951)
);

AND2x4_ASAP7_75t_L g2952 ( 
.A(n_2553),
.B(n_2460),
.Y(n_2952)
);

OR2x2_ASAP7_75t_L g2953 ( 
.A(n_2498),
.B(n_1882),
.Y(n_2953)
);

NOR2xp33_ASAP7_75t_L g2954 ( 
.A(n_2751),
.B(n_1167),
.Y(n_2954)
);

INVxp33_ASAP7_75t_L g2955 ( 
.A(n_2490),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2669),
.Y(n_2956)
);

INVx3_ASAP7_75t_L g2957 ( 
.A(n_2524),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2737),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_L g2959 ( 
.A(n_2755),
.B(n_1168),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2607),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2506),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2513),
.Y(n_2962)
);

HB1xp67_ASAP7_75t_L g2963 ( 
.A(n_2632),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2570),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2524),
.Y(n_2965)
);

INVx4_ASAP7_75t_L g2966 ( 
.A(n_2730),
.Y(n_2966)
);

INVx4_ASAP7_75t_L g2967 ( 
.A(n_2731),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2633),
.B(n_1552),
.Y(n_2968)
);

INVx4_ASAP7_75t_L g2969 ( 
.A(n_2520),
.Y(n_2969)
);

AND2x4_ASAP7_75t_L g2970 ( 
.A(n_2516),
.B(n_2408),
.Y(n_2970)
);

AND2x6_ASAP7_75t_L g2971 ( 
.A(n_2515),
.B(n_1750),
.Y(n_2971)
);

BUFx6f_ASAP7_75t_L g2972 ( 
.A(n_2531),
.Y(n_2972)
);

INVx4_ASAP7_75t_L g2973 ( 
.A(n_2527),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2560),
.Y(n_2974)
);

CKINVDCx5p33_ASAP7_75t_R g2975 ( 
.A(n_2468),
.Y(n_2975)
);

INVx2_ASAP7_75t_SL g2976 ( 
.A(n_2641),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2548),
.B(n_1552),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2478),
.B(n_2552),
.Y(n_2978)
);

INVx4_ASAP7_75t_L g2979 ( 
.A(n_2532),
.Y(n_2979)
);

INVx8_ASAP7_75t_L g2980 ( 
.A(n_2469),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2531),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2606),
.B(n_2143),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2534),
.Y(n_2983)
);

AND2x6_ASAP7_75t_L g2984 ( 
.A(n_2569),
.B(n_1766),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2503),
.B(n_2504),
.Y(n_2985)
);

INVxp67_ASAP7_75t_L g2986 ( 
.A(n_2476),
.Y(n_2986)
);

INVx2_ASAP7_75t_SL g2987 ( 
.A(n_2643),
.Y(n_2987)
);

AND2x6_ASAP7_75t_L g2988 ( 
.A(n_2579),
.B(n_1766),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2505),
.B(n_2166),
.Y(n_2989)
);

INVx3_ASAP7_75t_L g2990 ( 
.A(n_2534),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2547),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2572),
.B(n_1552),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2510),
.B(n_2167),
.Y(n_2993)
);

CKINVDCx5p33_ASAP7_75t_R g2994 ( 
.A(n_2470),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2619),
.B(n_1170),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2555),
.B(n_1590),
.Y(n_2996)
);

BUFx6f_ASAP7_75t_L g2997 ( 
.A(n_2547),
.Y(n_2997)
);

INVx3_ASAP7_75t_L g2998 ( 
.A(n_2592),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2592),
.Y(n_2999)
);

INVx1_ASAP7_75t_SL g3000 ( 
.A(n_2522),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2611),
.Y(n_3001)
);

BUFx3_ASAP7_75t_L g3002 ( 
.A(n_2487),
.Y(n_3002)
);

INVx4_ASAP7_75t_L g3003 ( 
.A(n_2533),
.Y(n_3003)
);

INVx2_ASAP7_75t_SL g3004 ( 
.A(n_2611),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2639),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2616),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2639),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2645),
.Y(n_3008)
);

BUFx3_ASAP7_75t_L g3009 ( 
.A(n_2645),
.Y(n_3009)
);

AOI22xp5_ASAP7_75t_L g3010 ( 
.A1(n_2561),
.A2(n_2274),
.B1(n_2169),
.B2(n_2177),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2647),
.Y(n_3011)
);

INVx3_ASAP7_75t_L g3012 ( 
.A(n_2647),
.Y(n_3012)
);

OAI221xp5_ASAP7_75t_L g3013 ( 
.A1(n_2691),
.A2(n_1101),
.B1(n_1107),
.B2(n_1095),
.C(n_1085),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2672),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2672),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2618),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2941),
.B(n_2512),
.Y(n_3017)
);

INVx2_ASAP7_75t_SL g3018 ( 
.A(n_2813),
.Y(n_3018)
);

AND2x2_ASAP7_75t_L g3019 ( 
.A(n_2876),
.B(n_2477),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_2797),
.B(n_2585),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2859),
.Y(n_3021)
);

INVx2_ASAP7_75t_SL g3022 ( 
.A(n_2898),
.Y(n_3022)
);

OAI221xp5_ASAP7_75t_L g3023 ( 
.A1(n_3013),
.A2(n_2700),
.B1(n_2624),
.B2(n_2623),
.C(n_2688),
.Y(n_3023)
);

NOR2xp67_ASAP7_75t_SL g3024 ( 
.A(n_2926),
.B(n_2536),
.Y(n_3024)
);

INVxp67_ASAP7_75t_SL g3025 ( 
.A(n_2863),
.Y(n_3025)
);

CKINVDCx5p33_ASAP7_75t_R g3026 ( 
.A(n_2769),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2873),
.B(n_2542),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2945),
.B(n_2956),
.Y(n_3028)
);

AOI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2942),
.A2(n_2839),
.B1(n_2890),
.B2(n_2878),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2836),
.Y(n_3030)
);

AND2x6_ASAP7_75t_SL g3031 ( 
.A(n_2995),
.B(n_2933),
.Y(n_3031)
);

BUFx2_ASAP7_75t_L g3032 ( 
.A(n_2947),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2855),
.B(n_2621),
.Y(n_3033)
);

NOR2xp33_ASAP7_75t_L g3034 ( 
.A(n_2883),
.B(n_2653),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2862),
.B(n_2545),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2864),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_SL g3037 ( 
.A(n_2835),
.B(n_2644),
.Y(n_3037)
);

AOI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_2880),
.A2(n_2637),
.B(n_2625),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2888),
.B(n_2491),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_2793),
.B(n_2521),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2868),
.Y(n_3041)
);

NOR2xp33_ASAP7_75t_L g3042 ( 
.A(n_2834),
.B(n_2655),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2773),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2771),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2865),
.B(n_2571),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2775),
.Y(n_3046)
);

NOR3xp33_ASAP7_75t_L g3047 ( 
.A(n_2858),
.B(n_2517),
.C(n_2525),
.Y(n_3047)
);

NOR2x1p5_ASAP7_75t_L g3048 ( 
.A(n_2814),
.B(n_2479),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_SL g3049 ( 
.A(n_2820),
.B(n_2574),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2772),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_SL g3051 ( 
.A1(n_2816),
.A2(n_2588),
.B1(n_2576),
.B2(n_2580),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_SL g3052 ( 
.A(n_2872),
.B(n_2587),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2922),
.B(n_2589),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2869),
.B(n_2596),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2986),
.B(n_2597),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2877),
.B(n_2598),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2779),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_SL g3058 ( 
.A(n_2770),
.B(n_2609),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2861),
.B(n_2610),
.Y(n_3059)
);

NOR3xp33_ASAP7_75t_L g3060 ( 
.A(n_2939),
.B(n_2573),
.C(n_2657),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2780),
.Y(n_3061)
);

NOR2xp33_ASAP7_75t_L g3062 ( 
.A(n_2901),
.B(n_2955),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_SL g3063 ( 
.A(n_2860),
.B(n_2617),
.Y(n_3063)
);

OR2x2_ASAP7_75t_L g3064 ( 
.A(n_2827),
.B(n_2658),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2782),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2875),
.B(n_2620),
.Y(n_3066)
);

AOI22xp33_ASAP7_75t_SL g3067 ( 
.A1(n_2822),
.A2(n_2635),
.B1(n_2636),
.B2(n_2584),
.Y(n_3067)
);

BUFx6f_ASAP7_75t_SL g3068 ( 
.A(n_2908),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2784),
.B(n_2642),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2795),
.B(n_2664),
.Y(n_3070)
);

AOI22xp5_ASAP7_75t_L g3071 ( 
.A1(n_2822),
.A2(n_2557),
.B1(n_2677),
.B2(n_2554),
.Y(n_3071)
);

OAI221xp5_ASAP7_75t_L g3072 ( 
.A1(n_2902),
.A2(n_2472),
.B1(n_1122),
.B2(n_1130),
.C(n_1119),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2783),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2897),
.B(n_2675),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2899),
.B(n_2543),
.Y(n_3075)
);

NOR2xp67_ASAP7_75t_L g3076 ( 
.A(n_2985),
.B(n_2495),
.Y(n_3076)
);

INVx2_ASAP7_75t_SL g3077 ( 
.A(n_2823),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2808),
.Y(n_3078)
);

CKINVDCx5p33_ASAP7_75t_R g3079 ( 
.A(n_2776),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2900),
.B(n_2544),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2802),
.B(n_2530),
.Y(n_3081)
);

CKINVDCx5p33_ASAP7_75t_R g3082 ( 
.A(n_2975),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2803),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2817),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2806),
.B(n_2708),
.Y(n_3085)
);

NAND3xp33_ASAP7_75t_L g3086 ( 
.A(n_2954),
.B(n_2546),
.C(n_2687),
.Y(n_3086)
);

AOI22xp5_ASAP7_75t_L g3087 ( 
.A1(n_2822),
.A2(n_2550),
.B1(n_2652),
.B2(n_2640),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2809),
.Y(n_3088)
);

OAI22xp5_ASAP7_75t_L g3089 ( 
.A1(n_2791),
.A2(n_2568),
.B1(n_1421),
.B2(n_1441),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2819),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2818),
.Y(n_3091)
);

NAND2xp33_ASAP7_75t_L g3092 ( 
.A(n_2805),
.B(n_2660),
.Y(n_3092)
);

NOR3xp33_ASAP7_75t_L g3093 ( 
.A(n_2959),
.B(n_2648),
.C(n_2615),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_2904),
.B(n_2717),
.Y(n_3094)
);

INVx3_ASAP7_75t_L g3095 ( 
.A(n_2798),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2824),
.B(n_2825),
.Y(n_3096)
);

AND2x2_ASAP7_75t_L g3097 ( 
.A(n_2996),
.B(n_2676),
.Y(n_3097)
);

BUFx8_ASAP7_75t_L g3098 ( 
.A(n_2908),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2830),
.Y(n_3099)
);

BUFx6f_ASAP7_75t_SL g3100 ( 
.A(n_2829),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2833),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2837),
.B(n_2717),
.Y(n_3102)
);

HB1xp67_ASAP7_75t_L g3103 ( 
.A(n_2926),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2840),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2841),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_L g3106 ( 
.A(n_2909),
.B(n_2724),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2847),
.Y(n_3107)
);

NOR2xp33_ASAP7_75t_L g3108 ( 
.A(n_2911),
.B(n_2724),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2799),
.B(n_2170),
.Y(n_3109)
);

INVxp67_ASAP7_75t_L g3110 ( 
.A(n_2788),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2958),
.B(n_2178),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2826),
.B(n_2781),
.Y(n_3112)
);

NOR2xp67_ASAP7_75t_L g3113 ( 
.A(n_2786),
.B(n_2497),
.Y(n_3113)
);

INVx1_ASAP7_75t_SL g3114 ( 
.A(n_3000),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2781),
.B(n_2184),
.Y(n_3115)
);

INVx2_ASAP7_75t_SL g3116 ( 
.A(n_2977),
.Y(n_3116)
);

AOI22xp33_ASAP7_75t_L g3117 ( 
.A1(n_2971),
.A2(n_2407),
.B1(n_2441),
.B2(n_2205),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2781),
.B(n_2185),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2838),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2989),
.B(n_2186),
.Y(n_3120)
);

BUFx5_ASAP7_75t_L g3121 ( 
.A(n_2805),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2993),
.B(n_2191),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2910),
.B(n_2198),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_SL g3124 ( 
.A(n_2994),
.B(n_2482),
.Y(n_3124)
);

INVx2_ASAP7_75t_SL g3125 ( 
.A(n_2948),
.Y(n_3125)
);

AOI22xp33_ASAP7_75t_L g3126 ( 
.A1(n_2971),
.A2(n_1421),
.B1(n_1441),
.B2(n_1414),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2928),
.B(n_2200),
.Y(n_3127)
);

NOR2xp33_ASAP7_75t_L g3128 ( 
.A(n_2912),
.B(n_2500),
.Y(n_3128)
);

AOI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2805),
.A2(n_2202),
.B1(n_2211),
.B2(n_2207),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2848),
.Y(n_3130)
);

HB1xp67_ASAP7_75t_L g3131 ( 
.A(n_2948),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_2992),
.B(n_2502),
.Y(n_3132)
);

INVx3_ASAP7_75t_L g3133 ( 
.A(n_2777),
.Y(n_3133)
);

INVx2_ASAP7_75t_SL g3134 ( 
.A(n_2972),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2857),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2982),
.B(n_2213),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2892),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2914),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_2915),
.B(n_2759),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2887),
.B(n_2815),
.Y(n_3140)
);

NOR2xp33_ASAP7_75t_L g3141 ( 
.A(n_2917),
.B(n_1414),
.Y(n_3141)
);

AOI22xp33_ASAP7_75t_L g3142 ( 
.A1(n_2971),
.A2(n_1450),
.B1(n_1457),
.B2(n_1445),
.Y(n_3142)
);

NOR3xp33_ASAP7_75t_L g3143 ( 
.A(n_2879),
.B(n_2608),
.C(n_2488),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2930),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2960),
.Y(n_3145)
);

NAND2xp33_ASAP7_75t_L g3146 ( 
.A(n_2920),
.B(n_2274),
.Y(n_3146)
);

OAI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_2894),
.A2(n_1450),
.B1(n_1457),
.B2(n_1445),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2952),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2964),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2887),
.B(n_2218),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2903),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2916),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2970),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_2925),
.B(n_2927),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_2936),
.B(n_2804),
.Y(n_3155)
);

INVx2_ASAP7_75t_SL g3156 ( 
.A(n_2972),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_SL g3157 ( 
.A(n_2804),
.B(n_2759),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2887),
.B(n_2221),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2965),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2886),
.B(n_2233),
.Y(n_3160)
);

INVxp33_ASAP7_75t_L g3161 ( 
.A(n_2874),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2981),
.Y(n_3162)
);

INVxp67_ASAP7_75t_L g3163 ( 
.A(n_2907),
.Y(n_3163)
);

NOR2xp33_ASAP7_75t_L g3164 ( 
.A(n_2969),
.B(n_2953),
.Y(n_3164)
);

OAI22xp33_ASAP7_75t_L g3165 ( 
.A1(n_3010),
.A2(n_1468),
.B1(n_1506),
.B2(n_1459),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2921),
.Y(n_3166)
);

NOR2xp33_ASAP7_75t_L g3167 ( 
.A(n_2831),
.B(n_1459),
.Y(n_3167)
);

NOR3xp33_ASAP7_75t_L g3168 ( 
.A(n_2918),
.B(n_2681),
.C(n_2680),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_L g3169 ( 
.A(n_2796),
.B(n_1468),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2920),
.B(n_2235),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2920),
.B(n_2236),
.Y(n_3171)
);

AOI22xp33_ASAP7_75t_L g3172 ( 
.A1(n_2787),
.A2(n_1521),
.B1(n_1523),
.B2(n_1506),
.Y(n_3172)
);

BUFx6f_ASAP7_75t_L g3173 ( 
.A(n_2777),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2938),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_SL g3175 ( 
.A(n_2845),
.B(n_2258),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2937),
.B(n_2940),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2983),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2937),
.B(n_2262),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_SL g3179 ( 
.A(n_2846),
.B(n_2237),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2961),
.Y(n_3180)
);

NAND2xp33_ASAP7_75t_L g3181 ( 
.A(n_2937),
.B(n_2940),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_R g3182 ( 
.A(n_2929),
.B(n_2650),
.Y(n_3182)
);

INVx2_ASAP7_75t_SL g3183 ( 
.A(n_2997),
.Y(n_3183)
);

INVxp67_ASAP7_75t_SL g3184 ( 
.A(n_2778),
.Y(n_3184)
);

INVx2_ASAP7_75t_SL g3185 ( 
.A(n_2997),
.Y(n_3185)
);

NOR2xp33_ASAP7_75t_L g3186 ( 
.A(n_2800),
.B(n_1521),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2940),
.B(n_2248),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2962),
.B(n_2415),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_2974),
.Y(n_3189)
);

NOR2xp33_ASAP7_75t_L g3190 ( 
.A(n_2978),
.B(n_1523),
.Y(n_3190)
);

INVxp67_ASAP7_75t_L g3191 ( 
.A(n_2934),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_L g3192 ( 
.A(n_2850),
.B(n_1530),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_3006),
.B(n_2420),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2991),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3016),
.B(n_2454),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2812),
.Y(n_3196)
);

INVx2_ASAP7_75t_SL g3197 ( 
.A(n_2851),
.Y(n_3197)
);

CKINVDCx5p33_ASAP7_75t_R g3198 ( 
.A(n_2811),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_2932),
.B(n_1590),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_SL g3200 ( 
.A(n_2867),
.B(n_1530),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2999),
.Y(n_3201)
);

NOR2xp33_ASAP7_75t_L g3202 ( 
.A(n_2944),
.B(n_1617),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2924),
.B(n_2457),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2931),
.B(n_2763),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2957),
.B(n_2162),
.Y(n_3205)
);

AOI22xp33_ASAP7_75t_L g3206 ( 
.A1(n_2889),
.A2(n_1649),
.B1(n_1671),
.B2(n_1617),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2990),
.B(n_1172),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_3001),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_2866),
.B(n_1590),
.Y(n_3209)
);

AOI22xp33_ASAP7_75t_L g3210 ( 
.A1(n_2895),
.A2(n_1671),
.B1(n_1674),
.B2(n_1649),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2998),
.B(n_1175),
.Y(n_3211)
);

INVxp67_ASAP7_75t_L g3212 ( 
.A(n_2935),
.Y(n_3212)
);

NAND3xp33_ASAP7_75t_L g3213 ( 
.A(n_2913),
.B(n_1177),
.C(n_1176),
.Y(n_3213)
);

NOR2xp33_ASAP7_75t_L g3214 ( 
.A(n_2966),
.B(n_1674),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_2967),
.B(n_1701),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_2896),
.B(n_1633),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3012),
.B(n_1178),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2905),
.B(n_1179),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_SL g3219 ( 
.A(n_2919),
.B(n_1701),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3043),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3028),
.B(n_2923),
.Y(n_3221)
);

INVx3_ASAP7_75t_L g3222 ( 
.A(n_3125),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_3034),
.B(n_2843),
.Y(n_3223)
);

AOI22xp5_ASAP7_75t_L g3224 ( 
.A1(n_3053),
.A2(n_2976),
.B1(n_2943),
.B2(n_2968),
.Y(n_3224)
);

A2O1A1Ixp33_ASAP7_75t_L g3225 ( 
.A1(n_3154),
.A2(n_2906),
.B(n_2946),
.C(n_2801),
.Y(n_3225)
);

OAI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_3059),
.A2(n_2856),
.B(n_3005),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3066),
.B(n_3004),
.Y(n_3227)
);

AOI22xp5_ASAP7_75t_L g3228 ( 
.A1(n_3019),
.A2(n_2950),
.B1(n_2987),
.B2(n_2821),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_3017),
.B(n_3035),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3029),
.B(n_3007),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3030),
.Y(n_3231)
);

OAI22xp5_ASAP7_75t_L g3232 ( 
.A1(n_3206),
.A2(n_2854),
.B1(n_2963),
.B2(n_2951),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3062),
.B(n_3008),
.Y(n_3233)
);

BUFx2_ASAP7_75t_L g3234 ( 
.A(n_3032),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_3120),
.B(n_3011),
.Y(n_3235)
);

A2O1A1Ixp33_ASAP7_75t_L g3236 ( 
.A1(n_3042),
.A2(n_3015),
.B(n_3014),
.C(n_2790),
.Y(n_3236)
);

NOR2xp33_ASAP7_75t_L g3237 ( 
.A(n_3064),
.B(n_2949),
.Y(n_3237)
);

INVx3_ASAP7_75t_L g3238 ( 
.A(n_3173),
.Y(n_3238)
);

BUFx6f_ASAP7_75t_L g3239 ( 
.A(n_3173),
.Y(n_3239)
);

AOI21xp5_ASAP7_75t_L g3240 ( 
.A1(n_3136),
.A2(n_2774),
.B(n_2891),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_SL g3241 ( 
.A(n_3045),
.B(n_2871),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_3092),
.A2(n_2844),
.B(n_2785),
.Y(n_3242)
);

BUFx8_ASAP7_75t_L g3243 ( 
.A(n_3068),
.Y(n_3243)
);

OAI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3038),
.A2(n_2870),
.B(n_2882),
.Y(n_3244)
);

INVx3_ASAP7_75t_L g3245 ( 
.A(n_3173),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_3122),
.B(n_3123),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3127),
.B(n_2885),
.Y(n_3247)
);

A2O1A1Ixp33_ASAP7_75t_L g3248 ( 
.A1(n_3141),
.A2(n_3009),
.B(n_2893),
.C(n_2849),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3044),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3096),
.B(n_2828),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3046),
.B(n_2778),
.Y(n_3251)
);

OAI22xp5_ASAP7_75t_L g3252 ( 
.A1(n_3033),
.A2(n_2794),
.B1(n_2807),
.B2(n_2789),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3057),
.B(n_2789),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_3025),
.A2(n_2807),
.B(n_2794),
.Y(n_3254)
);

OAI22xp5_ASAP7_75t_L g3255 ( 
.A1(n_3022),
.A2(n_2842),
.B1(n_2852),
.B2(n_2832),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_3061),
.B(n_2832),
.Y(n_3256)
);

BUFx4f_ASAP7_75t_L g3257 ( 
.A(n_3077),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3065),
.B(n_2842),
.Y(n_3258)
);

AOI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_3205),
.A2(n_2853),
.B(n_2852),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3083),
.Y(n_3260)
);

OAI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_3140),
.A2(n_3112),
.B(n_3109),
.Y(n_3261)
);

NOR2xp33_ASAP7_75t_L g3262 ( 
.A(n_3020),
.B(n_2884),
.Y(n_3262)
);

AO21x1_ASAP7_75t_L g3263 ( 
.A1(n_3027),
.A2(n_1135),
.B(n_1115),
.Y(n_3263)
);

O2A1O1Ixp5_ASAP7_75t_L g3264 ( 
.A1(n_3063),
.A2(n_1880),
.B(n_1896),
.C(n_1776),
.Y(n_3264)
);

AOI22xp33_ASAP7_75t_L g3265 ( 
.A1(n_3023),
.A2(n_3041),
.B1(n_3036),
.B2(n_3072),
.Y(n_3265)
);

BUFx2_ASAP7_75t_L g3266 ( 
.A(n_3018),
.Y(n_3266)
);

AOI21xp5_ASAP7_75t_L g3267 ( 
.A1(n_3058),
.A2(n_2853),
.B(n_2973),
.Y(n_3267)
);

O2A1O1Ixp33_ASAP7_75t_L g3268 ( 
.A1(n_3052),
.A2(n_1143),
.B(n_1145),
.C(n_1137),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_3040),
.B(n_3002),
.Y(n_3269)
);

AOI21xp5_ASAP7_75t_L g3270 ( 
.A1(n_3095),
.A2(n_3003),
.B(n_2979),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3088),
.Y(n_3271)
);

BUFx3_ASAP7_75t_L g3272 ( 
.A(n_3098),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_3090),
.B(n_2984),
.Y(n_3273)
);

CKINVDCx20_ASAP7_75t_R g3274 ( 
.A(n_3198),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3050),
.Y(n_3275)
);

NOR2xp33_ASAP7_75t_L g3276 ( 
.A(n_3190),
.B(n_2792),
.Y(n_3276)
);

OAI21xp5_ASAP7_75t_L g3277 ( 
.A1(n_3099),
.A2(n_2988),
.B(n_2984),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3101),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3104),
.B(n_2984),
.Y(n_3279)
);

OAI321xp33_ASAP7_75t_L g3280 ( 
.A1(n_3126),
.A2(n_1161),
.A3(n_1150),
.B1(n_1171),
.B2(n_1158),
.C(n_1149),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_3095),
.A2(n_2810),
.B(n_2980),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_3054),
.B(n_1711),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_3056),
.A2(n_1174),
.B(n_1173),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3105),
.Y(n_3284)
);

AND2x4_ASAP7_75t_L g3285 ( 
.A(n_3196),
.B(n_2988),
.Y(n_3285)
);

AOI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_3069),
.A2(n_1184),
.B(n_1183),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3107),
.B(n_2988),
.Y(n_3287)
);

O2A1O1Ixp5_ASAP7_75t_L g3288 ( 
.A1(n_3175),
.A2(n_1880),
.B(n_1896),
.C(n_1776),
.Y(n_3288)
);

NOR2x1p5_ASAP7_75t_L g3289 ( 
.A(n_3026),
.B(n_2881),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_3110),
.B(n_1633),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3073),
.Y(n_3291)
);

AOI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_3070),
.A2(n_3181),
.B(n_3160),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3130),
.B(n_1180),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3081),
.A2(n_1194),
.B(n_1187),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3145),
.B(n_1182),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3149),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3085),
.A2(n_1198),
.B(n_1197),
.Y(n_3297)
);

NOR2xp33_ASAP7_75t_SL g3298 ( 
.A(n_3079),
.B(n_2662),
.Y(n_3298)
);

AO21x1_ASAP7_75t_L g3299 ( 
.A1(n_3150),
.A2(n_1212),
.B(n_1208),
.Y(n_3299)
);

INVx11_ASAP7_75t_L g3300 ( 
.A(n_3098),
.Y(n_3300)
);

AOI22xp33_ASAP7_75t_L g3301 ( 
.A1(n_3021),
.A2(n_3047),
.B1(n_3119),
.B2(n_3060),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3039),
.B(n_1186),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3078),
.Y(n_3303)
);

NAND2x1p5_ASAP7_75t_L g3304 ( 
.A(n_3197),
.B(n_1220),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3084),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3164),
.B(n_1188),
.Y(n_3306)
);

AOI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_3115),
.A2(n_1232),
.B(n_1222),
.Y(n_3307)
);

AOI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_3118),
.A2(n_1240),
.B(n_1236),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_SL g3309 ( 
.A(n_3051),
.B(n_1711),
.Y(n_3309)
);

OAI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_3117),
.A2(n_2182),
.B(n_1244),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3091),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3159),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3097),
.B(n_1190),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_3176),
.A2(n_1247),
.B(n_1241),
.Y(n_3314)
);

HB1xp67_ASAP7_75t_L g3315 ( 
.A(n_3103),
.Y(n_3315)
);

INVx3_ASAP7_75t_L g3316 ( 
.A(n_3100),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_3055),
.B(n_1191),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3162),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3177),
.Y(n_3319)
);

NOR2x2_ASAP7_75t_L g3320 ( 
.A(n_3135),
.B(n_1904),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3194),
.Y(n_3321)
);

OR2x2_ASAP7_75t_SL g3322 ( 
.A(n_3131),
.B(n_1904),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3199),
.B(n_1192),
.Y(n_3323)
);

AOI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_3139),
.A2(n_1250),
.B(n_1249),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_3163),
.B(n_1193),
.Y(n_3325)
);

AOI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_3049),
.A2(n_1265),
.B(n_1251),
.Y(n_3326)
);

NOR2xp67_ASAP7_75t_SL g3327 ( 
.A(n_3082),
.B(n_1916),
.Y(n_3327)
);

AND2x4_ASAP7_75t_L g3328 ( 
.A(n_3134),
.B(n_1269),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_SL g3329 ( 
.A(n_3116),
.B(n_1728),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3151),
.B(n_1199),
.Y(n_3330)
);

INVx3_ASAP7_75t_L g3331 ( 
.A(n_3133),
.Y(n_3331)
);

INVx3_ASAP7_75t_L g3332 ( 
.A(n_3156),
.Y(n_3332)
);

AOI22xp5_ASAP7_75t_L g3333 ( 
.A1(n_3191),
.A2(n_1738),
.B1(n_1768),
.B2(n_1728),
.Y(n_3333)
);

NOR3xp33_ASAP7_75t_L g3334 ( 
.A(n_3192),
.B(n_1202),
.C(n_1201),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3146),
.A2(n_1272),
.B(n_1271),
.Y(n_3335)
);

OR2x2_ASAP7_75t_L g3336 ( 
.A(n_3114),
.B(n_1204),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_3152),
.Y(n_3337)
);

OAI21xp33_ASAP7_75t_L g3338 ( 
.A1(n_3142),
.A2(n_3172),
.B(n_3210),
.Y(n_3338)
);

AOI22xp33_ASAP7_75t_L g3339 ( 
.A1(n_3089),
.A2(n_1768),
.B1(n_1792),
.B2(n_1738),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3166),
.B(n_1206),
.Y(n_3340)
);

NAND2xp33_ASAP7_75t_L g3341 ( 
.A(n_3121),
.B(n_1207),
.Y(n_3341)
);

O2A1O1Ixp33_ASAP7_75t_L g3342 ( 
.A1(n_3212),
.A2(n_3074),
.B(n_3218),
.C(n_3165),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3174),
.B(n_1209),
.Y(n_3343)
);

BUFx2_ASAP7_75t_L g3344 ( 
.A(n_3184),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3201),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3180),
.B(n_1211),
.Y(n_3346)
);

AOI21xp5_ASAP7_75t_L g3347 ( 
.A1(n_3170),
.A2(n_1274),
.B(n_1273),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3189),
.B(n_1213),
.Y(n_3348)
);

AOI21xp5_ASAP7_75t_L g3349 ( 
.A1(n_3171),
.A2(n_1284),
.B(n_1278),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3111),
.B(n_1214),
.Y(n_3350)
);

INVx3_ASAP7_75t_L g3351 ( 
.A(n_3183),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_3178),
.A2(n_1291),
.B(n_1287),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3187),
.A2(n_1306),
.B(n_1304),
.Y(n_3353)
);

INVx4_ASAP7_75t_L g3354 ( 
.A(n_3185),
.Y(n_3354)
);

AND2x2_ASAP7_75t_SL g3355 ( 
.A(n_3124),
.B(n_3093),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_3102),
.A2(n_1311),
.B(n_1309),
.Y(n_3356)
);

OAI22xp5_ASAP7_75t_L g3357 ( 
.A1(n_3208),
.A2(n_1799),
.B1(n_1833),
.B2(n_1792),
.Y(n_3357)
);

AND2x4_ASAP7_75t_L g3358 ( 
.A(n_3137),
.B(n_3138),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3094),
.B(n_1215),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_3067),
.B(n_1799),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3106),
.B(n_1218),
.Y(n_3361)
);

AOI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_3207),
.A2(n_1317),
.B(n_1314),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3108),
.B(n_1221),
.Y(n_3363)
);

NOR2xp33_ASAP7_75t_L g3364 ( 
.A(n_3167),
.B(n_3202),
.Y(n_3364)
);

AOI22xp33_ASAP7_75t_L g3365 ( 
.A1(n_3147),
.A2(n_1857),
.B1(n_1862),
.B2(n_1833),
.Y(n_3365)
);

AOI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3214),
.A2(n_1862),
.B1(n_1867),
.B2(n_1857),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3132),
.B(n_1633),
.Y(n_3367)
);

NOR2xp33_ASAP7_75t_L g3368 ( 
.A(n_3169),
.B(n_1867),
.Y(n_3368)
);

AOI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_3211),
.A2(n_1324),
.B(n_1321),
.Y(n_3369)
);

BUFx3_ASAP7_75t_L g3370 ( 
.A(n_3209),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3186),
.B(n_1226),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_R g3372 ( 
.A(n_3274),
.B(n_3031),
.Y(n_3372)
);

INVx3_ASAP7_75t_L g3373 ( 
.A(n_3257),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3220),
.Y(n_3374)
);

BUFx4f_ASAP7_75t_L g3375 ( 
.A(n_3239),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_3364),
.B(n_3161),
.Y(n_3376)
);

OR2x6_ASAP7_75t_L g3377 ( 
.A(n_3272),
.B(n_3113),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3246),
.B(n_3128),
.Y(n_3378)
);

BUFx2_ASAP7_75t_L g3379 ( 
.A(n_3234),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_3221),
.B(n_3217),
.Y(n_3380)
);

AND2x4_ASAP7_75t_SL g3381 ( 
.A(n_3315),
.B(n_3216),
.Y(n_3381)
);

O2A1O1Ixp33_ASAP7_75t_L g3382 ( 
.A1(n_3368),
.A2(n_3200),
.B(n_3215),
.C(n_3219),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3229),
.B(n_3076),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3233),
.B(n_3071),
.Y(n_3384)
);

OAI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_3366),
.A2(n_3087),
.B1(n_3213),
.B2(n_3086),
.Y(n_3385)
);

BUFx2_ASAP7_75t_L g3386 ( 
.A(n_3266),
.Y(n_3386)
);

AOI21xp5_ASAP7_75t_L g3387 ( 
.A1(n_3292),
.A2(n_3037),
.B(n_3075),
.Y(n_3387)
);

AND2x4_ASAP7_75t_L g3388 ( 
.A(n_3285),
.B(n_3048),
.Y(n_3388)
);

A2O1A1Ixp33_ASAP7_75t_L g3389 ( 
.A1(n_3342),
.A2(n_3158),
.B(n_3080),
.C(n_3188),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_L g3390 ( 
.A(n_3262),
.B(n_3155),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_3226),
.A2(n_3179),
.B(n_3203),
.Y(n_3391)
);

O2A1O1Ixp33_ASAP7_75t_L g3392 ( 
.A1(n_3241),
.A2(n_3143),
.B(n_3204),
.C(n_3168),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3306),
.B(n_3144),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3260),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3271),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3227),
.B(n_3148),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_3240),
.A2(n_3121),
.B(n_3193),
.Y(n_3397)
);

AOI21xp5_ASAP7_75t_L g3398 ( 
.A1(n_3261),
.A2(n_3121),
.B(n_3195),
.Y(n_3398)
);

CKINVDCx5p33_ASAP7_75t_R g3399 ( 
.A(n_3300),
.Y(n_3399)
);

NOR2xp33_ASAP7_75t_R g3400 ( 
.A(n_3298),
.B(n_3153),
.Y(n_3400)
);

OAI22xp5_ASAP7_75t_SL g3401 ( 
.A1(n_3339),
.A2(n_1879),
.B1(n_1886),
.B2(n_1871),
.Y(n_3401)
);

INVx3_ASAP7_75t_L g3402 ( 
.A(n_3354),
.Y(n_3402)
);

INVx3_ASAP7_75t_L g3403 ( 
.A(n_3354),
.Y(n_3403)
);

OR2x2_ASAP7_75t_L g3404 ( 
.A(n_3313),
.B(n_3157),
.Y(n_3404)
);

BUFx3_ASAP7_75t_L g3405 ( 
.A(n_3243),
.Y(n_3405)
);

OAI21xp33_ASAP7_75t_L g3406 ( 
.A1(n_3365),
.A2(n_1879),
.B(n_1871),
.Y(n_3406)
);

NAND3xp33_ASAP7_75t_L g3407 ( 
.A(n_3334),
.B(n_3024),
.C(n_3129),
.Y(n_3407)
);

A2O1A1Ixp33_ASAP7_75t_L g3408 ( 
.A1(n_3338),
.A2(n_1334),
.B(n_1335),
.C(n_1328),
.Y(n_3408)
);

O2A1O1Ixp33_ASAP7_75t_L g3409 ( 
.A1(n_3282),
.A2(n_1342),
.B(n_1345),
.C(n_1341),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_3278),
.Y(n_3410)
);

OR2x6_ASAP7_75t_L g3411 ( 
.A(n_3370),
.B(n_3182),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_3223),
.B(n_1886),
.Y(n_3412)
);

CKINVDCx14_ASAP7_75t_R g3413 ( 
.A(n_3269),
.Y(n_3413)
);

BUFx3_ASAP7_75t_L g3414 ( 
.A(n_3243),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_3276),
.B(n_1233),
.Y(n_3415)
);

CKINVDCx5p33_ASAP7_75t_R g3416 ( 
.A(n_3289),
.Y(n_3416)
);

AOI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_3341),
.A2(n_3121),
.B(n_1349),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3284),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3265),
.B(n_3121),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_SL g3420 ( 
.A(n_3224),
.B(n_1720),
.Y(n_3420)
);

AOI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_3225),
.A2(n_1351),
.B(n_1346),
.Y(n_3421)
);

BUFx2_ASAP7_75t_L g3422 ( 
.A(n_3239),
.Y(n_3422)
);

A2O1A1Ixp33_ASAP7_75t_L g3423 ( 
.A1(n_3242),
.A2(n_1354),
.B(n_1360),
.C(n_1353),
.Y(n_3423)
);

OAI21x1_ASAP7_75t_L g3424 ( 
.A1(n_3259),
.A2(n_1916),
.B(n_1919),
.Y(n_3424)
);

OAI22xp5_ASAP7_75t_L g3425 ( 
.A1(n_3301),
.A2(n_1237),
.B1(n_1238),
.B2(n_1235),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3296),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_3310),
.A2(n_1379),
.B(n_1374),
.Y(n_3427)
);

NOR2x1_ASAP7_75t_L g3428 ( 
.A(n_3247),
.B(n_1384),
.Y(n_3428)
);

BUFx2_ASAP7_75t_L g3429 ( 
.A(n_3239),
.Y(n_3429)
);

OAI22xp5_ASAP7_75t_L g3430 ( 
.A1(n_3230),
.A2(n_1245),
.B1(n_1246),
.B2(n_1239),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_R g3431 ( 
.A(n_3316),
.B(n_996),
.Y(n_3431)
);

A2O1A1Ixp33_ASAP7_75t_L g3432 ( 
.A1(n_3236),
.A2(n_1403),
.B(n_1404),
.C(n_1399),
.Y(n_3432)
);

AND2x4_ASAP7_75t_SL g3433 ( 
.A(n_3222),
.B(n_1720),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_3235),
.A2(n_1410),
.B(n_1405),
.Y(n_3434)
);

A2O1A1Ixp33_ASAP7_75t_L g3435 ( 
.A1(n_3280),
.A2(n_1437),
.B(n_1438),
.C(n_1423),
.Y(n_3435)
);

INVx3_ASAP7_75t_L g3436 ( 
.A(n_3332),
.Y(n_3436)
);

NOR2x1_ASAP7_75t_SL g3437 ( 
.A(n_3273),
.B(n_3279),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_SL g3438 ( 
.A(n_3237),
.B(n_1720),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_3232),
.B(n_3228),
.Y(n_3439)
);

BUFx6f_ASAP7_75t_L g3440 ( 
.A(n_3238),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3312),
.Y(n_3441)
);

INVx5_ASAP7_75t_L g3442 ( 
.A(n_3245),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3367),
.B(n_1769),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_SL g3444 ( 
.A(n_3358),
.B(n_1769),
.Y(n_3444)
);

CKINVDCx5p33_ASAP7_75t_R g3445 ( 
.A(n_3355),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3318),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3319),
.Y(n_3447)
);

OAI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_3264),
.A2(n_2182),
.B(n_1447),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3244),
.A2(n_1452),
.B(n_1440),
.Y(n_3449)
);

INVx3_ASAP7_75t_L g3450 ( 
.A(n_3351),
.Y(n_3450)
);

A2O1A1Ixp33_ASAP7_75t_L g3451 ( 
.A1(n_3371),
.A2(n_1454),
.B(n_1465),
.C(n_1453),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3350),
.B(n_1469),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3321),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3250),
.A2(n_1252),
.B1(n_1253),
.B2(n_1248),
.Y(n_3454)
);

NOR2xp33_ASAP7_75t_R g3455 ( 
.A(n_3331),
.B(n_1000),
.Y(n_3455)
);

INVxp67_ASAP7_75t_SL g3456 ( 
.A(n_3251),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3360),
.B(n_1769),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_R g3458 ( 
.A(n_3344),
.B(n_1002),
.Y(n_3458)
);

AOI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_3254),
.A2(n_1474),
.B(n_1471),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3359),
.B(n_1488),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3345),
.Y(n_3461)
);

OAI22xp5_ASAP7_75t_L g3462 ( 
.A1(n_3361),
.A2(n_1256),
.B1(n_1257),
.B2(n_1254),
.Y(n_3462)
);

BUFx6f_ASAP7_75t_L g3463 ( 
.A(n_3358),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3363),
.B(n_1490),
.Y(n_3464)
);

AO21x1_ASAP7_75t_L g3465 ( 
.A1(n_3314),
.A2(n_1499),
.B(n_1498),
.Y(n_3465)
);

O2A1O1Ixp5_ASAP7_75t_SL g3466 ( 
.A1(n_3277),
.A2(n_3252),
.B(n_3309),
.C(n_3329),
.Y(n_3466)
);

NOR3xp33_ASAP7_75t_SL g3467 ( 
.A(n_3357),
.B(n_1263),
.C(n_1260),
.Y(n_3467)
);

OAI22x1_ASAP7_75t_L g3468 ( 
.A1(n_3333),
.A2(n_1266),
.B1(n_1267),
.B2(n_1264),
.Y(n_3468)
);

AOI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_3263),
.A2(n_1846),
.B1(n_1865),
.B2(n_1813),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_3267),
.A2(n_1507),
.B(n_1504),
.Y(n_3470)
);

AND2x4_ASAP7_75t_L g3471 ( 
.A(n_3285),
.B(n_1508),
.Y(n_3471)
);

NOR2xp33_ASAP7_75t_L g3472 ( 
.A(n_3302),
.B(n_1268),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_SL g3473 ( 
.A(n_3323),
.B(n_1813),
.Y(n_3473)
);

O2A1O1Ixp33_ASAP7_75t_L g3474 ( 
.A1(n_3248),
.A2(n_1520),
.B(n_1522),
.C(n_1511),
.Y(n_3474)
);

A2O1A1Ixp33_ASAP7_75t_L g3475 ( 
.A1(n_3287),
.A2(n_1533),
.B(n_1539),
.C(n_1527),
.Y(n_3475)
);

A2O1A1Ixp33_ASAP7_75t_SL g3476 ( 
.A1(n_3327),
.A2(n_1544),
.B(n_1550),
.C(n_1543),
.Y(n_3476)
);

CKINVDCx5p33_ASAP7_75t_R g3477 ( 
.A(n_3281),
.Y(n_3477)
);

A2O1A1Ixp33_ASAP7_75t_L g3478 ( 
.A1(n_3317),
.A2(n_1574),
.B(n_1578),
.C(n_1563),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3231),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3294),
.B(n_1579),
.Y(n_3480)
);

AOI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_3335),
.A2(n_1591),
.B(n_1588),
.Y(n_3481)
);

OAI22xp5_ASAP7_75t_L g3482 ( 
.A1(n_3253),
.A2(n_1275),
.B1(n_1277),
.B2(n_1270),
.Y(n_3482)
);

A2O1A1Ixp33_ASAP7_75t_L g3483 ( 
.A1(n_3297),
.A2(n_3283),
.B(n_3286),
.C(n_3353),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_3336),
.B(n_1813),
.Y(n_3484)
);

BUFx2_ASAP7_75t_L g3485 ( 
.A(n_3322),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3270),
.A2(n_1614),
.B(n_1593),
.Y(n_3486)
);

OAI22xp5_ASAP7_75t_L g3487 ( 
.A1(n_3256),
.A2(n_1281),
.B1(n_1283),
.B2(n_1279),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3328),
.A2(n_1865),
.B1(n_1903),
.B2(n_1846),
.Y(n_3488)
);

BUFx6f_ASAP7_75t_L g3489 ( 
.A(n_3328),
.Y(n_3489)
);

NOR2xp67_ASAP7_75t_SL g3490 ( 
.A(n_3290),
.B(n_1285),
.Y(n_3490)
);

NAND3xp33_ASAP7_75t_L g3491 ( 
.A(n_3326),
.B(n_1294),
.C(n_1286),
.Y(n_3491)
);

INVx3_ASAP7_75t_SL g3492 ( 
.A(n_3320),
.Y(n_3492)
);

BUFx2_ASAP7_75t_L g3493 ( 
.A(n_3304),
.Y(n_3493)
);

BUFx6f_ASAP7_75t_L g3494 ( 
.A(n_3258),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3303),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3249),
.B(n_1846),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_SL g3497 ( 
.A(n_3275),
.B(n_1865),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_SL g3498 ( 
.A(n_3291),
.B(n_1903),
.Y(n_3498)
);

INVx4_ASAP7_75t_L g3499 ( 
.A(n_3311),
.Y(n_3499)
);

NOR2xp33_ASAP7_75t_L g3500 ( 
.A(n_3325),
.B(n_1298),
.Y(n_3500)
);

AOI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_3330),
.A2(n_3343),
.B(n_3340),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3337),
.Y(n_3502)
);

CKINVDCx5p33_ASAP7_75t_R g3503 ( 
.A(n_3305),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3293),
.B(n_1616),
.Y(n_3504)
);

AOI21x1_ASAP7_75t_L g3505 ( 
.A1(n_3299),
.A2(n_1623),
.B(n_1618),
.Y(n_3505)
);

NOR2xp33_ASAP7_75t_L g3506 ( 
.A(n_3295),
.B(n_1299),
.Y(n_3506)
);

AOI21xp5_ASAP7_75t_L g3507 ( 
.A1(n_3346),
.A2(n_1637),
.B(n_1636),
.Y(n_3507)
);

NOR2xp67_ASAP7_75t_SL g3508 ( 
.A(n_3348),
.B(n_1301),
.Y(n_3508)
);

BUFx12f_ASAP7_75t_L g3509 ( 
.A(n_3268),
.Y(n_3509)
);

OAI21x1_ASAP7_75t_L g3510 ( 
.A1(n_3288),
.A2(n_1909),
.B(n_1905),
.Y(n_3510)
);

CKINVDCx16_ASAP7_75t_R g3511 ( 
.A(n_3255),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3378),
.B(n_3356),
.Y(n_3512)
);

BUFx2_ASAP7_75t_L g3513 ( 
.A(n_3379),
.Y(n_3513)
);

NOR4xp25_ASAP7_75t_L g3514 ( 
.A(n_3382),
.B(n_1640),
.C(n_1641),
.D(n_1639),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3410),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_3501),
.A2(n_3369),
.B(n_3362),
.Y(n_3516)
);

INVxp67_ASAP7_75t_SL g3517 ( 
.A(n_3456),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3376),
.B(n_3307),
.Y(n_3518)
);

OAI21x1_ASAP7_75t_L g3519 ( 
.A1(n_3397),
.A2(n_3347),
.B(n_3308),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3441),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3415),
.B(n_3349),
.Y(n_3521)
);

BUFx2_ASAP7_75t_L g3522 ( 
.A(n_3386),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_R g3523 ( 
.A(n_3413),
.B(n_1006),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3384),
.B(n_3352),
.Y(n_3524)
);

AND2x2_ASAP7_75t_L g3525 ( 
.A(n_3443),
.B(n_3471),
.Y(n_3525)
);

CKINVDCx5p33_ASAP7_75t_R g3526 ( 
.A(n_3416),
.Y(n_3526)
);

AO31x2_ASAP7_75t_L g3527 ( 
.A1(n_3432),
.A2(n_3324),
.A3(n_1654),
.B(n_1658),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3447),
.Y(n_3528)
);

OAI22xp5_ASAP7_75t_L g3529 ( 
.A1(n_3390),
.A2(n_1303),
.B1(n_1305),
.B2(n_1302),
.Y(n_3529)
);

BUFx3_ASAP7_75t_L g3530 ( 
.A(n_3373),
.Y(n_3530)
);

INVx2_ASAP7_75t_SL g3531 ( 
.A(n_3440),
.Y(n_3531)
);

CKINVDCx8_ASAP7_75t_R g3532 ( 
.A(n_3399),
.Y(n_3532)
);

BUFx2_ASAP7_75t_L g3533 ( 
.A(n_3503),
.Y(n_3533)
);

AO31x2_ASAP7_75t_L g3534 ( 
.A1(n_3449),
.A2(n_1660),
.A3(n_1662),
.B(n_1645),
.Y(n_3534)
);

NOR2xp33_ASAP7_75t_L g3535 ( 
.A(n_3412),
.B(n_1307),
.Y(n_3535)
);

OAI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3439),
.A2(n_1668),
.B(n_1667),
.Y(n_3536)
);

OAI21x1_ASAP7_75t_L g3537 ( 
.A1(n_3398),
.A2(n_1679),
.B(n_1673),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3380),
.B(n_3406),
.Y(n_3538)
);

OAI21x1_ASAP7_75t_L g3539 ( 
.A1(n_3424),
.A2(n_1692),
.B(n_1681),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3472),
.B(n_1308),
.Y(n_3540)
);

OAI21x1_ASAP7_75t_L g3541 ( 
.A1(n_3510),
.A2(n_1703),
.B(n_1700),
.Y(n_3541)
);

INVx1_ASAP7_75t_SL g3542 ( 
.A(n_3381),
.Y(n_3542)
);

OAI21x1_ASAP7_75t_L g3543 ( 
.A1(n_3391),
.A2(n_1706),
.B(n_1705),
.Y(n_3543)
);

O2A1O1Ixp33_ASAP7_75t_SL g3544 ( 
.A1(n_3483),
.A2(n_1714),
.B(n_1716),
.C(n_1712),
.Y(n_3544)
);

NOR2xp33_ASAP7_75t_L g3545 ( 
.A(n_3445),
.B(n_1310),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_3511),
.B(n_1903),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3506),
.B(n_1312),
.Y(n_3547)
);

OAI21x1_ASAP7_75t_L g3548 ( 
.A1(n_3387),
.A2(n_1731),
.B(n_1730),
.Y(n_3548)
);

NOR2xp33_ASAP7_75t_L g3549 ( 
.A(n_3492),
.B(n_1313),
.Y(n_3549)
);

INVx3_ASAP7_75t_SL g3550 ( 
.A(n_3411),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3374),
.Y(n_3551)
);

OAI21x1_ASAP7_75t_L g3552 ( 
.A1(n_3417),
.A2(n_1740),
.B(n_1732),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3394),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_L g3554 ( 
.A(n_3401),
.B(n_1315),
.Y(n_3554)
);

OAI21x1_ASAP7_75t_L g3555 ( 
.A1(n_3421),
.A2(n_1748),
.B(n_1744),
.Y(n_3555)
);

HB1xp67_ASAP7_75t_L g3556 ( 
.A(n_3463),
.Y(n_3556)
);

BUFx6f_ASAP7_75t_L g3557 ( 
.A(n_3375),
.Y(n_3557)
);

CKINVDCx5p33_ASAP7_75t_R g3558 ( 
.A(n_3372),
.Y(n_3558)
);

OAI21x1_ASAP7_75t_L g3559 ( 
.A1(n_3505),
.A2(n_1754),
.B(n_1752),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3395),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3418),
.Y(n_3561)
);

AND2x2_ASAP7_75t_L g3562 ( 
.A(n_3471),
.B(n_1758),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_SL g3563 ( 
.A(n_3494),
.B(n_1918),
.Y(n_3563)
);

AO22x2_ASAP7_75t_L g3564 ( 
.A1(n_3420),
.A2(n_1765),
.B1(n_1767),
.B2(n_1763),
.Y(n_3564)
);

NAND3xp33_ASAP7_75t_L g3565 ( 
.A(n_3467),
.B(n_1318),
.C(n_1316),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3426),
.Y(n_3566)
);

INVx5_ASAP7_75t_L g3567 ( 
.A(n_3411),
.Y(n_3567)
);

INVx3_ASAP7_75t_L g3568 ( 
.A(n_3440),
.Y(n_3568)
);

OAI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_3466),
.A2(n_1774),
.B(n_1771),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3393),
.B(n_1319),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3419),
.A2(n_1783),
.B(n_1778),
.Y(n_3571)
);

OAI21x1_ASAP7_75t_L g3572 ( 
.A1(n_3474),
.A2(n_1789),
.B(n_1784),
.Y(n_3572)
);

AND2x2_ASAP7_75t_L g3573 ( 
.A(n_3457),
.B(n_1790),
.Y(n_3573)
);

NOR2xp67_ASAP7_75t_SL g3574 ( 
.A(n_3509),
.B(n_1320),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_3500),
.B(n_1323),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3396),
.B(n_1326),
.Y(n_3576)
);

OAI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_3389),
.A2(n_1809),
.B(n_1806),
.Y(n_3577)
);

AND2x2_ASAP7_75t_L g3578 ( 
.A(n_3485),
.B(n_1810),
.Y(n_3578)
);

OR2x2_ASAP7_75t_L g3579 ( 
.A(n_3460),
.B(n_1814),
.Y(n_3579)
);

AO21x2_ASAP7_75t_L g3580 ( 
.A1(n_3427),
.A2(n_1819),
.B(n_1816),
.Y(n_3580)
);

INVx4_ASAP7_75t_L g3581 ( 
.A(n_3442),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3464),
.B(n_1329),
.Y(n_3582)
);

BUFx6f_ASAP7_75t_L g3583 ( 
.A(n_3489),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3446),
.Y(n_3584)
);

AOI221xp5_ASAP7_75t_SL g3585 ( 
.A1(n_3385),
.A2(n_1831),
.B1(n_1837),
.B2(n_1829),
.C(n_1825),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3453),
.Y(n_3586)
);

AO31x2_ASAP7_75t_L g3587 ( 
.A1(n_3437),
.A2(n_1843),
.A3(n_1850),
.B(n_1840),
.Y(n_3587)
);

OR2x2_ASAP7_75t_L g3588 ( 
.A(n_3452),
.B(n_1853),
.Y(n_3588)
);

A2O1A1Ixp33_ASAP7_75t_L g3589 ( 
.A1(n_3392),
.A2(n_1856),
.B(n_1866),
.C(n_1854),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3461),
.Y(n_3590)
);

BUFx12f_ASAP7_75t_L g3591 ( 
.A(n_3405),
.Y(n_3591)
);

NOR2xp33_ASAP7_75t_L g3592 ( 
.A(n_3404),
.B(n_1330),
.Y(n_3592)
);

A2O1A1Ixp33_ASAP7_75t_L g3593 ( 
.A1(n_3407),
.A2(n_1876),
.B(n_1884),
.C(n_1868),
.Y(n_3593)
);

OAI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3383),
.A2(n_1893),
.B(n_1885),
.Y(n_3594)
);

OAI21x1_ASAP7_75t_L g3595 ( 
.A1(n_3470),
.A2(n_3459),
.B(n_3486),
.Y(n_3595)
);

INVx4_ASAP7_75t_L g3596 ( 
.A(n_3442),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3504),
.B(n_1331),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3495),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3473),
.A2(n_1900),
.B(n_1894),
.Y(n_3599)
);

NAND2x1p5_ASAP7_75t_L g3600 ( 
.A(n_3442),
.B(n_1911),
.Y(n_3600)
);

NOR2xp33_ASAP7_75t_L g3601 ( 
.A(n_3438),
.B(n_3494),
.Y(n_3601)
);

INVx3_ASAP7_75t_L g3602 ( 
.A(n_3463),
.Y(n_3602)
);

AOI21xp33_ASAP7_75t_L g3603 ( 
.A1(n_3462),
.A2(n_1913),
.B(n_1337),
.Y(n_3603)
);

OAI21x1_ASAP7_75t_L g3604 ( 
.A1(n_3448),
.A2(n_1013),
.B(n_1012),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3502),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3479),
.Y(n_3606)
);

OAI21x1_ASAP7_75t_L g3607 ( 
.A1(n_3434),
.A2(n_1018),
.B(n_1016),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_L g3608 ( 
.A(n_3484),
.B(n_1336),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3507),
.A2(n_1020),
.B(n_1019),
.Y(n_3609)
);

O2A1O1Ixp5_ASAP7_75t_SL g3610 ( 
.A1(n_3496),
.A2(n_1344),
.B(n_1347),
.C(n_1338),
.Y(n_3610)
);

OAI21x1_ASAP7_75t_L g3611 ( 
.A1(n_3481),
.A2(n_3465),
.B(n_3480),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3477),
.A2(n_1026),
.B(n_1023),
.Y(n_3612)
);

CKINVDCx6p67_ASAP7_75t_R g3613 ( 
.A(n_3414),
.Y(n_3613)
);

INVx5_ASAP7_75t_L g3614 ( 
.A(n_3377),
.Y(n_3614)
);

OAI21x1_ASAP7_75t_L g3615 ( 
.A1(n_3428),
.A2(n_1030),
.B(n_1029),
.Y(n_3615)
);

AO21x2_ASAP7_75t_L g3616 ( 
.A1(n_3423),
.A2(n_2182),
.B(n_1037),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_SL g3617 ( 
.A(n_3489),
.B(n_1914),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3499),
.Y(n_3618)
);

OA21x2_ASAP7_75t_L g3619 ( 
.A1(n_3408),
.A2(n_1358),
.B(n_1350),
.Y(n_3619)
);

BUFx4f_ASAP7_75t_L g3620 ( 
.A(n_3377),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3475),
.Y(n_3621)
);

CKINVDCx6p67_ASAP7_75t_R g3622 ( 
.A(n_3388),
.Y(n_3622)
);

OAI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_3575),
.A2(n_3491),
.B(n_3425),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3551),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3553),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3515),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3560),
.Y(n_3627)
);

HB1xp67_ASAP7_75t_L g3628 ( 
.A(n_3517),
.Y(n_3628)
);

OAI21x1_ASAP7_75t_SL g3629 ( 
.A1(n_3577),
.A2(n_3409),
.B(n_3469),
.Y(n_3629)
);

AOI221xp5_ASAP7_75t_L g3630 ( 
.A1(n_3603),
.A2(n_3468),
.B1(n_3430),
.B2(n_3451),
.C(n_3478),
.Y(n_3630)
);

OR2x6_ASAP7_75t_L g3631 ( 
.A(n_3533),
.B(n_3493),
.Y(n_3631)
);

OAI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_3521),
.A2(n_3498),
.B(n_3497),
.Y(n_3632)
);

AOI22xp33_ASAP7_75t_SL g3633 ( 
.A1(n_3564),
.A2(n_3458),
.B1(n_3400),
.B2(n_3431),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_3535),
.A2(n_3444),
.B1(n_3490),
.B2(n_3508),
.Y(n_3634)
);

NAND2x1p5_ASAP7_75t_L g3635 ( 
.A(n_3567),
.B(n_3614),
.Y(n_3635)
);

OAI21x1_ASAP7_75t_L g3636 ( 
.A1(n_3519),
.A2(n_3403),
.B(n_3402),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3538),
.B(n_3435),
.Y(n_3637)
);

CKINVDCx5p33_ASAP7_75t_R g3638 ( 
.A(n_3532),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3561),
.Y(n_3639)
);

BUFx3_ASAP7_75t_L g3640 ( 
.A(n_3530),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3573),
.B(n_3422),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3525),
.B(n_3429),
.Y(n_3642)
);

OAI21x1_ASAP7_75t_L g3643 ( 
.A1(n_3539),
.A2(n_3454),
.B(n_3450),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3605),
.Y(n_3644)
);

OAI22xp5_ASAP7_75t_L g3645 ( 
.A1(n_3554),
.A2(n_3547),
.B1(n_3608),
.B2(n_3540),
.Y(n_3645)
);

OAI21x1_ASAP7_75t_L g3646 ( 
.A1(n_3541),
.A2(n_3436),
.B(n_3482),
.Y(n_3646)
);

OAI21x1_ASAP7_75t_L g3647 ( 
.A1(n_3537),
.A2(n_3487),
.B(n_3488),
.Y(n_3647)
);

OAI222xp33_ASAP7_75t_L g3648 ( 
.A1(n_3546),
.A2(n_1416),
.B1(n_1390),
.B2(n_1430),
.C1(n_1398),
.C2(n_1380),
.Y(n_3648)
);

INVx1_ASAP7_75t_SL g3649 ( 
.A(n_3513),
.Y(n_3649)
);

OAI21x1_ASAP7_75t_L g3650 ( 
.A1(n_3548),
.A2(n_3476),
.B(n_3455),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3566),
.Y(n_3651)
);

NAND2x1p5_ASAP7_75t_L g3652 ( 
.A(n_3567),
.B(n_3388),
.Y(n_3652)
);

AND2x4_ASAP7_75t_L g3653 ( 
.A(n_3614),
.B(n_3433),
.Y(n_3653)
);

AND2x2_ASAP7_75t_L g3654 ( 
.A(n_3520),
.B(n_3528),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3606),
.Y(n_3655)
);

AOI221xp5_ASAP7_75t_L g3656 ( 
.A1(n_3514),
.A2(n_3529),
.B1(n_3594),
.B2(n_3585),
.C(n_3536),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3598),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3584),
.Y(n_3658)
);

BUFx6f_ASAP7_75t_L g3659 ( 
.A(n_3557),
.Y(n_3659)
);

AOI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_3516),
.A2(n_1371),
.B(n_1366),
.Y(n_3660)
);

OA21x2_ASAP7_75t_L g3661 ( 
.A1(n_3543),
.A2(n_1373),
.B(n_1372),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3586),
.Y(n_3662)
);

INVxp67_ASAP7_75t_SL g3663 ( 
.A(n_3590),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_R g3664 ( 
.A(n_3557),
.B(n_1035),
.Y(n_3664)
);

NAND2x1p5_ASAP7_75t_L g3665 ( 
.A(n_3581),
.B(n_1041),
.Y(n_3665)
);

O2A1O1Ixp33_ASAP7_75t_SL g3666 ( 
.A1(n_3589),
.A2(n_3),
.B(n_4),
.C(n_2),
.Y(n_3666)
);

INVx2_ASAP7_75t_SL g3667 ( 
.A(n_3568),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3512),
.B(n_1912),
.Y(n_3668)
);

NAND3xp33_ASAP7_75t_L g3669 ( 
.A(n_3592),
.B(n_1377),
.C(n_1375),
.Y(n_3669)
);

NOR2xp33_ASAP7_75t_SL g3670 ( 
.A(n_3558),
.B(n_1378),
.Y(n_3670)
);

A2O1A1Ixp33_ASAP7_75t_L g3671 ( 
.A1(n_3518),
.A2(n_1395),
.B(n_1408),
.C(n_1385),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3587),
.Y(n_3672)
);

CKINVDCx5p33_ASAP7_75t_R g3673 ( 
.A(n_3526),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3587),
.Y(n_3674)
);

INVx8_ASAP7_75t_L g3675 ( 
.A(n_3591),
.Y(n_3675)
);

NAND2x1p5_ASAP7_75t_L g3676 ( 
.A(n_3596),
.B(n_1042),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3602),
.Y(n_3677)
);

A2O1A1Ixp33_ASAP7_75t_L g3678 ( 
.A1(n_3571),
.A2(n_1400),
.B(n_1420),
.C(n_1388),
.Y(n_3678)
);

AOI22xp33_ASAP7_75t_L g3679 ( 
.A1(n_3564),
.A2(n_1382),
.B1(n_1383),
.B2(n_1381),
.Y(n_3679)
);

OR2x6_ASAP7_75t_L g3680 ( 
.A(n_3600),
.B(n_3612),
.Y(n_3680)
);

INVx1_ASAP7_75t_SL g3681 ( 
.A(n_3522),
.Y(n_3681)
);

BUFx2_ASAP7_75t_L g3682 ( 
.A(n_3556),
.Y(n_3682)
);

OAI21x1_ASAP7_75t_L g3683 ( 
.A1(n_3595),
.A2(n_1047),
.B(n_1045),
.Y(n_3683)
);

AOI22xp33_ASAP7_75t_L g3684 ( 
.A1(n_3621),
.A2(n_1389),
.B1(n_1391),
.B2(n_1387),
.Y(n_3684)
);

AND2x4_ASAP7_75t_L g3685 ( 
.A(n_3542),
.B(n_1048),
.Y(n_3685)
);

NAND2x1p5_ASAP7_75t_L g3686 ( 
.A(n_3620),
.B(n_1049),
.Y(n_3686)
);

OAI21xp5_ASAP7_75t_L g3687 ( 
.A1(n_3524),
.A2(n_3610),
.B(n_3582),
.Y(n_3687)
);

INVxp67_ASAP7_75t_SL g3688 ( 
.A(n_3618),
.Y(n_3688)
);

OA21x2_ASAP7_75t_L g3689 ( 
.A1(n_3604),
.A2(n_1393),
.B(n_1392),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3593),
.Y(n_3690)
);

CKINVDCx5p33_ASAP7_75t_R g3691 ( 
.A(n_3613),
.Y(n_3691)
);

AOI21x1_ASAP7_75t_L g3692 ( 
.A1(n_3559),
.A2(n_1396),
.B(n_1394),
.Y(n_3692)
);

AOI21x1_ASAP7_75t_L g3693 ( 
.A1(n_3569),
.A2(n_1401),
.B(n_1397),
.Y(n_3693)
);

INVx4_ASAP7_75t_L g3694 ( 
.A(n_3583),
.Y(n_3694)
);

AO31x2_ASAP7_75t_L g3695 ( 
.A1(n_3544),
.A2(n_6),
.A3(n_0),
.B(n_4),
.Y(n_3695)
);

OAI21x1_ASAP7_75t_L g3696 ( 
.A1(n_3611),
.A2(n_1051),
.B(n_1050),
.Y(n_3696)
);

OAI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3597),
.A2(n_1406),
.B(n_1402),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3565),
.A2(n_1415),
.B1(n_1417),
.B2(n_1407),
.Y(n_3698)
);

OR2x2_ASAP7_75t_L g3699 ( 
.A(n_3628),
.B(n_3550),
.Y(n_3699)
);

OAI21x1_ASAP7_75t_L g3700 ( 
.A1(n_3683),
.A2(n_3607),
.B(n_3609),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3657),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3663),
.Y(n_3702)
);

AOI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_3645),
.A2(n_3580),
.B(n_3616),
.Y(n_3703)
);

OAI21x1_ASAP7_75t_L g3704 ( 
.A1(n_3696),
.A2(n_3636),
.B(n_3672),
.Y(n_3704)
);

OAI21x1_ASAP7_75t_L g3705 ( 
.A1(n_3674),
.A2(n_3615),
.B(n_3552),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3624),
.Y(n_3706)
);

INVx2_ASAP7_75t_L g3707 ( 
.A(n_3655),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3654),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3625),
.Y(n_3709)
);

OAI21x1_ASAP7_75t_SL g3710 ( 
.A1(n_3629),
.A2(n_3599),
.B(n_3619),
.Y(n_3710)
);

AO31x2_ASAP7_75t_L g3711 ( 
.A1(n_3660),
.A2(n_3601),
.A3(n_3570),
.B(n_3576),
.Y(n_3711)
);

BUFx12f_ASAP7_75t_L g3712 ( 
.A(n_3638),
.Y(n_3712)
);

CKINVDCx11_ASAP7_75t_R g3713 ( 
.A(n_3675),
.Y(n_3713)
);

OAI21x1_ASAP7_75t_L g3714 ( 
.A1(n_3646),
.A2(n_3555),
.B(n_3572),
.Y(n_3714)
);

OR2x6_ASAP7_75t_L g3715 ( 
.A(n_3635),
.B(n_3583),
.Y(n_3715)
);

AO21x2_ASAP7_75t_L g3716 ( 
.A1(n_3687),
.A2(n_3523),
.B(n_3563),
.Y(n_3716)
);

HB1xp67_ASAP7_75t_L g3717 ( 
.A(n_3627),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3639),
.Y(n_3718)
);

INVx2_ASAP7_75t_SL g3719 ( 
.A(n_3640),
.Y(n_3719)
);

O2A1O1Ixp33_ASAP7_75t_L g3720 ( 
.A1(n_3648),
.A2(n_3617),
.B(n_3579),
.C(n_3588),
.Y(n_3720)
);

AOI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_3623),
.A2(n_3562),
.B(n_3545),
.Y(n_3721)
);

AO21x2_ASAP7_75t_L g3722 ( 
.A1(n_3632),
.A2(n_3549),
.B(n_3578),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3651),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3658),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3662),
.Y(n_3725)
);

NAND3xp33_ASAP7_75t_L g3726 ( 
.A(n_3656),
.B(n_3630),
.C(n_3669),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3626),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3642),
.B(n_3622),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3688),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3637),
.A2(n_3534),
.B(n_3527),
.Y(n_3730)
);

AND2x4_ASAP7_75t_L g3731 ( 
.A(n_3649),
.B(n_3531),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3644),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3682),
.Y(n_3733)
);

OAI22xp5_ASAP7_75t_L g3734 ( 
.A1(n_3633),
.A2(n_1424),
.B1(n_1427),
.B2(n_1419),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3695),
.Y(n_3735)
);

BUFx2_ASAP7_75t_L g3736 ( 
.A(n_3631),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3695),
.Y(n_3737)
);

OA21x2_ASAP7_75t_L g3738 ( 
.A1(n_3647),
.A2(n_3534),
.B(n_1429),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3681),
.Y(n_3739)
);

AOI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_3668),
.A2(n_3527),
.B(n_1431),
.Y(n_3740)
);

NOR2x1_ASAP7_75t_SL g3741 ( 
.A(n_3680),
.B(n_3574),
.Y(n_3741)
);

AOI21xp33_ASAP7_75t_SL g3742 ( 
.A1(n_3675),
.A2(n_1433),
.B(n_1428),
.Y(n_3742)
);

HB1xp67_ASAP7_75t_L g3743 ( 
.A(n_3631),
.Y(n_3743)
);

AOI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_3680),
.A2(n_1436),
.B(n_1435),
.Y(n_3744)
);

AOI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3692),
.A2(n_1442),
.B(n_1439),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3677),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3641),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_3690),
.B(n_1443),
.Y(n_3748)
);

BUFx3_ASAP7_75t_L g3749 ( 
.A(n_3659),
.Y(n_3749)
);

OAI22xp5_ASAP7_75t_L g3750 ( 
.A1(n_3634),
.A2(n_1446),
.B1(n_1448),
.B2(n_1444),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3666),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3685),
.B(n_1455),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3643),
.Y(n_3753)
);

OAI21x1_ASAP7_75t_L g3754 ( 
.A1(n_3650),
.A2(n_1055),
.B(n_1052),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3652),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3724),
.Y(n_3756)
);

OAI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3704),
.A2(n_3693),
.B(n_3689),
.Y(n_3757)
);

BUFx2_ASAP7_75t_L g3758 ( 
.A(n_3736),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3701),
.Y(n_3759)
);

HB1xp67_ASAP7_75t_L g3760 ( 
.A(n_3717),
.Y(n_3760)
);

HB1xp67_ASAP7_75t_L g3761 ( 
.A(n_3729),
.Y(n_3761)
);

INVx8_ASAP7_75t_L g3762 ( 
.A(n_3712),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3706),
.Y(n_3763)
);

BUFx2_ASAP7_75t_L g3764 ( 
.A(n_3736),
.Y(n_3764)
);

AOI22xp5_ASAP7_75t_L g3765 ( 
.A1(n_3726),
.A2(n_3679),
.B1(n_3653),
.B2(n_3686),
.Y(n_3765)
);

INVx2_ASAP7_75t_L g3766 ( 
.A(n_3707),
.Y(n_3766)
);

AO21x2_ASAP7_75t_L g3767 ( 
.A1(n_3753),
.A2(n_3671),
.B(n_3697),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3709),
.Y(n_3768)
);

OAI21x1_ASAP7_75t_L g3769 ( 
.A1(n_3714),
.A2(n_3661),
.B(n_3665),
.Y(n_3769)
);

HB1xp67_ASAP7_75t_L g3770 ( 
.A(n_3733),
.Y(n_3770)
);

OR2x2_ASAP7_75t_L g3771 ( 
.A(n_3702),
.B(n_3667),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3718),
.Y(n_3772)
);

INVx3_ASAP7_75t_L g3773 ( 
.A(n_3699),
.Y(n_3773)
);

HB1xp67_ASAP7_75t_L g3774 ( 
.A(n_3708),
.Y(n_3774)
);

OAI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_3721),
.A2(n_3678),
.B(n_3684),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3723),
.Y(n_3776)
);

BUFx3_ASAP7_75t_L g3777 ( 
.A(n_3749),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3743),
.B(n_3694),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3725),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3727),
.Y(n_3780)
);

HB1xp67_ASAP7_75t_L g3781 ( 
.A(n_3739),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3732),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3735),
.Y(n_3783)
);

BUFx3_ASAP7_75t_L g3784 ( 
.A(n_3713),
.Y(n_3784)
);

INVx3_ASAP7_75t_L g3785 ( 
.A(n_3755),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3747),
.B(n_3659),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3737),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3746),
.Y(n_3788)
);

BUFx3_ASAP7_75t_L g3789 ( 
.A(n_3731),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3722),
.Y(n_3790)
);

AO21x2_ASAP7_75t_L g3791 ( 
.A1(n_3703),
.A2(n_3664),
.B(n_3676),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3728),
.B(n_3691),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3738),
.Y(n_3793)
);

AOI21x1_ASAP7_75t_L g3794 ( 
.A1(n_3745),
.A2(n_3698),
.B(n_3670),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_3738),
.Y(n_3795)
);

AND2x4_ASAP7_75t_L g3796 ( 
.A(n_3741),
.B(n_3673),
.Y(n_3796)
);

AO21x2_ASAP7_75t_L g3797 ( 
.A1(n_3710),
.A2(n_6),
.B(n_7),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3751),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3730),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3705),
.Y(n_3800)
);

INVx4_ASAP7_75t_SL g3801 ( 
.A(n_3711),
.Y(n_3801)
);

BUFx2_ASAP7_75t_L g3802 ( 
.A(n_3715),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3719),
.B(n_7),
.Y(n_3803)
);

OAI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_3744),
.A2(n_1461),
.B(n_1456),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3715),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3716),
.Y(n_3806)
);

BUFx4f_ASAP7_75t_SL g3807 ( 
.A(n_3742),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3711),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3754),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3748),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3700),
.Y(n_3811)
);

INVx3_ASAP7_75t_L g3812 ( 
.A(n_3752),
.Y(n_3812)
);

OA21x2_ASAP7_75t_L g3813 ( 
.A1(n_3740),
.A2(n_1466),
.B(n_1464),
.Y(n_3813)
);

AO21x1_ASAP7_75t_SL g3814 ( 
.A1(n_3720),
.A2(n_8),
.B(n_9),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3775),
.A2(n_3734),
.B1(n_3750),
.B2(n_1906),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3758),
.B(n_9),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3773),
.Y(n_3817)
);

NOR3xp33_ASAP7_75t_L g3818 ( 
.A(n_3804),
.B(n_1470),
.C(n_1467),
.Y(n_3818)
);

AOI211xp5_ASAP7_75t_L g3819 ( 
.A1(n_3790),
.A2(n_1475),
.B(n_1477),
.C(n_1473),
.Y(n_3819)
);

AOI22xp33_ASAP7_75t_L g3820 ( 
.A1(n_3813),
.A2(n_1887),
.B1(n_1888),
.B2(n_1863),
.Y(n_3820)
);

OAI22xp5_ASAP7_75t_L g3821 ( 
.A1(n_3765),
.A2(n_1478),
.B1(n_1479),
.B2(n_1476),
.Y(n_3821)
);

NAND3xp33_ASAP7_75t_L g3822 ( 
.A(n_3813),
.B(n_1484),
.C(n_1482),
.Y(n_3822)
);

AOI221xp5_ASAP7_75t_L g3823 ( 
.A1(n_3810),
.A2(n_1489),
.B1(n_1492),
.B2(n_1486),
.C(n_1485),
.Y(n_3823)
);

AOI21xp5_ASAP7_75t_L g3824 ( 
.A1(n_3791),
.A2(n_1496),
.B(n_1495),
.Y(n_3824)
);

OAI22xp5_ASAP7_75t_L g3825 ( 
.A1(n_3805),
.A2(n_1505),
.B1(n_1509),
.B2(n_1501),
.Y(n_3825)
);

OAI22xp33_ASAP7_75t_L g3826 ( 
.A1(n_3812),
.A2(n_1513),
.B1(n_1515),
.B2(n_1510),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_R g3827 ( 
.A(n_3784),
.B(n_10),
.Y(n_3827)
);

INVx4_ASAP7_75t_L g3828 ( 
.A(n_3762),
.Y(n_3828)
);

INVxp67_ASAP7_75t_SL g3829 ( 
.A(n_3760),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3781),
.B(n_1517),
.Y(n_3830)
);

OAI22xp33_ASAP7_75t_L g3831 ( 
.A1(n_3812),
.A2(n_1524),
.B1(n_1526),
.B2(n_1519),
.Y(n_3831)
);

OAI22xp33_ASAP7_75t_L g3832 ( 
.A1(n_3764),
.A2(n_3802),
.B1(n_3773),
.B2(n_3794),
.Y(n_3832)
);

AOI221xp5_ASAP7_75t_L g3833 ( 
.A1(n_3808),
.A2(n_1536),
.B1(n_1537),
.B2(n_1532),
.C(n_1531),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3763),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3763),
.Y(n_3835)
);

OAI22xp5_ASAP7_75t_L g3836 ( 
.A1(n_3789),
.A2(n_1542),
.B1(n_1545),
.B2(n_1541),
.Y(n_3836)
);

OAI22xp5_ASAP7_75t_L g3837 ( 
.A1(n_3798),
.A2(n_1547),
.B1(n_1548),
.B2(n_1546),
.Y(n_3837)
);

OAI22xp5_ASAP7_75t_L g3838 ( 
.A1(n_3796),
.A2(n_1553),
.B1(n_1554),
.B2(n_1551),
.Y(n_3838)
);

HB1xp67_ASAP7_75t_L g3839 ( 
.A(n_3761),
.Y(n_3839)
);

CKINVDCx5p33_ASAP7_75t_R g3840 ( 
.A(n_3762),
.Y(n_3840)
);

INVx2_ASAP7_75t_L g3841 ( 
.A(n_3768),
.Y(n_3841)
);

INVxp67_ASAP7_75t_L g3842 ( 
.A(n_3770),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3772),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3772),
.Y(n_3844)
);

AOI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3767),
.A2(n_1556),
.B1(n_1557),
.B2(n_1555),
.Y(n_3845)
);

AOI22xp33_ASAP7_75t_SL g3846 ( 
.A1(n_3797),
.A2(n_1559),
.B1(n_1560),
.B2(n_1558),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3776),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3782),
.B(n_1562),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3817),
.B(n_3778),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3829),
.B(n_3788),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3834),
.Y(n_3851)
);

INVx3_ASAP7_75t_SL g3852 ( 
.A(n_3840),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3835),
.Y(n_3853)
);

OR2x2_ASAP7_75t_L g3854 ( 
.A(n_3839),
.B(n_3774),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3842),
.B(n_3796),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3844),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3847),
.B(n_3779),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3843),
.Y(n_3858)
);

AOI22xp33_ASAP7_75t_L g3859 ( 
.A1(n_3818),
.A2(n_3814),
.B1(n_3806),
.B2(n_3809),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3841),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3828),
.B(n_3785),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3816),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3848),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3830),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3828),
.B(n_3785),
.Y(n_3865)
);

NOR2xp33_ASAP7_75t_L g3866 ( 
.A(n_3838),
.B(n_3792),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3827),
.B(n_3786),
.Y(n_3867)
);

OR2x2_ASAP7_75t_L g3868 ( 
.A(n_3832),
.B(n_3799),
.Y(n_3868)
);

HB1xp67_ASAP7_75t_L g3869 ( 
.A(n_3845),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3824),
.B(n_3801),
.Y(n_3870)
);

INVx1_ASAP7_75t_SL g3871 ( 
.A(n_3846),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3821),
.B(n_3801),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3822),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3836),
.Y(n_3874)
);

NOR2xp67_ASAP7_75t_L g3875 ( 
.A(n_3820),
.B(n_3811),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3819),
.B(n_3777),
.Y(n_3876)
);

OAI222xp33_ASAP7_75t_L g3877 ( 
.A1(n_3815),
.A2(n_3794),
.B1(n_3771),
.B2(n_3809),
.C1(n_3793),
.C2(n_3795),
.Y(n_3877)
);

INVxp67_ASAP7_75t_SL g3878 ( 
.A(n_3826),
.Y(n_3878)
);

OR2x2_ASAP7_75t_L g3879 ( 
.A(n_3825),
.B(n_3756),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3837),
.B(n_3759),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3831),
.B(n_3780),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3851),
.Y(n_3882)
);

OR2x2_ASAP7_75t_L g3883 ( 
.A(n_3854),
.B(n_3766),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3855),
.B(n_3783),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3861),
.B(n_3787),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3865),
.B(n_3803),
.Y(n_3886)
);

BUFx2_ASAP7_75t_L g3887 ( 
.A(n_3867),
.Y(n_3887)
);

BUFx2_ASAP7_75t_L g3888 ( 
.A(n_3870),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3851),
.Y(n_3889)
);

NAND3xp33_ASAP7_75t_L g3890 ( 
.A(n_3875),
.B(n_3833),
.C(n_3823),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3858),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3863),
.B(n_3793),
.Y(n_3892)
);

OAI21xp5_ASAP7_75t_SL g3893 ( 
.A1(n_3871),
.A2(n_3807),
.B(n_3811),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3849),
.B(n_3769),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3862),
.B(n_3800),
.Y(n_3895)
);

OAI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3875),
.A2(n_1565),
.B1(n_1566),
.B2(n_1564),
.Y(n_3896)
);

AND2x2_ASAP7_75t_L g3897 ( 
.A(n_3864),
.B(n_3757),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3881),
.B(n_1567),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3853),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3853),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3857),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_3860),
.B(n_3872),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3850),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3860),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3856),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3880),
.B(n_1569),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3868),
.B(n_12),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3852),
.B(n_14),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3873),
.B(n_1570),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3879),
.Y(n_3910)
);

OR2x2_ASAP7_75t_L g3911 ( 
.A(n_3878),
.B(n_14),
.Y(n_3911)
);

AOI221xp5_ASAP7_75t_L g3912 ( 
.A1(n_3869),
.A2(n_1576),
.B1(n_1577),
.B2(n_1575),
.C(n_1573),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3876),
.B(n_15),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3874),
.B(n_15),
.Y(n_3914)
);

AND2x2_ASAP7_75t_L g3915 ( 
.A(n_3866),
.B(n_3859),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3871),
.B(n_16),
.Y(n_3916)
);

INVx2_ASAP7_75t_L g3917 ( 
.A(n_3887),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3907),
.B(n_1581),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3888),
.B(n_3877),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3902),
.B(n_16),
.Y(n_3920)
);

INVx2_ASAP7_75t_SL g3921 ( 
.A(n_3886),
.Y(n_3921)
);

NOR3xp33_ASAP7_75t_SL g3922 ( 
.A(n_3893),
.B(n_1583),
.C(n_1582),
.Y(n_3922)
);

OR2x2_ASAP7_75t_L g3923 ( 
.A(n_3910),
.B(n_17),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3910),
.B(n_1584),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3882),
.Y(n_3925)
);

OAI321xp33_ASAP7_75t_L g3926 ( 
.A1(n_3890),
.A2(n_22),
.A3(n_25),
.B1(n_18),
.B2(n_19),
.C(n_24),
.Y(n_3926)
);

AOI22xp5_ASAP7_75t_L g3927 ( 
.A1(n_3915),
.A2(n_1589),
.B1(n_1594),
.B2(n_1585),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3903),
.B(n_1597),
.Y(n_3928)
);

BUFx3_ASAP7_75t_L g3929 ( 
.A(n_3908),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3901),
.B(n_1598),
.Y(n_3930)
);

INVxp67_ASAP7_75t_L g3931 ( 
.A(n_3911),
.Y(n_3931)
);

INVx2_ASAP7_75t_SL g3932 ( 
.A(n_3884),
.Y(n_3932)
);

AND2x2_ASAP7_75t_L g3933 ( 
.A(n_3885),
.B(n_19),
.Y(n_3933)
);

OAI31xp33_ASAP7_75t_L g3934 ( 
.A1(n_3896),
.A2(n_26),
.A3(n_22),
.B(n_24),
.Y(n_3934)
);

AOI22xp5_ASAP7_75t_L g3935 ( 
.A1(n_3916),
.A2(n_1601),
.B1(n_1602),
.B2(n_1600),
.Y(n_3935)
);

OR2x2_ASAP7_75t_L g3936 ( 
.A(n_3892),
.B(n_26),
.Y(n_3936)
);

HB1xp67_ASAP7_75t_L g3937 ( 
.A(n_3882),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3889),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3883),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3899),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3900),
.Y(n_3941)
);

AND2x2_ASAP7_75t_SL g3942 ( 
.A(n_3913),
.B(n_27),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3894),
.B(n_27),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3897),
.B(n_28),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3891),
.B(n_3895),
.Y(n_3945)
);

INVx3_ASAP7_75t_L g3946 ( 
.A(n_3905),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3904),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_SL g3948 ( 
.A(n_3898),
.B(n_1606),
.Y(n_3948)
);

HB1xp67_ASAP7_75t_L g3949 ( 
.A(n_3905),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3937),
.Y(n_3950)
);

INVx3_ASAP7_75t_L g3951 ( 
.A(n_3929),
.Y(n_3951)
);

INVx4_ASAP7_75t_L g3952 ( 
.A(n_3923),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3917),
.B(n_3914),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3925),
.Y(n_3954)
);

INVx1_ASAP7_75t_SL g3955 ( 
.A(n_3942),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3925),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3931),
.B(n_3906),
.Y(n_3957)
);

AOI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3948),
.A2(n_3909),
.B(n_3912),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3927),
.B(n_3920),
.Y(n_3959)
);

OR2x2_ASAP7_75t_L g3960 ( 
.A(n_3939),
.B(n_29),
.Y(n_3960)
);

NAND3xp33_ASAP7_75t_L g3961 ( 
.A(n_3934),
.B(n_1608),
.C(n_1607),
.Y(n_3961)
);

AND2x2_ASAP7_75t_L g3962 ( 
.A(n_3921),
.B(n_30),
.Y(n_3962)
);

OR2x2_ASAP7_75t_L g3963 ( 
.A(n_3936),
.B(n_30),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3932),
.B(n_31),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3943),
.B(n_31),
.Y(n_3965)
);

OR2x2_ASAP7_75t_L g3966 ( 
.A(n_3924),
.B(n_32),
.Y(n_3966)
);

AND2x2_ASAP7_75t_L g3967 ( 
.A(n_3944),
.B(n_32),
.Y(n_3967)
);

INVx1_ASAP7_75t_SL g3968 ( 
.A(n_3933),
.Y(n_3968)
);

OR2x2_ASAP7_75t_L g3969 ( 
.A(n_3919),
.B(n_33),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3945),
.B(n_33),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3928),
.B(n_1611),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3949),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3940),
.Y(n_3973)
);

INVx1_ASAP7_75t_SL g3974 ( 
.A(n_3918),
.Y(n_3974)
);

NOR2x1_ASAP7_75t_L g3975 ( 
.A(n_3946),
.B(n_34),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3940),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3922),
.B(n_35),
.Y(n_3977)
);

NOR2x1_ASAP7_75t_L g3978 ( 
.A(n_3946),
.B(n_36),
.Y(n_3978)
);

OR2x2_ASAP7_75t_L g3979 ( 
.A(n_3930),
.B(n_37),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3938),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3947),
.B(n_38),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_3935),
.B(n_3941),
.Y(n_3982)
);

HB1xp67_ASAP7_75t_L g3983 ( 
.A(n_3926),
.Y(n_3983)
);

NAND4xp25_ASAP7_75t_L g3984 ( 
.A(n_3917),
.B(n_1917),
.C(n_1915),
.D(n_1613),
.Y(n_3984)
);

OR2x2_ASAP7_75t_L g3985 ( 
.A(n_3931),
.B(n_38),
.Y(n_3985)
);

AOI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3919),
.A2(n_1615),
.B1(n_1619),
.B2(n_1612),
.Y(n_3986)
);

INVx3_ASAP7_75t_L g3987 ( 
.A(n_3929),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3929),
.Y(n_3988)
);

OR2x2_ASAP7_75t_L g3989 ( 
.A(n_3931),
.B(n_39),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3937),
.Y(n_3990)
);

AND2x4_ASAP7_75t_L g3991 ( 
.A(n_3929),
.B(n_42),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3929),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3937),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3937),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3955),
.B(n_1620),
.Y(n_3995)
);

AND2x2_ASAP7_75t_SL g3996 ( 
.A(n_3983),
.B(n_43),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3954),
.Y(n_3997)
);

AND2x4_ASAP7_75t_L g3998 ( 
.A(n_3951),
.B(n_44),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3968),
.B(n_1621),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3952),
.B(n_1624),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3952),
.B(n_1625),
.Y(n_4001)
);

AND2x2_ASAP7_75t_L g4002 ( 
.A(n_3987),
.B(n_45),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3956),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3988),
.Y(n_4004)
);

OAI22xp33_ASAP7_75t_L g4005 ( 
.A1(n_3969),
.A2(n_1652),
.B1(n_1665),
.B2(n_1642),
.Y(n_4005)
);

INVx1_ASAP7_75t_SL g4006 ( 
.A(n_3975),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_3953),
.B(n_3978),
.Y(n_4007)
);

OR2x2_ASAP7_75t_L g4008 ( 
.A(n_3957),
.B(n_46),
.Y(n_4008)
);

NOR2xp33_ASAP7_75t_L g4009 ( 
.A(n_3992),
.B(n_1626),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3974),
.B(n_1627),
.Y(n_4010)
);

OR2x2_ASAP7_75t_L g4011 ( 
.A(n_3982),
.B(n_3960),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3973),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3986),
.B(n_1628),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3970),
.B(n_1631),
.Y(n_4014)
);

AND2x2_ASAP7_75t_L g4015 ( 
.A(n_3962),
.B(n_46),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3959),
.B(n_1632),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3967),
.B(n_3965),
.Y(n_4017)
);

BUFx2_ASAP7_75t_L g4018 ( 
.A(n_3972),
.Y(n_4018)
);

NAND2x1p5_ASAP7_75t_L g4019 ( 
.A(n_3991),
.B(n_48),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3964),
.B(n_47),
.Y(n_4020)
);

OR2x6_ASAP7_75t_L g4021 ( 
.A(n_3991),
.B(n_48),
.Y(n_4021)
);

OR2x2_ASAP7_75t_L g4022 ( 
.A(n_3950),
.B(n_49),
.Y(n_4022)
);

OR2x2_ASAP7_75t_L g4023 ( 
.A(n_3990),
.B(n_49),
.Y(n_4023)
);

INVx1_ASAP7_75t_SL g4024 ( 
.A(n_3963),
.Y(n_4024)
);

INVx1_ASAP7_75t_SL g4025 ( 
.A(n_3985),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3981),
.B(n_50),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3976),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3989),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3993),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3958),
.B(n_3994),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3979),
.B(n_51),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3980),
.Y(n_4032)
);

HB1xp67_ASAP7_75t_L g4033 ( 
.A(n_3966),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3971),
.Y(n_4034)
);

INVx2_ASAP7_75t_SL g4035 ( 
.A(n_3977),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3961),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3984),
.B(n_1635),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3954),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3955),
.B(n_1638),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3955),
.B(n_52),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3955),
.B(n_53),
.Y(n_4041)
);

INVxp67_ASAP7_75t_L g4042 ( 
.A(n_3975),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3954),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3955),
.B(n_1643),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_3955),
.B(n_53),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3954),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3954),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3955),
.B(n_1644),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3955),
.B(n_1646),
.Y(n_4049)
);

INVxp67_ASAP7_75t_SL g4050 ( 
.A(n_3975),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3955),
.B(n_55),
.Y(n_4051)
);

OR2x2_ASAP7_75t_L g4052 ( 
.A(n_3969),
.B(n_58),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3955),
.B(n_58),
.Y(n_4053)
);

INVx2_ASAP7_75t_L g4054 ( 
.A(n_3951),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_3955),
.B(n_59),
.Y(n_4055)
);

HB1xp67_ASAP7_75t_L g4056 ( 
.A(n_3955),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3955),
.B(n_59),
.Y(n_4057)
);

NAND2x1_ASAP7_75t_L g4058 ( 
.A(n_3952),
.B(n_60),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_3951),
.Y(n_4059)
);

NOR2xp33_ASAP7_75t_SL g4060 ( 
.A(n_4006),
.B(n_1650),
.Y(n_4060)
);

OAI22xp5_ASAP7_75t_L g4061 ( 
.A1(n_4050),
.A2(n_1648),
.B1(n_1651),
.B2(n_1647),
.Y(n_4061)
);

NAND3xp33_ASAP7_75t_L g4062 ( 
.A(n_4042),
.B(n_1655),
.C(n_1653),
.Y(n_4062)
);

AND2x2_ASAP7_75t_L g4063 ( 
.A(n_4056),
.B(n_1656),
.Y(n_4063)
);

OAI211xp5_ASAP7_75t_L g4064 ( 
.A1(n_4030),
.A2(n_1661),
.B(n_1663),
.C(n_1659),
.Y(n_4064)
);

AOI31xp33_ASAP7_75t_L g4065 ( 
.A1(n_4019),
.A2(n_1669),
.A3(n_1672),
.B(n_1664),
.Y(n_4065)
);

NOR2x1_ASAP7_75t_L g4066 ( 
.A(n_4058),
.B(n_60),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_SL g4067 ( 
.A1(n_3996),
.A2(n_1678),
.B1(n_1680),
.B2(n_1675),
.Y(n_4067)
);

AOI22xp5_ASAP7_75t_L g4068 ( 
.A1(n_4035),
.A2(n_1684),
.B1(n_1685),
.B2(n_1682),
.Y(n_4068)
);

OAI31xp33_ASAP7_75t_L g4069 ( 
.A1(n_4007),
.A2(n_64),
.A3(n_61),
.B(n_62),
.Y(n_4069)
);

OAI31xp33_ASAP7_75t_L g4070 ( 
.A1(n_4018),
.A2(n_65),
.A3(n_62),
.B(n_64),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_4040),
.Y(n_4071)
);

OAI32xp33_ASAP7_75t_L g4072 ( 
.A1(n_4011),
.A2(n_1691),
.A3(n_1693),
.B1(n_1690),
.B2(n_1688),
.Y(n_4072)
);

OAI22xp5_ASAP7_75t_L g4073 ( 
.A1(n_4054),
.A2(n_1696),
.B1(n_1697),
.B2(n_1695),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_4041),
.Y(n_4074)
);

OR2x2_ASAP7_75t_L g4075 ( 
.A(n_4024),
.B(n_65),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4045),
.Y(n_4076)
);

NOR2xp33_ASAP7_75t_L g4077 ( 
.A(n_4059),
.B(n_1698),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_4058),
.Y(n_4078)
);

OAI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_4017),
.A2(n_1702),
.B(n_1699),
.Y(n_4079)
);

OAI21xp33_ASAP7_75t_L g4080 ( 
.A1(n_4004),
.A2(n_1708),
.B(n_1704),
.Y(n_4080)
);

OAI22xp33_ASAP7_75t_L g4081 ( 
.A1(n_4025),
.A2(n_1710),
.B1(n_1713),
.B2(n_1709),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_4051),
.B(n_1715),
.Y(n_4082)
);

AOI22xp33_ASAP7_75t_L g4083 ( 
.A1(n_4034),
.A2(n_4028),
.B1(n_4033),
.B2(n_4036),
.Y(n_4083)
);

AOI32xp33_ASAP7_75t_L g4084 ( 
.A1(n_4053),
.A2(n_1721),
.A3(n_1722),
.B1(n_1719),
.B2(n_1718),
.Y(n_4084)
);

INVxp67_ASAP7_75t_L g4085 ( 
.A(n_4055),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_4057),
.Y(n_4086)
);

AND3x1_ASAP7_75t_L g4087 ( 
.A(n_4029),
.B(n_68),
.C(n_69),
.Y(n_4087)
);

AND2x4_ASAP7_75t_L g4088 ( 
.A(n_3998),
.B(n_69),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_4022),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_4005),
.B(n_4031),
.Y(n_4090)
);

OAI22xp5_ASAP7_75t_L g4091 ( 
.A1(n_4008),
.A2(n_1726),
.B1(n_1729),
.B2(n_1725),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_4021),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_4002),
.B(n_1733),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4023),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_4015),
.B(n_4020),
.Y(n_4095)
);

HB1xp67_ASAP7_75t_L g4096 ( 
.A(n_4021),
.Y(n_4096)
);

INVx2_ASAP7_75t_L g4097 ( 
.A(n_3998),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_4052),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3997),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_4003),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_4026),
.Y(n_4101)
);

OR2x2_ASAP7_75t_L g4102 ( 
.A(n_3995),
.B(n_68),
.Y(n_4102)
);

OAI222xp33_ASAP7_75t_L g4103 ( 
.A1(n_4032),
.A2(n_1742),
.B1(n_1739),
.B2(n_1743),
.C1(n_1741),
.C2(n_1737),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4038),
.Y(n_4104)
);

AOI21xp33_ASAP7_75t_L g4105 ( 
.A1(n_4000),
.A2(n_1746),
.B(n_1745),
.Y(n_4105)
);

OAI211xp5_ASAP7_75t_L g4106 ( 
.A1(n_4012),
.A2(n_1749),
.B(n_1751),
.C(n_1747),
.Y(n_4106)
);

OAI21xp33_ASAP7_75t_L g4107 ( 
.A1(n_4027),
.A2(n_1756),
.B(n_1755),
.Y(n_4107)
);

AND2x4_ASAP7_75t_L g4108 ( 
.A(n_4043),
.B(n_71),
.Y(n_4108)
);

INVx2_ASAP7_75t_SL g4109 ( 
.A(n_4046),
.Y(n_4109)
);

OAI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_4016),
.A2(n_1761),
.B(n_1759),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_4039),
.B(n_1764),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_4009),
.B(n_1770),
.Y(n_4112)
);

NAND2x1p5_ASAP7_75t_L g4113 ( 
.A(n_4047),
.B(n_70),
.Y(n_4113)
);

INVxp33_ASAP7_75t_L g4114 ( 
.A(n_4010),
.Y(n_4114)
);

AOI21x1_ASAP7_75t_L g4115 ( 
.A1(n_4044),
.A2(n_72),
.B(n_73),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3999),
.Y(n_4116)
);

INVx2_ASAP7_75t_SL g4117 ( 
.A(n_4001),
.Y(n_4117)
);

AND2x2_ASAP7_75t_L g4118 ( 
.A(n_4014),
.B(n_1773),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_4048),
.B(n_1781),
.Y(n_4119)
);

OR2x2_ASAP7_75t_L g4120 ( 
.A(n_4049),
.B(n_74),
.Y(n_4120)
);

NAND2xp33_ASAP7_75t_L g4121 ( 
.A(n_4037),
.B(n_1782),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4013),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4056),
.Y(n_4123)
);

AOI22xp5_ASAP7_75t_L g4124 ( 
.A1(n_3996),
.A2(n_1794),
.B1(n_1795),
.B2(n_1787),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4056),
.Y(n_4125)
);

OAI21xp5_ASAP7_75t_L g4126 ( 
.A1(n_4042),
.A2(n_1800),
.B(n_1798),
.Y(n_4126)
);

NAND2x1_ASAP7_75t_L g4127 ( 
.A(n_4018),
.B(n_74),
.Y(n_4127)
);

INVx1_ASAP7_75t_SL g4128 ( 
.A(n_4006),
.Y(n_4128)
);

NAND3xp33_ASAP7_75t_L g4129 ( 
.A(n_4042),
.B(n_1802),
.C(n_1801),
.Y(n_4129)
);

INVxp67_ASAP7_75t_L g4130 ( 
.A(n_4056),
.Y(n_4130)
);

AND2x2_ASAP7_75t_L g4131 ( 
.A(n_4056),
.B(n_1803),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_4056),
.Y(n_4132)
);

AOI21xp33_ASAP7_75t_L g4133 ( 
.A1(n_4056),
.A2(n_1805),
.B(n_1804),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_4019),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4056),
.B(n_1812),
.Y(n_4135)
);

OAI22xp5_ASAP7_75t_L g4136 ( 
.A1(n_4050),
.A2(n_1817),
.B1(n_1821),
.B2(n_1815),
.Y(n_4136)
);

OAI22xp33_ASAP7_75t_L g4137 ( 
.A1(n_4050),
.A2(n_1823),
.B1(n_1824),
.B2(n_1822),
.Y(n_4137)
);

OAI22xp5_ASAP7_75t_L g4138 ( 
.A1(n_4050),
.A2(n_1827),
.B1(n_1828),
.B2(n_1826),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4056),
.Y(n_4139)
);

OR2x2_ASAP7_75t_L g4140 ( 
.A(n_4056),
.B(n_75),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4056),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_4019),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4056),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4056),
.Y(n_4144)
);

NOR2x1_ASAP7_75t_L g4145 ( 
.A(n_4058),
.B(n_75),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_4019),
.Y(n_4146)
);

AOI221xp5_ASAP7_75t_L g4147 ( 
.A1(n_4130),
.A2(n_1838),
.B1(n_1839),
.B2(n_1835),
.C(n_1834),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_4096),
.Y(n_4148)
);

OR2x2_ASAP7_75t_L g4149 ( 
.A(n_4128),
.B(n_76),
.Y(n_4149)
);

NOR2x1_ASAP7_75t_L g4150 ( 
.A(n_4066),
.B(n_77),
.Y(n_4150)
);

A2O1A1Ixp33_ASAP7_75t_L g4151 ( 
.A1(n_4069),
.A2(n_1844),
.B(n_1845),
.C(n_1842),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_4123),
.Y(n_4152)
);

OAI22xp5_ASAP7_75t_L g4153 ( 
.A1(n_4083),
.A2(n_1848),
.B1(n_1849),
.B2(n_1847),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4125),
.Y(n_4154)
);

AOI22xp33_ASAP7_75t_L g4155 ( 
.A1(n_4132),
.A2(n_1852),
.B1(n_1892),
.B2(n_1851),
.Y(n_4155)
);

AOI22xp5_ASAP7_75t_L g4156 ( 
.A1(n_4139),
.A2(n_1855),
.B1(n_1859),
.B2(n_1858),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_4078),
.B(n_1860),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_4092),
.B(n_1889),
.Y(n_4158)
);

O2A1O1Ixp33_ASAP7_75t_L g4159 ( 
.A1(n_4127),
.A2(n_81),
.B(n_78),
.C(n_80),
.Y(n_4159)
);

O2A1O1Ixp33_ASAP7_75t_L g4160 ( 
.A1(n_4145),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_4160)
);

OAI322xp33_ASAP7_75t_L g4161 ( 
.A1(n_4141),
.A2(n_1897),
.A3(n_1891),
.B1(n_1898),
.B2(n_1901),
.C1(n_1895),
.C2(n_1890),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4143),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4144),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4097),
.B(n_1907),
.Y(n_4164)
);

OAI21xp5_ASAP7_75t_L g4165 ( 
.A1(n_4085),
.A2(n_1908),
.B(n_83),
.Y(n_4165)
);

INVx1_ASAP7_75t_SL g4166 ( 
.A(n_4140),
.Y(n_4166)
);

AND2x2_ASAP7_75t_L g4167 ( 
.A(n_4095),
.B(n_84),
.Y(n_4167)
);

INVx3_ASAP7_75t_SL g4168 ( 
.A(n_4088),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_4134),
.B(n_86),
.Y(n_4169)
);

NAND4xp25_ASAP7_75t_SL g4170 ( 
.A(n_4071),
.B(n_88),
.C(n_86),
.D(n_87),
.Y(n_4170)
);

INVxp67_ASAP7_75t_SL g4171 ( 
.A(n_4113),
.Y(n_4171)
);

OAI31xp33_ASAP7_75t_L g4172 ( 
.A1(n_4060),
.A2(n_90),
.A3(n_88),
.B(n_89),
.Y(n_4172)
);

OAI21xp5_ASAP7_75t_L g4173 ( 
.A1(n_4067),
.A2(n_4146),
.B(n_4142),
.Y(n_4173)
);

A2O1A1Ixp33_ASAP7_75t_L g4174 ( 
.A1(n_4070),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_4174)
);

AND2x2_ASAP7_75t_L g4175 ( 
.A(n_4074),
.B(n_91),
.Y(n_4175)
);

AND2x2_ASAP7_75t_L g4176 ( 
.A(n_4076),
.B(n_92),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4086),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_4101),
.B(n_93),
.Y(n_4178)
);

AOI21xp5_ASAP7_75t_L g4179 ( 
.A1(n_4065),
.A2(n_93),
.B(n_94),
.Y(n_4179)
);

INVx2_ASAP7_75t_L g4180 ( 
.A(n_4088),
.Y(n_4180)
);

OAI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_4087),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_4181)
);

OR2x2_ASAP7_75t_L g4182 ( 
.A(n_4089),
.B(n_96),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4075),
.Y(n_4183)
);

OAI221xp5_ASAP7_75t_L g4184 ( 
.A1(n_4094),
.A2(n_100),
.B1(n_97),
.B2(n_99),
.C(n_101),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4108),
.Y(n_4185)
);

OAI31xp33_ASAP7_75t_L g4186 ( 
.A1(n_4064),
.A2(n_102),
.A3(n_97),
.B(n_99),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4108),
.Y(n_4187)
);

OA21x2_ASAP7_75t_L g4188 ( 
.A1(n_4133),
.A2(n_102),
.B(n_103),
.Y(n_4188)
);

OAI21xp33_ASAP7_75t_L g4189 ( 
.A1(n_4090),
.A2(n_103),
.B(n_104),
.Y(n_4189)
);

OAI22xp5_ASAP7_75t_L g4190 ( 
.A1(n_4124),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_4190)
);

AND2x2_ASAP7_75t_L g4191 ( 
.A(n_4098),
.B(n_105),
.Y(n_4191)
);

AOI322xp5_ASAP7_75t_L g4192 ( 
.A1(n_4109),
.A2(n_112),
.A3(n_111),
.B1(n_109),
.B2(n_107),
.C1(n_108),
.C2(n_110),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_4063),
.B(n_108),
.Y(n_4193)
);

HB1xp67_ASAP7_75t_L g4194 ( 
.A(n_4115),
.Y(n_4194)
);

OAI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_4116),
.A2(n_113),
.B1(n_110),
.B2(n_111),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4102),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4120),
.Y(n_4197)
);

NOR2xp33_ASAP7_75t_L g4198 ( 
.A(n_4114),
.B(n_114),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4099),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4100),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4104),
.Y(n_4201)
);

OAI322xp33_ASAP7_75t_L g4202 ( 
.A1(n_4135),
.A2(n_119),
.A3(n_118),
.B1(n_116),
.B2(n_114),
.C1(n_115),
.C2(n_117),
.Y(n_4202)
);

INVx1_ASAP7_75t_SL g4203 ( 
.A(n_4131),
.Y(n_4203)
);

NOR2xp33_ASAP7_75t_L g4204 ( 
.A(n_4082),
.B(n_117),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_4117),
.Y(n_4205)
);

AND2x2_ASAP7_75t_L g4206 ( 
.A(n_4122),
.B(n_121),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_4093),
.Y(n_4207)
);

INVxp67_ASAP7_75t_L g4208 ( 
.A(n_4077),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_L g4209 ( 
.A(n_4103),
.B(n_122),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4118),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4068),
.Y(n_4211)
);

CKINVDCx14_ASAP7_75t_R g4212 ( 
.A(n_4111),
.Y(n_4212)
);

OAI22xp5_ASAP7_75t_L g4213 ( 
.A1(n_4062),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_4213)
);

OR2x2_ASAP7_75t_L g4214 ( 
.A(n_4091),
.B(n_4129),
.Y(n_4214)
);

AOI22xp33_ASAP7_75t_L g4215 ( 
.A1(n_4080),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_4215)
);

BUFx3_ASAP7_75t_L g4216 ( 
.A(n_4119),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4084),
.B(n_125),
.Y(n_4217)
);

O2A1O1Ixp33_ASAP7_75t_SL g4218 ( 
.A1(n_4137),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_4218)
);

HB1xp67_ASAP7_75t_L g4219 ( 
.A(n_4126),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4073),
.Y(n_4220)
);

AOI22xp33_ASAP7_75t_L g4221 ( 
.A1(n_4107),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_4079),
.B(n_131),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4081),
.B(n_133),
.Y(n_4223)
);

AOI322xp5_ASAP7_75t_L g4224 ( 
.A1(n_4112),
.A2(n_139),
.A3(n_138),
.B1(n_135),
.B2(n_133),
.C1(n_134),
.C2(n_136),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4061),
.Y(n_4225)
);

OR2x2_ASAP7_75t_L g4226 ( 
.A(n_4136),
.B(n_134),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_4138),
.Y(n_4227)
);

AOI22xp5_ASAP7_75t_L g4228 ( 
.A1(n_4121),
.A2(n_139),
.B1(n_135),
.B2(n_138),
.Y(n_4228)
);

AOI21xp33_ASAP7_75t_SL g4229 ( 
.A1(n_4106),
.A2(n_140),
.B(n_141),
.Y(n_4229)
);

OAI31xp33_ASAP7_75t_L g4230 ( 
.A1(n_4105),
.A2(n_142),
.A3(n_140),
.B(n_141),
.Y(n_4230)
);

OAI22xp5_ASAP7_75t_L g4231 ( 
.A1(n_4110),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_4231)
);

OAI222xp33_ASAP7_75t_L g4232 ( 
.A1(n_4072),
.A2(n_145),
.B1(n_149),
.B2(n_143),
.C1(n_144),
.C2(n_146),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4096),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_4128),
.B(n_145),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_4128),
.B(n_146),
.Y(n_4235)
);

INVxp67_ASAP7_75t_L g4236 ( 
.A(n_4066),
.Y(n_4236)
);

OR2x2_ASAP7_75t_L g4237 ( 
.A(n_4128),
.B(n_150),
.Y(n_4237)
);

OAI22xp33_ASAP7_75t_L g4238 ( 
.A1(n_4128),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4096),
.Y(n_4239)
);

O2A1O1Ixp5_ASAP7_75t_L g4240 ( 
.A1(n_4078),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_4078),
.Y(n_4241)
);

AOI22xp5_ASAP7_75t_L g4242 ( 
.A1(n_4128),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_4242)
);

AND2x2_ASAP7_75t_L g4243 ( 
.A(n_4128),
.B(n_156),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4128),
.B(n_158),
.Y(n_4244)
);

AOI221xp5_ASAP7_75t_L g4245 ( 
.A1(n_4130),
.A2(n_183),
.B1(n_192),
.B2(n_171),
.C(n_159),
.Y(n_4245)
);

AOI221xp5_ASAP7_75t_L g4246 ( 
.A1(n_4130),
.A2(n_183),
.B1(n_192),
.B2(n_171),
.C(n_159),
.Y(n_4246)
);

AOI321xp33_ASAP7_75t_L g4247 ( 
.A1(n_4123),
.A2(n_163),
.A3(n_168),
.B1(n_160),
.B2(n_161),
.C(n_165),
.Y(n_4247)
);

INVxp67_ASAP7_75t_SL g4248 ( 
.A(n_4066),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4096),
.Y(n_4249)
);

O2A1O1Ixp33_ASAP7_75t_L g4250 ( 
.A1(n_4069),
.A2(n_163),
.B(n_160),
.C(n_161),
.Y(n_4250)
);

NOR4xp25_ASAP7_75t_L g4251 ( 
.A(n_4128),
.B(n_172),
.C(n_169),
.D(n_170),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_4128),
.B(n_169),
.Y(n_4252)
);

INVxp67_ASAP7_75t_L g4253 ( 
.A(n_4066),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4128),
.B(n_170),
.Y(n_4254)
);

NOR2xp33_ASAP7_75t_L g4255 ( 
.A(n_4128),
.B(n_173),
.Y(n_4255)
);

OAI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_4066),
.A2(n_173),
.B(n_174),
.Y(n_4256)
);

OAI21xp5_ASAP7_75t_L g4257 ( 
.A1(n_4066),
.A2(n_174),
.B(n_176),
.Y(n_4257)
);

OR2x2_ASAP7_75t_L g4258 ( 
.A(n_4128),
.B(n_178),
.Y(n_4258)
);

INVx1_ASAP7_75t_SL g4259 ( 
.A(n_4128),
.Y(n_4259)
);

OAI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_4130),
.A2(n_181),
.B1(n_178),
.B2(n_179),
.Y(n_4260)
);

NAND4xp25_ASAP7_75t_SL g4261 ( 
.A(n_4128),
.B(n_186),
.C(n_184),
.D(n_185),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4096),
.Y(n_4262)
);

AOI221xp5_ASAP7_75t_L g4263 ( 
.A1(n_4130),
.A2(n_205),
.B1(n_214),
.B2(n_194),
.C(n_184),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_4128),
.B(n_185),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_4128),
.B(n_186),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_4069),
.A2(n_188),
.B(n_189),
.Y(n_4266)
);

OAI22xp5_ASAP7_75t_L g4267 ( 
.A1(n_4130),
.A2(n_193),
.B1(n_190),
.B2(n_191),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4096),
.Y(n_4268)
);

INVx1_ASAP7_75t_SL g4269 ( 
.A(n_4128),
.Y(n_4269)
);

INVxp67_ASAP7_75t_L g4270 ( 
.A(n_4066),
.Y(n_4270)
);

OAI22xp33_ASAP7_75t_L g4271 ( 
.A1(n_4128),
.A2(n_194),
.B1(n_190),
.B2(n_191),
.Y(n_4271)
);

INVx2_ASAP7_75t_SL g4272 ( 
.A(n_4078),
.Y(n_4272)
);

AND2x2_ASAP7_75t_L g4273 ( 
.A(n_4128),
.B(n_195),
.Y(n_4273)
);

AOI21xp33_ASAP7_75t_SL g4274 ( 
.A1(n_4069),
.A2(n_196),
.B(n_200),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4096),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4128),
.B(n_196),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4096),
.Y(n_4277)
);

AOI221xp5_ASAP7_75t_L g4278 ( 
.A1(n_4130),
.A2(n_220),
.B1(n_230),
.B2(n_209),
.C(n_200),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4096),
.Y(n_4279)
);

INVxp67_ASAP7_75t_L g4280 ( 
.A(n_4066),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4078),
.Y(n_4281)
);

AOI22xp33_ASAP7_75t_L g4282 ( 
.A1(n_4123),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_4282)
);

NOR2xp33_ASAP7_75t_L g4283 ( 
.A(n_4128),
.B(n_201),
.Y(n_4283)
);

AOI21xp33_ASAP7_75t_L g4284 ( 
.A1(n_4128),
.A2(n_204),
.B(n_206),
.Y(n_4284)
);

OAI222xp33_ASAP7_75t_L g4285 ( 
.A1(n_4128),
.A2(n_208),
.B1(n_211),
.B2(n_206),
.C1(n_207),
.C2(n_210),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4096),
.Y(n_4286)
);

AOI32xp33_ASAP7_75t_L g4287 ( 
.A1(n_4087),
.A2(n_215),
.A3(n_211),
.B1(n_213),
.B2(n_216),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_4128),
.B(n_213),
.Y(n_4288)
);

AOI22xp5_ASAP7_75t_L g4289 ( 
.A1(n_4128),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4096),
.Y(n_4290)
);

XOR2x2_ASAP7_75t_L g4291 ( 
.A(n_4066),
.B(n_218),
.Y(n_4291)
);

INVx2_ASAP7_75t_SL g4292 ( 
.A(n_4078),
.Y(n_4292)
);

OAI221xp5_ASAP7_75t_L g4293 ( 
.A1(n_4069),
.A2(n_222),
.B1(n_218),
.B2(n_221),
.C(n_224),
.Y(n_4293)
);

INVx2_ASAP7_75t_SL g4294 ( 
.A(n_4078),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_4128),
.B(n_222),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4096),
.Y(n_4296)
);

OR2x2_ASAP7_75t_L g4297 ( 
.A(n_4259),
.B(n_4269),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4248),
.B(n_224),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4168),
.B(n_225),
.Y(n_4299)
);

OAI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_4236),
.A2(n_4253),
.B1(n_4280),
.B2(n_4270),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_SL g4301 ( 
.A(n_4251),
.B(n_225),
.Y(n_4301)
);

INVxp67_ASAP7_75t_L g4302 ( 
.A(n_4150),
.Y(n_4302)
);

HB1xp67_ASAP7_75t_L g4303 ( 
.A(n_4291),
.Y(n_4303)
);

A2O1A1O1Ixp25_ASAP7_75t_L g4304 ( 
.A1(n_4247),
.A2(n_245),
.B(n_253),
.C(n_236),
.D(n_226),
.Y(n_4304)
);

AOI31xp33_ASAP7_75t_L g4305 ( 
.A1(n_4171),
.A2(n_4212),
.A3(n_4194),
.B(n_4166),
.Y(n_4305)
);

AOI22xp5_ASAP7_75t_L g4306 ( 
.A1(n_4148),
.A2(n_231),
.B1(n_228),
.B2(n_229),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_4272),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4234),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4243),
.Y(n_4309)
);

AOI221xp5_ASAP7_75t_L g4310 ( 
.A1(n_4274),
.A2(n_981),
.B1(n_982),
.B2(n_980),
.C(n_978),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4233),
.B(n_229),
.Y(n_4311)
);

AND2x4_ASAP7_75t_L g4312 ( 
.A(n_4292),
.B(n_984),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4273),
.Y(n_4313)
);

NAND2xp33_ASAP7_75t_SL g4314 ( 
.A(n_4294),
.B(n_231),
.Y(n_4314)
);

AOI22xp5_ASAP7_75t_L g4315 ( 
.A1(n_4239),
.A2(n_987),
.B1(n_988),
.B2(n_986),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4295),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_4287),
.B(n_232),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_4180),
.B(n_232),
.Y(n_4318)
);

OAI21xp33_ASAP7_75t_SL g4319 ( 
.A1(n_4185),
.A2(n_233),
.B(n_234),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_4241),
.B(n_233),
.Y(n_4320)
);

AND2x4_ASAP7_75t_L g4321 ( 
.A(n_4187),
.B(n_988),
.Y(n_4321)
);

AND2x2_ASAP7_75t_L g4322 ( 
.A(n_4249),
.B(n_4262),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_4281),
.Y(n_4323)
);

AOI22xp33_ASAP7_75t_L g4324 ( 
.A1(n_4268),
.A2(n_4277),
.B1(n_4279),
.B2(n_4275),
.Y(n_4324)
);

INVx2_ASAP7_75t_L g4325 ( 
.A(n_4149),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_4286),
.B(n_234),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4290),
.B(n_235),
.Y(n_4327)
);

OAI22xp5_ASAP7_75t_L g4328 ( 
.A1(n_4293),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4237),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4296),
.B(n_237),
.Y(n_4330)
);

NOR2x1_ASAP7_75t_L g4331 ( 
.A(n_4285),
.B(n_239),
.Y(n_4331)
);

AOI221xp5_ASAP7_75t_L g4332 ( 
.A1(n_4250),
.A2(n_242),
.B1(n_239),
.B2(n_240),
.C(n_243),
.Y(n_4332)
);

AOI22xp5_ASAP7_75t_L g4333 ( 
.A1(n_4255),
.A2(n_243),
.B1(n_240),
.B2(n_242),
.Y(n_4333)
);

OAI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_4266),
.A2(n_246),
.B(n_245),
.Y(n_4334)
);

NAND2xp33_ASAP7_75t_L g4335 ( 
.A(n_4181),
.B(n_244),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_4167),
.B(n_4283),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4205),
.B(n_246),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4258),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4235),
.Y(n_4339)
);

NOR2xp33_ASAP7_75t_L g4340 ( 
.A(n_4189),
.B(n_247),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_4203),
.B(n_247),
.Y(n_4341)
);

NAND2xp33_ASAP7_75t_L g4342 ( 
.A(n_4183),
.B(n_248),
.Y(n_4342)
);

OAI31xp33_ASAP7_75t_L g4343 ( 
.A1(n_4151),
.A2(n_251),
.A3(n_249),
.B(n_250),
.Y(n_4343)
);

OR2x2_ASAP7_75t_L g4344 ( 
.A(n_4244),
.B(n_251),
.Y(n_4344)
);

OAI332xp33_ASAP7_75t_L g4345 ( 
.A1(n_4152),
.A2(n_4163),
.A3(n_4162),
.B1(n_4154),
.B2(n_4177),
.B3(n_4201),
.C1(n_4200),
.C2(n_4199),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4252),
.Y(n_4346)
);

OR2x6_ASAP7_75t_L g4347 ( 
.A(n_4179),
.B(n_252),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_4254),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_4240),
.A2(n_254),
.B(n_253),
.Y(n_4349)
);

NOR2xp33_ASAP7_75t_L g4350 ( 
.A(n_4264),
.B(n_252),
.Y(n_4350)
);

O2A1O1Ixp33_ASAP7_75t_L g4351 ( 
.A1(n_4160),
.A2(n_256),
.B(n_254),
.C(n_255),
.Y(n_4351)
);

OAI22xp5_ASAP7_75t_L g4352 ( 
.A1(n_4174),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_4352)
);

OAI21xp33_ASAP7_75t_L g4353 ( 
.A1(n_4173),
.A2(n_258),
.B(n_259),
.Y(n_4353)
);

AO21x1_ASAP7_75t_L g4354 ( 
.A1(n_4238),
.A2(n_259),
.B(n_260),
.Y(n_4354)
);

AOI22xp5_ASAP7_75t_L g4355 ( 
.A1(n_4261),
.A2(n_980),
.B1(n_984),
.B2(n_977),
.Y(n_4355)
);

OAI22xp5_ASAP7_75t_L g4356 ( 
.A1(n_4242),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_4356)
);

AOI21xp33_ASAP7_75t_SL g4357 ( 
.A1(n_4271),
.A2(n_987),
.B(n_985),
.Y(n_4357)
);

OAI22xp33_ASAP7_75t_L g4358 ( 
.A1(n_4289),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_4358)
);

AOI21xp33_ASAP7_75t_SL g4359 ( 
.A1(n_4256),
.A2(n_265),
.B(n_266),
.Y(n_4359)
);

NAND3xp33_ASAP7_75t_L g4360 ( 
.A(n_4186),
.B(n_265),
.C(n_267),
.Y(n_4360)
);

AOI32xp33_ASAP7_75t_L g4361 ( 
.A1(n_4225),
.A2(n_269),
.A3(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_4361)
);

NOR2xp33_ASAP7_75t_L g4362 ( 
.A(n_4265),
.B(n_268),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4276),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4288),
.Y(n_4364)
);

INVxp67_ASAP7_75t_L g4365 ( 
.A(n_4198),
.Y(n_4365)
);

INVxp67_ASAP7_75t_L g4366 ( 
.A(n_4209),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_4191),
.B(n_271),
.Y(n_4367)
);

OAI22xp5_ASAP7_75t_L g4368 ( 
.A1(n_4282),
.A2(n_274),
.B1(n_271),
.B2(n_272),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_4182),
.Y(n_4369)
);

AOI22xp33_ASAP7_75t_L g4370 ( 
.A1(n_4216),
.A2(n_275),
.B1(n_272),
.B2(n_274),
.Y(n_4370)
);

AOI22xp5_ASAP7_75t_L g4371 ( 
.A1(n_4227),
.A2(n_976),
.B1(n_985),
.B2(n_975),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4175),
.Y(n_4372)
);

XNOR2x1_ASAP7_75t_L g4373 ( 
.A(n_4257),
.B(n_277),
.Y(n_4373)
);

AOI22xp5_ASAP7_75t_L g4374 ( 
.A1(n_4211),
.A2(n_976),
.B1(n_989),
.B2(n_975),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4176),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_4158),
.B(n_277),
.Y(n_4376)
);

NOR2xp33_ASAP7_75t_L g4377 ( 
.A(n_4284),
.B(n_278),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_4206),
.B(n_279),
.Y(n_4378)
);

OAI21xp5_ASAP7_75t_SL g4379 ( 
.A1(n_4208),
.A2(n_280),
.B(n_281),
.Y(n_4379)
);

AOI322xp5_ASAP7_75t_L g4380 ( 
.A1(n_4219),
.A2(n_286),
.A3(n_285),
.B1(n_283),
.B2(n_281),
.C1(n_282),
.C2(n_284),
.Y(n_4380)
);

AOI321xp33_ASAP7_75t_L g4381 ( 
.A1(n_4196),
.A2(n_968),
.A3(n_966),
.B1(n_969),
.B2(n_967),
.C(n_965),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_4197),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_4210),
.Y(n_4383)
);

HB1xp67_ASAP7_75t_L g4384 ( 
.A(n_4188),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_4229),
.B(n_287),
.Y(n_4385)
);

AOI21xp5_ASAP7_75t_L g4386 ( 
.A1(n_4153),
.A2(n_288),
.B(n_289),
.Y(n_4386)
);

AOI21xp33_ASAP7_75t_SL g4387 ( 
.A1(n_4188),
.A2(n_973),
.B(n_971),
.Y(n_4387)
);

OR2x2_ASAP7_75t_L g4388 ( 
.A(n_4178),
.B(n_291),
.Y(n_4388)
);

OAI22xp5_ASAP7_75t_SL g4389 ( 
.A1(n_4220),
.A2(n_294),
.B1(n_291),
.B2(n_292),
.Y(n_4389)
);

AND2x2_ASAP7_75t_L g4390 ( 
.A(n_4207),
.B(n_292),
.Y(n_4390)
);

OAI32xp33_ASAP7_75t_L g4391 ( 
.A1(n_4214),
.A2(n_315),
.A3(n_324),
.B1(n_305),
.B2(n_294),
.Y(n_4391)
);

AOI211x1_ASAP7_75t_L g4392 ( 
.A1(n_4232),
.A2(n_4165),
.B(n_4170),
.C(n_4169),
.Y(n_4392)
);

OAI222xp33_ASAP7_75t_L g4393 ( 
.A1(n_4184),
.A2(n_297),
.B1(n_301),
.B2(n_295),
.C1(n_296),
.C2(n_299),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_4159),
.A2(n_296),
.B(n_299),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4193),
.Y(n_4395)
);

AND2x4_ASAP7_75t_L g4396 ( 
.A(n_4222),
.B(n_960),
.Y(n_4396)
);

AOI22xp5_ASAP7_75t_L g4397 ( 
.A1(n_4245),
.A2(n_964),
.B1(n_965),
.B2(n_963),
.Y(n_4397)
);

O2A1O1Ixp33_ASAP7_75t_L g4398 ( 
.A1(n_4218),
.A2(n_303),
.B(n_301),
.C(n_302),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_4204),
.B(n_302),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4164),
.Y(n_4400)
);

NOR3xp33_ASAP7_75t_L g4401 ( 
.A(n_4161),
.B(n_303),
.C(n_305),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4157),
.Y(n_4402)
);

O2A1O1Ixp33_ASAP7_75t_L g4403 ( 
.A1(n_4202),
.A2(n_309),
.B(n_306),
.C(n_308),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_4172),
.B(n_308),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4192),
.B(n_311),
.Y(n_4405)
);

A2O1A1Ixp33_ASAP7_75t_SL g4406 ( 
.A1(n_4230),
.A2(n_313),
.B(n_311),
.C(n_312),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4260),
.Y(n_4407)
);

AOI22xp5_ASAP7_75t_L g4408 ( 
.A1(n_4246),
.A2(n_316),
.B1(n_312),
.B2(n_314),
.Y(n_4408)
);

O2A1O1Ixp33_ASAP7_75t_L g4409 ( 
.A1(n_4267),
.A2(n_319),
.B(n_314),
.C(n_318),
.Y(n_4409)
);

AOI222xp33_ASAP7_75t_L g4410 ( 
.A1(n_4263),
.A2(n_321),
.B1(n_323),
.B2(n_318),
.C1(n_320),
.C2(n_322),
.Y(n_4410)
);

NOR2xp33_ASAP7_75t_L g4411 ( 
.A(n_4217),
.B(n_320),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_4278),
.B(n_321),
.Y(n_4412)
);

AND2x2_ASAP7_75t_L g4413 ( 
.A(n_4155),
.B(n_322),
.Y(n_4413)
);

AOI21xp5_ASAP7_75t_L g4414 ( 
.A1(n_4223),
.A2(n_323),
.B(n_325),
.Y(n_4414)
);

INVx1_ASAP7_75t_SL g4415 ( 
.A(n_4226),
.Y(n_4415)
);

INVx3_ASAP7_75t_SL g4416 ( 
.A(n_4297),
.Y(n_4416)
);

AOI21xp5_ASAP7_75t_L g4417 ( 
.A1(n_4305),
.A2(n_4147),
.B(n_4156),
.Y(n_4417)
);

OAI21xp5_ASAP7_75t_SL g4418 ( 
.A1(n_4324),
.A2(n_4228),
.B(n_4221),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4302),
.Y(n_4419)
);

NOR4xp25_ASAP7_75t_L g4420 ( 
.A(n_4300),
.B(n_4213),
.C(n_4195),
.D(n_4231),
.Y(n_4420)
);

AOI211xp5_ASAP7_75t_L g4421 ( 
.A1(n_4301),
.A2(n_4190),
.B(n_4224),
.C(n_4215),
.Y(n_4421)
);

OAI211xp5_ASAP7_75t_L g4422 ( 
.A1(n_4304),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_4422)
);

O2A1O1Ixp33_ASAP7_75t_L g4423 ( 
.A1(n_4406),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_4423)
);

AOI221xp5_ASAP7_75t_L g4424 ( 
.A1(n_4392),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.C(n_332),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4299),
.Y(n_4425)
);

NAND4xp25_ASAP7_75t_L g4426 ( 
.A(n_4336),
.B(n_332),
.C(n_330),
.D(n_331),
.Y(n_4426)
);

NOR2xp33_ASAP7_75t_L g4427 ( 
.A(n_4303),
.B(n_4319),
.Y(n_4427)
);

AOI211xp5_ASAP7_75t_L g4428 ( 
.A1(n_4354),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_4428)
);

AOI21xp33_ASAP7_75t_L g4429 ( 
.A1(n_4415),
.A2(n_335),
.B(n_336),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4322),
.Y(n_4430)
);

AOI22xp33_ASAP7_75t_L g4431 ( 
.A1(n_4331),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_4431)
);

AOI211xp5_ASAP7_75t_L g4432 ( 
.A1(n_4403),
.A2(n_4387),
.B(n_4353),
.C(n_4349),
.Y(n_4432)
);

AOI211x1_ASAP7_75t_L g4433 ( 
.A1(n_4317),
.A2(n_4334),
.B(n_4360),
.C(n_4394),
.Y(n_4433)
);

NOR3xp33_ASAP7_75t_L g4434 ( 
.A(n_4366),
.B(n_338),
.C(n_340),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_4312),
.B(n_341),
.Y(n_4435)
);

NAND3xp33_ASAP7_75t_L g4436 ( 
.A(n_4384),
.B(n_341),
.C(n_344),
.Y(n_4436)
);

NAND2xp67_ASAP7_75t_SL g4437 ( 
.A(n_4310),
.B(n_344),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4312),
.B(n_345),
.Y(n_4438)
);

AOI211xp5_ASAP7_75t_SL g4439 ( 
.A1(n_4345),
.A2(n_348),
.B(n_345),
.C(n_347),
.Y(n_4439)
);

AOI21xp33_ASAP7_75t_SL g4440 ( 
.A1(n_4398),
.A2(n_349),
.B(n_348),
.Y(n_4440)
);

AOI221x1_ASAP7_75t_SL g4441 ( 
.A1(n_4407),
.A2(n_350),
.B1(n_347),
.B2(n_349),
.C(n_353),
.Y(n_4441)
);

NAND4xp25_ASAP7_75t_L g4442 ( 
.A(n_4308),
.B(n_356),
.C(n_353),
.D(n_355),
.Y(n_4442)
);

AOI21xp33_ASAP7_75t_L g4443 ( 
.A1(n_4329),
.A2(n_356),
.B(n_358),
.Y(n_4443)
);

OAI22xp33_ASAP7_75t_L g4444 ( 
.A1(n_4405),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_4444)
);

AOI21xp5_ASAP7_75t_L g4445 ( 
.A1(n_4342),
.A2(n_361),
.B(n_362),
.Y(n_4445)
);

AOI21xp33_ASAP7_75t_L g4446 ( 
.A1(n_4382),
.A2(n_361),
.B(n_363),
.Y(n_4446)
);

OAI211xp5_ASAP7_75t_L g4447 ( 
.A1(n_4381),
.A2(n_365),
.B(n_363),
.C(n_364),
.Y(n_4447)
);

AO21x1_ASAP7_75t_L g4448 ( 
.A1(n_4314),
.A2(n_973),
.B(n_366),
.Y(n_4448)
);

NOR3xp33_ASAP7_75t_L g4449 ( 
.A(n_4365),
.B(n_366),
.C(n_368),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_4321),
.Y(n_4450)
);

O2A1O1Ixp33_ASAP7_75t_L g4451 ( 
.A1(n_4351),
.A2(n_370),
.B(n_368),
.C(n_369),
.Y(n_4451)
);

AOI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_4401),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_4452)
);

OAI21xp5_ASAP7_75t_L g4453 ( 
.A1(n_4414),
.A2(n_4335),
.B(n_4373),
.Y(n_4453)
);

NAND4xp25_ASAP7_75t_L g4454 ( 
.A(n_4309),
.B(n_374),
.C(n_371),
.D(n_372),
.Y(n_4454)
);

OAI21xp33_ASAP7_75t_L g4455 ( 
.A1(n_4313),
.A2(n_374),
.B(n_375),
.Y(n_4455)
);

NOR2xp33_ASAP7_75t_L g4456 ( 
.A(n_4316),
.B(n_375),
.Y(n_4456)
);

AOI221xp5_ASAP7_75t_L g4457 ( 
.A1(n_4357),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.C(n_380),
.Y(n_4457)
);

AOI221xp5_ASAP7_75t_L g4458 ( 
.A1(n_4307),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.C(n_381),
.Y(n_4458)
);

NOR3xp33_ASAP7_75t_L g4459 ( 
.A(n_4325),
.B(n_382),
.C(n_384),
.Y(n_4459)
);

AOI221xp5_ASAP7_75t_L g4460 ( 
.A1(n_4352),
.A2(n_386),
.B1(n_382),
.B2(n_385),
.C(n_389),
.Y(n_4460)
);

NAND4xp25_ASAP7_75t_L g4461 ( 
.A(n_4372),
.B(n_390),
.C(n_385),
.D(n_389),
.Y(n_4461)
);

AOI221xp5_ASAP7_75t_L g4462 ( 
.A1(n_4359),
.A2(n_394),
.B1(n_391),
.B2(n_393),
.C(n_395),
.Y(n_4462)
);

OAI211xp5_ASAP7_75t_L g4463 ( 
.A1(n_4410),
.A2(n_400),
.B(n_395),
.C(n_397),
.Y(n_4463)
);

OAI22xp33_ASAP7_75t_L g4464 ( 
.A1(n_4397),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_4355),
.B(n_403),
.Y(n_4465)
);

OAI21xp5_ASAP7_75t_SL g4466 ( 
.A1(n_4375),
.A2(n_404),
.B(n_405),
.Y(n_4466)
);

AOI22xp5_ASAP7_75t_L g4467 ( 
.A1(n_4411),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_4467)
);

NAND4xp25_ASAP7_75t_SL g4468 ( 
.A(n_4332),
.B(n_409),
.C(n_406),
.D(n_407),
.Y(n_4468)
);

NAND4xp75_ASAP7_75t_L g4469 ( 
.A(n_4323),
.B(n_412),
.C(n_410),
.D(n_411),
.Y(n_4469)
);

AOI221xp5_ASAP7_75t_L g4470 ( 
.A1(n_4393),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.C(n_416),
.Y(n_4470)
);

AOI21xp5_ASAP7_75t_L g4471 ( 
.A1(n_4298),
.A2(n_414),
.B(n_415),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_SL g4472 ( 
.A(n_4338),
.B(n_416),
.Y(n_4472)
);

AOI21xp5_ASAP7_75t_L g4473 ( 
.A1(n_4412),
.A2(n_418),
.B(n_421),
.Y(n_4473)
);

AOI221xp5_ASAP7_75t_L g4474 ( 
.A1(n_4358),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.C(n_424),
.Y(n_4474)
);

AOI221xp5_ASAP7_75t_L g4475 ( 
.A1(n_4391),
.A2(n_425),
.B1(n_422),
.B2(n_424),
.C(n_427),
.Y(n_4475)
);

A2O1A1Ixp33_ASAP7_75t_L g4476 ( 
.A1(n_4409),
.A2(n_435),
.B(n_444),
.C(n_425),
.Y(n_4476)
);

NAND3xp33_ASAP7_75t_L g4477 ( 
.A(n_4369),
.B(n_427),
.C(n_428),
.Y(n_4477)
);

OAI22xp5_ASAP7_75t_L g4478 ( 
.A1(n_4408),
.A2(n_431),
.B1(n_428),
.B2(n_429),
.Y(n_4478)
);

AND3x1_ASAP7_75t_L g4479 ( 
.A(n_4343),
.B(n_431),
.C(n_432),
.Y(n_4479)
);

AOI22xp5_ASAP7_75t_L g4480 ( 
.A1(n_4383),
.A2(n_437),
.B1(n_433),
.B2(n_434),
.Y(n_4480)
);

NOR4xp25_ASAP7_75t_L g4481 ( 
.A(n_4339),
.B(n_440),
.C(n_438),
.D(n_439),
.Y(n_4481)
);

NOR3xp33_ASAP7_75t_L g4482 ( 
.A(n_4346),
.B(n_4363),
.C(n_4348),
.Y(n_4482)
);

AOI221xp5_ASAP7_75t_L g4483 ( 
.A1(n_4328),
.A2(n_440),
.B1(n_438),
.B2(n_439),
.C(n_441),
.Y(n_4483)
);

AOI222xp33_ASAP7_75t_L g4484 ( 
.A1(n_4389),
.A2(n_444),
.B1(n_446),
.B2(n_442),
.C1(n_443),
.C2(n_445),
.Y(n_4484)
);

AOI222xp33_ASAP7_75t_L g4485 ( 
.A1(n_4364),
.A2(n_448),
.B1(n_450),
.B2(n_443),
.C1(n_447),
.C2(n_449),
.Y(n_4485)
);

OAI211xp5_ASAP7_75t_L g4486 ( 
.A1(n_4380),
.A2(n_451),
.B(n_447),
.C(n_450),
.Y(n_4486)
);

NOR2x1_ASAP7_75t_L g4487 ( 
.A(n_4379),
.B(n_451),
.Y(n_4487)
);

NAND3xp33_ASAP7_75t_L g4488 ( 
.A(n_4326),
.B(n_453),
.C(n_455),
.Y(n_4488)
);

OAI21xp33_ASAP7_75t_L g4489 ( 
.A1(n_4395),
.A2(n_455),
.B(n_456),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_4396),
.B(n_458),
.Y(n_4490)
);

NAND3xp33_ASAP7_75t_SL g4491 ( 
.A(n_4361),
.B(n_461),
.C(n_460),
.Y(n_4491)
);

NOR3xp33_ASAP7_75t_L g4492 ( 
.A(n_4402),
.B(n_459),
.C(n_461),
.Y(n_4492)
);

OAI22xp33_ASAP7_75t_L g4493 ( 
.A1(n_4404),
.A2(n_465),
.B1(n_462),
.B2(n_463),
.Y(n_4493)
);

AOI22xp5_ASAP7_75t_L g4494 ( 
.A1(n_4311),
.A2(n_469),
.B1(n_465),
.B2(n_467),
.Y(n_4494)
);

NOR2xp33_ASAP7_75t_L g4495 ( 
.A(n_4385),
.B(n_469),
.Y(n_4495)
);

NOR3xp33_ASAP7_75t_L g4496 ( 
.A(n_4400),
.B(n_470),
.C(n_471),
.Y(n_4496)
);

O2A1O1Ixp33_ASAP7_75t_L g4497 ( 
.A1(n_4356),
.A2(n_473),
.B(n_470),
.C(n_472),
.Y(n_4497)
);

OAI21xp5_ASAP7_75t_SL g4498 ( 
.A1(n_4330),
.A2(n_472),
.B(n_473),
.Y(n_4498)
);

AOI21xp5_ASAP7_75t_L g4499 ( 
.A1(n_4318),
.A2(n_4347),
.B(n_4327),
.Y(n_4499)
);

OAI221xp5_ASAP7_75t_L g4500 ( 
.A1(n_4347),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.C(n_478),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4321),
.Y(n_4501)
);

A2O1A1Ixp33_ASAP7_75t_L g4502 ( 
.A1(n_4377),
.A2(n_478),
.B(n_474),
.C(n_475),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4337),
.Y(n_4503)
);

A2O1A1Ixp33_ASAP7_75t_L g4504 ( 
.A1(n_4340),
.A2(n_4386),
.B(n_4362),
.C(n_4350),
.Y(n_4504)
);

AOI221xp5_ASAP7_75t_L g4505 ( 
.A1(n_4368),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.C(n_483),
.Y(n_4505)
);

OAI221xp5_ASAP7_75t_L g4506 ( 
.A1(n_4320),
.A2(n_4370),
.B1(n_4341),
.B2(n_4333),
.C(n_4315),
.Y(n_4506)
);

OAI221xp5_ASAP7_75t_L g4507 ( 
.A1(n_4306),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.C(n_485),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4396),
.B(n_485),
.Y(n_4508)
);

AOI21xp5_ASAP7_75t_L g4509 ( 
.A1(n_4399),
.A2(n_487),
.B(n_488),
.Y(n_4509)
);

AOI221xp5_ASAP7_75t_SL g4510 ( 
.A1(n_4378),
.A2(n_491),
.B1(n_487),
.B2(n_489),
.C(n_492),
.Y(n_4510)
);

NAND4xp25_ASAP7_75t_L g4511 ( 
.A(n_4371),
.B(n_492),
.C(n_489),
.D(n_491),
.Y(n_4511)
);

NAND3xp33_ASAP7_75t_L g4512 ( 
.A(n_4374),
.B(n_494),
.C(n_495),
.Y(n_4512)
);

NOR2xp33_ASAP7_75t_L g4513 ( 
.A(n_4367),
.B(n_494),
.Y(n_4513)
);

AOI22xp5_ASAP7_75t_L g4514 ( 
.A1(n_4390),
.A2(n_497),
.B1(n_495),
.B2(n_496),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_4413),
.B(n_496),
.Y(n_4515)
);

OAI32xp33_ASAP7_75t_L g4516 ( 
.A1(n_4344),
.A2(n_502),
.A3(n_497),
.B1(n_498),
.B2(n_503),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4376),
.B(n_498),
.Y(n_4517)
);

NOR4xp25_ASAP7_75t_L g4518 ( 
.A(n_4388),
.B(n_505),
.C(n_503),
.D(n_504),
.Y(n_4518)
);

NOR2xp67_ASAP7_75t_SL g4519 ( 
.A(n_4297),
.B(n_504),
.Y(n_4519)
);

AOI222xp33_ASAP7_75t_L g4520 ( 
.A1(n_4302),
.A2(n_510),
.B1(n_512),
.B2(n_508),
.C1(n_509),
.C2(n_511),
.Y(n_4520)
);

NOR2xp67_ASAP7_75t_L g4521 ( 
.A(n_4302),
.B(n_508),
.Y(n_4521)
);

OAI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_4302),
.A2(n_510),
.B(n_512),
.Y(n_4522)
);

AOI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_4305),
.A2(n_513),
.B(n_514),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4297),
.Y(n_4524)
);

NAND4xp75_ASAP7_75t_L g4525 ( 
.A(n_4322),
.B(n_519),
.C(n_516),
.D(n_518),
.Y(n_4525)
);

AOI21xp5_ASAP7_75t_SL g4526 ( 
.A1(n_4398),
.A2(n_516),
.B(n_520),
.Y(n_4526)
);

AOI22xp33_ASAP7_75t_L g4527 ( 
.A1(n_4303),
.A2(n_525),
.B1(n_523),
.B2(n_524),
.Y(n_4527)
);

OA21x2_ASAP7_75t_L g4528 ( 
.A1(n_4384),
.A2(n_524),
.B(n_525),
.Y(n_4528)
);

AOI211xp5_ASAP7_75t_L g4529 ( 
.A1(n_4300),
.A2(n_528),
.B(n_526),
.C(n_527),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4302),
.B(n_528),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4297),
.Y(n_4531)
);

NAND4xp25_ASAP7_75t_L g4532 ( 
.A(n_4324),
.B(n_532),
.C(n_530),
.D(n_531),
.Y(n_4532)
);

OAI21xp33_ASAP7_75t_SL g4533 ( 
.A1(n_4305),
.A2(n_530),
.B(n_532),
.Y(n_4533)
);

NOR2xp67_ASAP7_75t_L g4534 ( 
.A(n_4302),
.B(n_533),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4297),
.Y(n_4535)
);

AOI222xp33_ASAP7_75t_L g4536 ( 
.A1(n_4302),
.A2(n_536),
.B1(n_538),
.B2(n_533),
.C1(n_534),
.C2(n_537),
.Y(n_4536)
);

O2A1O1Ixp33_ASAP7_75t_SL g4537 ( 
.A1(n_4301),
.A2(n_537),
.B(n_534),
.C(n_536),
.Y(n_4537)
);

NOR2x1_ASAP7_75t_L g4538 ( 
.A(n_4297),
.B(n_539),
.Y(n_4538)
);

AOI21xp5_ASAP7_75t_L g4539 ( 
.A1(n_4305),
.A2(n_540),
.B(n_543),
.Y(n_4539)
);

A2O1A1Ixp33_ASAP7_75t_L g4540 ( 
.A1(n_4398),
.A2(n_544),
.B(n_540),
.C(n_543),
.Y(n_4540)
);

AOI221xp5_ASAP7_75t_L g4541 ( 
.A1(n_4305),
.A2(n_549),
.B1(n_545),
.B2(n_546),
.C(n_550),
.Y(n_4541)
);

OAI22xp5_ASAP7_75t_L g4542 ( 
.A1(n_4324),
.A2(n_553),
.B1(n_551),
.B2(n_552),
.Y(n_4542)
);

NOR3xp33_ASAP7_75t_L g4543 ( 
.A(n_4305),
.B(n_551),
.C(n_552),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4297),
.Y(n_4544)
);

OAI21xp5_ASAP7_75t_SL g4545 ( 
.A1(n_4305),
.A2(n_553),
.B(n_555),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4297),
.Y(n_4546)
);

AOI221xp5_ASAP7_75t_L g4547 ( 
.A1(n_4305),
.A2(n_559),
.B1(n_555),
.B2(n_556),
.C(n_560),
.Y(n_4547)
);

A2O1A1Ixp33_ASAP7_75t_L g4548 ( 
.A1(n_4398),
.A2(n_562),
.B(n_559),
.C(n_561),
.Y(n_4548)
);

AOI21xp33_ASAP7_75t_L g4549 ( 
.A1(n_4305),
.A2(n_563),
.B(n_564),
.Y(n_4549)
);

AOI211xp5_ASAP7_75t_SL g4550 ( 
.A1(n_4305),
.A2(n_565),
.B(n_563),
.C(n_564),
.Y(n_4550)
);

OAI211xp5_ASAP7_75t_L g4551 ( 
.A1(n_4304),
.A2(n_570),
.B(n_566),
.C(n_569),
.Y(n_4551)
);

AOI22xp5_ASAP7_75t_L g4552 ( 
.A1(n_4322),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_4552)
);

NOR2xp33_ASAP7_75t_L g4553 ( 
.A(n_4302),
.B(n_571),
.Y(n_4553)
);

OAI21xp33_ASAP7_75t_SL g4554 ( 
.A1(n_4305),
.A2(n_573),
.B(n_574),
.Y(n_4554)
);

OAI211xp5_ASAP7_75t_SL g4555 ( 
.A1(n_4324),
.A2(n_576),
.B(n_574),
.C(n_575),
.Y(n_4555)
);

OAI21xp33_ASAP7_75t_L g4556 ( 
.A1(n_4324),
.A2(n_575),
.B(n_577),
.Y(n_4556)
);

AOI21xp5_ASAP7_75t_L g4557 ( 
.A1(n_4305),
.A2(n_577),
.B(n_578),
.Y(n_4557)
);

AOI21xp5_ASAP7_75t_L g4558 ( 
.A1(n_4305),
.A2(n_579),
.B(n_581),
.Y(n_4558)
);

AOI22xp5_ASAP7_75t_L g4559 ( 
.A1(n_4322),
.A2(n_584),
.B1(n_581),
.B2(n_582),
.Y(n_4559)
);

OAI21xp33_ASAP7_75t_L g4560 ( 
.A1(n_4324),
.A2(n_585),
.B(n_587),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4302),
.B(n_585),
.Y(n_4561)
);

NAND4xp25_ASAP7_75t_L g4562 ( 
.A(n_4324),
.B(n_590),
.C(n_588),
.D(n_589),
.Y(n_4562)
);

OAI221xp5_ASAP7_75t_L g4563 ( 
.A1(n_4324),
.A2(n_590),
.B1(n_588),
.B2(n_589),
.C(n_592),
.Y(n_4563)
);

AND2x4_ASAP7_75t_L g4564 ( 
.A(n_4312),
.B(n_592),
.Y(n_4564)
);

AOI211xp5_ASAP7_75t_SL g4565 ( 
.A1(n_4549),
.A2(n_595),
.B(n_593),
.C(n_594),
.Y(n_4565)
);

AOI21xp33_ASAP7_75t_L g4566 ( 
.A1(n_4427),
.A2(n_4554),
.B(n_4533),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4538),
.Y(n_4567)
);

OAI21x1_ASAP7_75t_SL g4568 ( 
.A1(n_4448),
.A2(n_593),
.B(n_594),
.Y(n_4568)
);

AOI21xp5_ASAP7_75t_L g4569 ( 
.A1(n_4423),
.A2(n_595),
.B(n_596),
.Y(n_4569)
);

AOI21xp33_ASAP7_75t_SL g4570 ( 
.A1(n_4416),
.A2(n_597),
.B(n_598),
.Y(n_4570)
);

NOR2xp33_ASAP7_75t_L g4571 ( 
.A(n_4501),
.B(n_597),
.Y(n_4571)
);

AOI22xp5_ASAP7_75t_L g4572 ( 
.A1(n_4422),
.A2(n_601),
.B1(n_599),
.B2(n_600),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_L g4573 ( 
.A(n_4450),
.B(n_599),
.Y(n_4573)
);

OAI322xp33_ASAP7_75t_L g4574 ( 
.A1(n_4523),
.A2(n_610),
.A3(n_609),
.B1(n_607),
.B2(n_601),
.C1(n_605),
.C2(n_608),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4521),
.Y(n_4575)
);

AOI221xp5_ASAP7_75t_L g4576 ( 
.A1(n_4543),
.A2(n_609),
.B1(n_605),
.B2(n_607),
.C(n_610),
.Y(n_4576)
);

NOR2xp33_ASAP7_75t_L g4577 ( 
.A(n_4545),
.B(n_4447),
.Y(n_4577)
);

AOI31xp33_ASAP7_75t_L g4578 ( 
.A1(n_4550),
.A2(n_614),
.A3(n_611),
.B(n_612),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4534),
.Y(n_4579)
);

AOI221xp5_ASAP7_75t_L g4580 ( 
.A1(n_4420),
.A2(n_615),
.B1(n_612),
.B2(n_614),
.C(n_616),
.Y(n_4580)
);

OAI221xp5_ASAP7_75t_L g4581 ( 
.A1(n_4439),
.A2(n_619),
.B1(n_616),
.B2(n_618),
.C(n_620),
.Y(n_4581)
);

AOI311xp33_ASAP7_75t_L g4582 ( 
.A1(n_4419),
.A2(n_620),
.A3(n_618),
.B(n_619),
.C(n_621),
.Y(n_4582)
);

AOI221xp5_ASAP7_75t_L g4583 ( 
.A1(n_4424),
.A2(n_624),
.B1(n_621),
.B2(n_623),
.C(n_625),
.Y(n_4583)
);

AOI322xp5_ASAP7_75t_L g4584 ( 
.A1(n_4491),
.A2(n_630),
.A3(n_628),
.B1(n_625),
.B2(n_623),
.C1(n_624),
.C2(n_626),
.Y(n_4584)
);

OAI211xp5_ASAP7_75t_L g4585 ( 
.A1(n_4551),
.A2(n_633),
.B(n_628),
.C(n_632),
.Y(n_4585)
);

OAI21xp33_ASAP7_75t_SL g4586 ( 
.A1(n_4524),
.A2(n_634),
.B(n_635),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4564),
.Y(n_4587)
);

OAI21xp5_ASAP7_75t_L g4588 ( 
.A1(n_4539),
.A2(n_636),
.B(n_637),
.Y(n_4588)
);

INVxp67_ASAP7_75t_L g4589 ( 
.A(n_4519),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4528),
.Y(n_4590)
);

XOR2xp5_ASAP7_75t_L g4591 ( 
.A(n_4535),
.B(n_636),
.Y(n_4591)
);

OR2x2_ASAP7_75t_L g4592 ( 
.A(n_4518),
.B(n_637),
.Y(n_4592)
);

OAI32xp33_ASAP7_75t_L g4593 ( 
.A1(n_4430),
.A2(n_4546),
.A3(n_4544),
.B1(n_4531),
.B2(n_4482),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4528),
.Y(n_4594)
);

OR2x2_ASAP7_75t_L g4595 ( 
.A(n_4481),
.B(n_638),
.Y(n_4595)
);

A2O1A1Ixp33_ASAP7_75t_L g4596 ( 
.A1(n_4441),
.A2(n_642),
.B(n_638),
.C(n_640),
.Y(n_4596)
);

INVx3_ASAP7_75t_L g4597 ( 
.A(n_4564),
.Y(n_4597)
);

AOI21xp33_ASAP7_75t_SL g4598 ( 
.A1(n_4542),
.A2(n_640),
.B(n_642),
.Y(n_4598)
);

OAI21xp5_ASAP7_75t_L g4599 ( 
.A1(n_4557),
.A2(n_643),
.B(n_644),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4469),
.Y(n_4600)
);

OA21x2_ASAP7_75t_SL g4601 ( 
.A1(n_4472),
.A2(n_643),
.B(n_645),
.Y(n_4601)
);

AOI21xp33_ASAP7_75t_L g4602 ( 
.A1(n_4432),
.A2(n_647),
.B(n_648),
.Y(n_4602)
);

OAI22xp33_ASAP7_75t_L g4603 ( 
.A1(n_4452),
.A2(n_650),
.B1(n_647),
.B2(n_648),
.Y(n_4603)
);

AOI22xp5_ASAP7_75t_L g4604 ( 
.A1(n_4479),
.A2(n_654),
.B1(n_651),
.B2(n_653),
.Y(n_4604)
);

NAND4xp25_ASAP7_75t_L g4605 ( 
.A(n_4433),
.B(n_655),
.C(n_651),
.D(n_653),
.Y(n_4605)
);

HB1xp67_ASAP7_75t_L g4606 ( 
.A(n_4525),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4431),
.B(n_655),
.Y(n_4607)
);

AOI21xp5_ASAP7_75t_L g4608 ( 
.A1(n_4558),
.A2(n_656),
.B(n_657),
.Y(n_4608)
);

A2O1A1Ixp33_ASAP7_75t_SL g4609 ( 
.A1(n_4425),
.A2(n_659),
.B(n_656),
.C(n_658),
.Y(n_4609)
);

OAI21xp33_ASAP7_75t_L g4610 ( 
.A1(n_4418),
.A2(n_659),
.B(n_660),
.Y(n_4610)
);

OAI22xp5_ASAP7_75t_L g4611 ( 
.A1(n_4421),
.A2(n_666),
.B1(n_662),
.B2(n_665),
.Y(n_4611)
);

AOI22x1_ASAP7_75t_L g4612 ( 
.A1(n_4417),
.A2(n_668),
.B1(n_662),
.B2(n_667),
.Y(n_4612)
);

NOR4xp25_ASAP7_75t_L g4613 ( 
.A(n_4504),
.B(n_670),
.C(n_668),
.D(n_669),
.Y(n_4613)
);

NAND5xp2_ASAP7_75t_L g4614 ( 
.A(n_4503),
.B(n_671),
.C(n_669),
.D(n_670),
.E(n_672),
.Y(n_4614)
);

AOI322xp5_ASAP7_75t_L g4615 ( 
.A1(n_4541),
.A2(n_4547),
.A3(n_4444),
.B1(n_4487),
.B2(n_4556),
.C1(n_4560),
.C2(n_4493),
.Y(n_4615)
);

AOI221xp5_ASAP7_75t_L g4616 ( 
.A1(n_4440),
.A2(n_673),
.B1(n_671),
.B2(n_672),
.C(n_674),
.Y(n_4616)
);

AOI211xp5_ASAP7_75t_L g4617 ( 
.A1(n_4526),
.A2(n_675),
.B(n_673),
.C(n_674),
.Y(n_4617)
);

AOI221xp5_ASAP7_75t_L g4618 ( 
.A1(n_4537),
.A2(n_678),
.B1(n_676),
.B2(n_677),
.C(n_679),
.Y(n_4618)
);

O2A1O1Ixp33_ASAP7_75t_L g4619 ( 
.A1(n_4540),
.A2(n_679),
.B(n_676),
.C(n_678),
.Y(n_4619)
);

AOI22xp33_ASAP7_75t_SL g4620 ( 
.A1(n_4463),
.A2(n_682),
.B1(n_680),
.B2(n_681),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4435),
.Y(n_4621)
);

INVxp67_ASAP7_75t_L g4622 ( 
.A(n_4553),
.Y(n_4622)
);

AOI22xp5_ASAP7_75t_L g4623 ( 
.A1(n_4468),
.A2(n_4486),
.B1(n_4555),
.B2(n_4532),
.Y(n_4623)
);

NAND3xp33_ASAP7_75t_L g4624 ( 
.A(n_4428),
.B(n_681),
.C(n_682),
.Y(n_4624)
);

AOI322xp5_ASAP7_75t_L g4625 ( 
.A1(n_4510),
.A2(n_683),
.A3(n_684),
.B1(n_685),
.B2(n_686),
.C1(n_687),
.C2(n_689),
.Y(n_4625)
);

NAND4xp25_ASAP7_75t_SL g4626 ( 
.A(n_4499),
.B(n_687),
.C(n_683),
.D(n_684),
.Y(n_4626)
);

OAI22xp5_ASAP7_75t_L g4627 ( 
.A1(n_4563),
.A2(n_698),
.B1(n_691),
.B2(n_696),
.Y(n_4627)
);

NOR2x1_ASAP7_75t_L g4628 ( 
.A(n_4436),
.B(n_696),
.Y(n_4628)
);

XNOR2xp5_ASAP7_75t_L g4629 ( 
.A(n_4426),
.B(n_698),
.Y(n_4629)
);

AOI221xp5_ASAP7_75t_L g4630 ( 
.A1(n_4453),
.A2(n_703),
.B1(n_700),
.B2(n_702),
.C(n_705),
.Y(n_4630)
);

NAND2x1_ASAP7_75t_L g4631 ( 
.A(n_4438),
.B(n_4490),
.Y(n_4631)
);

AOI22xp5_ASAP7_75t_L g4632 ( 
.A1(n_4562),
.A2(n_706),
.B1(n_700),
.B2(n_703),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4484),
.B(n_4520),
.Y(n_4633)
);

NAND2x1p5_ASAP7_75t_L g4634 ( 
.A(n_4445),
.B(n_706),
.Y(n_4634)
);

OAI22xp5_ASAP7_75t_L g4635 ( 
.A1(n_4527),
.A2(n_710),
.B1(n_707),
.B2(n_708),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_4536),
.B(n_711),
.Y(n_4636)
);

OAI21xp33_ASAP7_75t_L g4637 ( 
.A1(n_4506),
.A2(n_712),
.B(n_714),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4522),
.B(n_712),
.Y(n_4638)
);

XOR2x2_ASAP7_75t_L g4639 ( 
.A(n_4470),
.B(n_714),
.Y(n_4639)
);

AOI221xp5_ASAP7_75t_SL g4640 ( 
.A1(n_4473),
.A2(n_717),
.B1(n_715),
.B2(n_716),
.C(n_718),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4508),
.Y(n_4641)
);

AOI221xp5_ASAP7_75t_L g4642 ( 
.A1(n_4451),
.A2(n_720),
.B1(n_717),
.B2(n_719),
.C(n_722),
.Y(n_4642)
);

NOR2x1_ASAP7_75t_SL g4643 ( 
.A(n_4498),
.B(n_719),
.Y(n_4643)
);

HB1xp67_ASAP7_75t_L g4644 ( 
.A(n_4530),
.Y(n_4644)
);

OAI21xp5_ASAP7_75t_L g4645 ( 
.A1(n_4548),
.A2(n_720),
.B(n_722),
.Y(n_4645)
);

OAI21xp33_ASAP7_75t_L g4646 ( 
.A1(n_4511),
.A2(n_723),
.B(n_724),
.Y(n_4646)
);

AOI21xp33_ASAP7_75t_L g4647 ( 
.A1(n_4497),
.A2(n_724),
.B(n_725),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_SL g4648 ( 
.A(n_4475),
.B(n_726),
.Y(n_4648)
);

OAI21xp33_ASAP7_75t_L g4649 ( 
.A1(n_4561),
.A2(n_726),
.B(n_727),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4434),
.B(n_4495),
.Y(n_4650)
);

AOI21xp33_ASAP7_75t_SL g4651 ( 
.A1(n_4459),
.A2(n_727),
.B(n_728),
.Y(n_4651)
);

OAI221xp5_ASAP7_75t_L g4652 ( 
.A1(n_4529),
.A2(n_730),
.B1(n_728),
.B2(n_729),
.C(n_731),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4590),
.Y(n_4653)
);

NOR2xp33_ASAP7_75t_R g4654 ( 
.A(n_4626),
.B(n_4465),
.Y(n_4654)
);

NOR2x1_ASAP7_75t_L g4655 ( 
.A(n_4594),
.B(n_4477),
.Y(n_4655)
);

INVxp67_ASAP7_75t_L g4656 ( 
.A(n_4614),
.Y(n_4656)
);

AOI211xp5_ASAP7_75t_L g4657 ( 
.A1(n_4566),
.A2(n_4464),
.B(n_4429),
.C(n_4478),
.Y(n_4657)
);

OAI21x1_ASAP7_75t_SL g4658 ( 
.A1(n_4568),
.A2(n_4471),
.B(n_4509),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4597),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_4587),
.B(n_4513),
.Y(n_4660)
);

OAI221xp5_ASAP7_75t_L g4661 ( 
.A1(n_4572),
.A2(n_4466),
.B1(n_4476),
.B2(n_4457),
.C(n_4483),
.Y(n_4661)
);

NOR2xp33_ASAP7_75t_L g4662 ( 
.A(n_4597),
.B(n_4581),
.Y(n_4662)
);

INVx2_ASAP7_75t_SL g4663 ( 
.A(n_4575),
.Y(n_4663)
);

NAND3xp33_ASAP7_75t_L g4664 ( 
.A(n_4617),
.B(n_4462),
.C(n_4512),
.Y(n_4664)
);

AOI22xp5_ASAP7_75t_L g4665 ( 
.A1(n_4577),
.A2(n_4589),
.B1(n_4610),
.B2(n_4585),
.Y(n_4665)
);

OAI22xp33_ASAP7_75t_L g4666 ( 
.A1(n_4578),
.A2(n_4507),
.B1(n_4488),
.B2(n_4442),
.Y(n_4666)
);

OAI21xp33_ASAP7_75t_L g4667 ( 
.A1(n_4623),
.A2(n_4455),
.B(n_4489),
.Y(n_4667)
);

INVx3_ASAP7_75t_L g4668 ( 
.A(n_4579),
.Y(n_4668)
);

OAI22xp5_ASAP7_75t_L g4669 ( 
.A1(n_4604),
.A2(n_4502),
.B1(n_4467),
.B2(n_4515),
.Y(n_4669)
);

OAI22xp5_ASAP7_75t_L g4670 ( 
.A1(n_4632),
.A2(n_4517),
.B1(n_4514),
.B2(n_4552),
.Y(n_4670)
);

INVx2_ASAP7_75t_SL g4671 ( 
.A(n_4567),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4634),
.Y(n_4672)
);

OAI22xp5_ASAP7_75t_L g4673 ( 
.A1(n_4620),
.A2(n_4559),
.B1(n_4456),
.B2(n_4494),
.Y(n_4673)
);

OAI221xp5_ASAP7_75t_L g4674 ( 
.A1(n_4580),
.A2(n_4474),
.B1(n_4460),
.B2(n_4505),
.C(n_4458),
.Y(n_4674)
);

BUFx2_ASAP7_75t_L g4675 ( 
.A(n_4586),
.Y(n_4675)
);

OAI221xp5_ASAP7_75t_L g4676 ( 
.A1(n_4637),
.A2(n_4449),
.B1(n_4496),
.B2(n_4492),
.C(n_4446),
.Y(n_4676)
);

AOI322xp5_ASAP7_75t_L g4677 ( 
.A1(n_4633),
.A2(n_4443),
.A3(n_4480),
.B1(n_4437),
.B2(n_4454),
.C1(n_4461),
.C2(n_4485),
.Y(n_4677)
);

AOI221xp5_ASAP7_75t_L g4678 ( 
.A1(n_4593),
.A2(n_4516),
.B1(n_4500),
.B2(n_736),
.C(n_732),
.Y(n_4678)
);

OAI221xp5_ASAP7_75t_L g4679 ( 
.A1(n_4588),
.A2(n_736),
.B1(n_732),
.B2(n_735),
.C(n_737),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4643),
.Y(n_4680)
);

A2O1A1Ixp33_ASAP7_75t_L g4681 ( 
.A1(n_4609),
.A2(n_738),
.B(n_735),
.C(n_737),
.Y(n_4681)
);

OR2x2_ASAP7_75t_L g4682 ( 
.A(n_4613),
.B(n_738),
.Y(n_4682)
);

O2A1O1Ixp33_ASAP7_75t_SL g4683 ( 
.A1(n_4596),
.A2(n_741),
.B(n_739),
.C(n_740),
.Y(n_4683)
);

INVxp67_ASAP7_75t_L g4684 ( 
.A(n_4571),
.Y(n_4684)
);

NAND3xp33_ASAP7_75t_L g4685 ( 
.A(n_4565),
.B(n_741),
.C(n_742),
.Y(n_4685)
);

INVx2_ASAP7_75t_SL g4686 ( 
.A(n_4628),
.Y(n_4686)
);

AOI22xp5_ASAP7_75t_L g4687 ( 
.A1(n_4600),
.A2(n_745),
.B1(n_743),
.B2(n_744),
.Y(n_4687)
);

OAI22xp33_ASAP7_75t_SL g4688 ( 
.A1(n_4595),
.A2(n_746),
.B1(n_743),
.B2(n_744),
.Y(n_4688)
);

INVx1_ASAP7_75t_SL g4689 ( 
.A(n_4592),
.Y(n_4689)
);

OAI22xp33_ASAP7_75t_L g4690 ( 
.A1(n_4605),
.A2(n_748),
.B1(n_746),
.B2(n_747),
.Y(n_4690)
);

AOI21xp33_ASAP7_75t_L g4691 ( 
.A1(n_4631),
.A2(n_748),
.B(n_749),
.Y(n_4691)
);

NAND4xp25_ASAP7_75t_SL g4692 ( 
.A(n_4615),
.B(n_752),
.C(n_750),
.D(n_751),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4591),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4606),
.Y(n_4694)
);

OA22x2_ASAP7_75t_L g4695 ( 
.A1(n_4599),
.A2(n_754),
.B1(n_752),
.B2(n_753),
.Y(n_4695)
);

AOI221xp5_ASAP7_75t_L g4696 ( 
.A1(n_4602),
.A2(n_757),
.B1(n_754),
.B2(n_756),
.C(n_759),
.Y(n_4696)
);

AOI21xp5_ASAP7_75t_L g4697 ( 
.A1(n_4569),
.A2(n_756),
.B(n_759),
.Y(n_4697)
);

OAI21xp5_ASAP7_75t_L g4698 ( 
.A1(n_4624),
.A2(n_761),
.B(n_762),
.Y(n_4698)
);

AOI21xp5_ASAP7_75t_L g4699 ( 
.A1(n_4608),
.A2(n_762),
.B(n_763),
.Y(n_4699)
);

NAND4xp25_ASAP7_75t_L g4700 ( 
.A(n_4601),
.B(n_765),
.C(n_763),
.D(n_764),
.Y(n_4700)
);

AOI22xp33_ASAP7_75t_SL g4701 ( 
.A1(n_4612),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.Y(n_4701)
);

AOI21xp33_ASAP7_75t_L g4702 ( 
.A1(n_4622),
.A2(n_768),
.B(n_769),
.Y(n_4702)
);

AOI21xp5_ASAP7_75t_L g4703 ( 
.A1(n_4648),
.A2(n_770),
.B(n_771),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4573),
.Y(n_4704)
);

OAI21xp33_ASAP7_75t_L g4705 ( 
.A1(n_4650),
.A2(n_4646),
.B(n_4636),
.Y(n_4705)
);

CKINVDCx5p33_ASAP7_75t_R g4706 ( 
.A(n_4629),
.Y(n_4706)
);

AOI32xp33_ASAP7_75t_L g4707 ( 
.A1(n_4582),
.A2(n_774),
.A3(n_770),
.B1(n_773),
.B2(n_775),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4638),
.Y(n_4708)
);

AOI22xp5_ASAP7_75t_L g4709 ( 
.A1(n_4611),
.A2(n_777),
.B1(n_775),
.B2(n_776),
.Y(n_4709)
);

CKINVDCx5p33_ASAP7_75t_R g4710 ( 
.A(n_4639),
.Y(n_4710)
);

AO22x1_ASAP7_75t_L g4711 ( 
.A1(n_4655),
.A2(n_4645),
.B1(n_4635),
.B2(n_4607),
.Y(n_4711)
);

OAI211xp5_ASAP7_75t_L g4712 ( 
.A1(n_4665),
.A2(n_4678),
.B(n_4667),
.C(n_4657),
.Y(n_4712)
);

NOR2x1_ASAP7_75t_L g4713 ( 
.A(n_4675),
.B(n_4574),
.Y(n_4713)
);

OAI22xp33_ASAP7_75t_L g4714 ( 
.A1(n_4680),
.A2(n_4652),
.B1(n_4627),
.B2(n_4641),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4659),
.Y(n_4715)
);

BUFx2_ASAP7_75t_L g4716 ( 
.A(n_4672),
.Y(n_4716)
);

AOI21xp33_ASAP7_75t_L g4717 ( 
.A1(n_4662),
.A2(n_4621),
.B(n_4619),
.Y(n_4717)
);

AOI221xp5_ASAP7_75t_L g4718 ( 
.A1(n_4683),
.A2(n_4647),
.B1(n_4598),
.B2(n_4651),
.C(n_4583),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4653),
.Y(n_4719)
);

NOR2xp33_ASAP7_75t_L g4720 ( 
.A(n_4656),
.B(n_4570),
.Y(n_4720)
);

OAI211xp5_ASAP7_75t_SL g4721 ( 
.A1(n_4705),
.A2(n_4644),
.B(n_4584),
.C(n_4625),
.Y(n_4721)
);

NOR4xp75_ASAP7_75t_L g4722 ( 
.A(n_4676),
.B(n_4649),
.C(n_4640),
.D(n_4616),
.Y(n_4722)
);

CKINVDCx5p33_ASAP7_75t_R g4723 ( 
.A(n_4710),
.Y(n_4723)
);

OAI31xp33_ASAP7_75t_L g4724 ( 
.A1(n_4681),
.A2(n_4688),
.A3(n_4692),
.B(n_4666),
.Y(n_4724)
);

NOR3x1_ASAP7_75t_L g4725 ( 
.A(n_4685),
.B(n_4618),
.C(n_4576),
.Y(n_4725)
);

AOI221xp5_ASAP7_75t_L g4726 ( 
.A1(n_4707),
.A2(n_4642),
.B1(n_4603),
.B2(n_4630),
.C(n_778),
.Y(n_4726)
);

BUFx3_ASAP7_75t_L g4727 ( 
.A(n_4668),
.Y(n_4727)
);

A2O1A1Ixp33_ASAP7_75t_SL g4728 ( 
.A1(n_4668),
.A2(n_779),
.B(n_776),
.C(n_777),
.Y(n_4728)
);

AOI22xp33_ASAP7_75t_L g4729 ( 
.A1(n_4694),
.A2(n_783),
.B1(n_780),
.B2(n_782),
.Y(n_4729)
);

AOI211xp5_ASAP7_75t_L g4730 ( 
.A1(n_4690),
.A2(n_785),
.B(n_782),
.C(n_784),
.Y(n_4730)
);

AOI31xp33_ASAP7_75t_L g4731 ( 
.A1(n_4701),
.A2(n_791),
.A3(n_786),
.B(n_787),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4695),
.Y(n_4732)
);

XOR2x2_ASAP7_75t_L g4733 ( 
.A(n_4664),
.B(n_786),
.Y(n_4733)
);

AOI22xp5_ASAP7_75t_L g4734 ( 
.A1(n_4689),
.A2(n_4671),
.B1(n_4663),
.B2(n_4673),
.Y(n_4734)
);

AOI22xp33_ASAP7_75t_L g4735 ( 
.A1(n_4686),
.A2(n_793),
.B1(n_787),
.B2(n_792),
.Y(n_4735)
);

NAND3xp33_ASAP7_75t_L g4736 ( 
.A(n_4677),
.B(n_792),
.C(n_793),
.Y(n_4736)
);

OAI211xp5_ASAP7_75t_L g4737 ( 
.A1(n_4654),
.A2(n_796),
.B(n_794),
.C(n_795),
.Y(n_4737)
);

INVxp67_ASAP7_75t_L g4738 ( 
.A(n_4682),
.Y(n_4738)
);

OAI211xp5_ASAP7_75t_SL g4739 ( 
.A1(n_4684),
.A2(n_797),
.B(n_795),
.C(n_796),
.Y(n_4739)
);

AOI21xp33_ASAP7_75t_L g4740 ( 
.A1(n_4658),
.A2(n_798),
.B(n_799),
.Y(n_4740)
);

INVx3_ASAP7_75t_L g4741 ( 
.A(n_4660),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4699),
.B(n_799),
.Y(n_4742)
);

AOI22xp5_ASAP7_75t_L g4743 ( 
.A1(n_4706),
.A2(n_803),
.B1(n_801),
.B2(n_802),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4687),
.Y(n_4744)
);

AOI22xp33_ASAP7_75t_L g4745 ( 
.A1(n_4700),
.A2(n_807),
.B1(n_801),
.B2(n_804),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4727),
.Y(n_4746)
);

INVxp67_ASAP7_75t_L g4747 ( 
.A(n_4713),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4716),
.Y(n_4748)
);

OR2x2_ASAP7_75t_L g4749 ( 
.A(n_4741),
.B(n_4693),
.Y(n_4749)
);

NOR3xp33_ASAP7_75t_L g4750 ( 
.A(n_4712),
.B(n_4708),
.C(n_4704),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4741),
.B(n_4698),
.Y(n_4751)
);

NOR2xp67_ASAP7_75t_L g4752 ( 
.A(n_4737),
.B(n_4697),
.Y(n_4752)
);

NOR2xp33_ASAP7_75t_L g4753 ( 
.A(n_4721),
.B(n_4661),
.Y(n_4753)
);

NOR2x1_ASAP7_75t_L g4754 ( 
.A(n_4736),
.B(n_4679),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4731),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4733),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4732),
.Y(n_4757)
);

BUFx6f_ASAP7_75t_L g4758 ( 
.A(n_4715),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4723),
.Y(n_4759)
);

AO22x2_ASAP7_75t_L g4760 ( 
.A1(n_4719),
.A2(n_4669),
.B1(n_4670),
.B2(n_4703),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4720),
.Y(n_4761)
);

NOR2x1_ASAP7_75t_L g4762 ( 
.A(n_4739),
.B(n_4674),
.Y(n_4762)
);

NOR2x1_ASAP7_75t_L g4763 ( 
.A(n_4742),
.B(n_4691),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4748),
.Y(n_4764)
);

NOR2x1_ASAP7_75t_L g4765 ( 
.A(n_4755),
.B(n_4744),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4760),
.Y(n_4766)
);

INVx2_ASAP7_75t_L g4767 ( 
.A(n_4758),
.Y(n_4767)
);

HB1xp67_ASAP7_75t_L g4768 ( 
.A(n_4752),
.Y(n_4768)
);

NOR3xp33_ASAP7_75t_L g4769 ( 
.A(n_4747),
.B(n_4717),
.C(n_4738),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4760),
.Y(n_4770)
);

OR2x2_ASAP7_75t_L g4771 ( 
.A(n_4749),
.B(n_4745),
.Y(n_4771)
);

AND2x4_ASAP7_75t_L g4772 ( 
.A(n_4746),
.B(n_4734),
.Y(n_4772)
);

AOI22xp33_ASAP7_75t_R g4773 ( 
.A1(n_4757),
.A2(n_4722),
.B1(n_4724),
.B2(n_4725),
.Y(n_4773)
);

NOR2x1_ASAP7_75t_L g4774 ( 
.A(n_4751),
.B(n_4714),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4758),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4772),
.B(n_4711),
.Y(n_4776)
);

OAI21xp5_ASAP7_75t_SL g4777 ( 
.A1(n_4774),
.A2(n_4718),
.B(n_4753),
.Y(n_4777)
);

INVx1_ASAP7_75t_SL g4778 ( 
.A(n_4771),
.Y(n_4778)
);

OAI311xp33_ASAP7_75t_L g4779 ( 
.A1(n_4766),
.A2(n_4761),
.A3(n_4726),
.B1(n_4756),
.C1(n_4696),
.Y(n_4779)
);

AOI211xp5_ASAP7_75t_L g4780 ( 
.A1(n_4769),
.A2(n_4740),
.B(n_4750),
.C(n_4759),
.Y(n_4780)
);

AOI221xp5_ASAP7_75t_L g4781 ( 
.A1(n_4770),
.A2(n_4730),
.B1(n_4728),
.B2(n_4702),
.C(n_4735),
.Y(n_4781)
);

OAI221xp5_ASAP7_75t_SL g4782 ( 
.A1(n_4764),
.A2(n_4709),
.B1(n_4729),
.B2(n_4743),
.C(n_4762),
.Y(n_4782)
);

NAND4xp25_ASAP7_75t_L g4783 ( 
.A(n_4765),
.B(n_4754),
.C(n_4763),
.D(n_808),
.Y(n_4783)
);

NOR3xp33_ASAP7_75t_L g4784 ( 
.A(n_4768),
.B(n_804),
.C(n_807),
.Y(n_4784)
);

NAND4xp25_ASAP7_75t_L g4785 ( 
.A(n_4780),
.B(n_4775),
.C(n_4767),
.D(n_4773),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4776),
.Y(n_4786)
);

AND2x4_ASAP7_75t_L g4787 ( 
.A(n_4778),
.B(n_808),
.Y(n_4787)
);

OAI21xp5_ASAP7_75t_L g4788 ( 
.A1(n_4777),
.A2(n_809),
.B(n_811),
.Y(n_4788)
);

OAI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4788),
.A2(n_4783),
.B(n_4781),
.Y(n_4789)
);

BUFx2_ASAP7_75t_L g4790 ( 
.A(n_4787),
.Y(n_4790)
);

XNOR2xp5_ASAP7_75t_L g4791 ( 
.A(n_4785),
.B(n_4786),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4790),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4792),
.Y(n_4793)
);

AOI21xp5_ASAP7_75t_L g4794 ( 
.A1(n_4793),
.A2(n_4791),
.B(n_4779),
.Y(n_4794)
);

AOI22xp5_ASAP7_75t_L g4795 ( 
.A1(n_4794),
.A2(n_4784),
.B1(n_4789),
.B2(n_4782),
.Y(n_4795)
);

INVx2_ASAP7_75t_L g4796 ( 
.A(n_4795),
.Y(n_4796)
);

AOI22xp33_ASAP7_75t_L g4797 ( 
.A1(n_4796),
.A2(n_813),
.B1(n_809),
.B2(n_812),
.Y(n_4797)
);

AOI22xp5_ASAP7_75t_L g4798 ( 
.A1(n_4797),
.A2(n_815),
.B1(n_812),
.B2(n_814),
.Y(n_4798)
);

AOI22xp33_ASAP7_75t_L g4799 ( 
.A1(n_4797),
.A2(n_821),
.B1(n_814),
.B2(n_820),
.Y(n_4799)
);

OA22x2_ASAP7_75t_L g4800 ( 
.A1(n_4798),
.A2(n_822),
.B1(n_820),
.B2(n_821),
.Y(n_4800)
);

AO21x2_ASAP7_75t_L g4801 ( 
.A1(n_4799),
.A2(n_826),
.B(n_827),
.Y(n_4801)
);

AOI221xp5_ASAP7_75t_L g4802 ( 
.A1(n_4801),
.A2(n_828),
.B1(n_829),
.B2(n_830),
.C(n_831),
.Y(n_4802)
);

AOI211xp5_ASAP7_75t_L g4803 ( 
.A1(n_4802),
.A2(n_4800),
.B(n_832),
.C(n_831),
.Y(n_4803)
);


endmodule