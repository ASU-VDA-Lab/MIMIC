module fake_jpeg_11686_n_91 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx11_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_52),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_36),
.B1(n_31),
.B2(n_35),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_37),
.B1(n_12),
.B2(n_15),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_33),
.C(n_2),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_28),
.B1(n_26),
.B2(n_33),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_63),
.B1(n_37),
.B2(n_7),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_44),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_26),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_58),
.Y(n_71)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_5),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_5),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_76),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_66),
.B(n_62),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_6),
.B(n_8),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_10),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

XOR2x2_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_77),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_78),
.C(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_75),
.C(n_80),
.Y(n_87)
);

AOI31xp33_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_84),
.A3(n_82),
.B(n_73),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_82),
.C(n_73),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_11),
.C(n_19),
.Y(n_90)
);

XNOR2x2_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_21),
.Y(n_91)
);


endmodule