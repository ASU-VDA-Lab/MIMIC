module fake_netlist_5_685_n_1250 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1250);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1250;

wire n_924;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_659;
wire n_1182;
wire n_579;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_187;
wire n_1189;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_254;
wire n_1233;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_252;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_261;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_222;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_315;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_212;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_210;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_205;
wire n_1136;
wire n_754;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_202;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_522;
wire n_400;
wire n_930;
wire n_181;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_277;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_246;
wire n_1042;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_533;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_31),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_3),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_65),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_62),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_2),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_17),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_54),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_1),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_8),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_2),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_24),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_55),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_105),
.Y(n_193)
);

BUFx8_ASAP7_75t_SL g194 ( 
.A(n_78),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_161),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_101),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_136),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_144),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_116),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_3),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_66),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_43),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_85),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_47),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_75),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_53),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_12),
.Y(n_214)
);

BUFx8_ASAP7_75t_SL g215 ( 
.A(n_157),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_68),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_6),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_50),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_130),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_46),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_25),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_148),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_133),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_59),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_15),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_1),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_15),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_88),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_140),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_143),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_139),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_6),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_27),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_110),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_152),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_77),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_154),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_74),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_51),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_60),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_99),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_103),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_32),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_119),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_146),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_138),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_18),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_160),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_145),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_35),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_56),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_76),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_81),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_176),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_71),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_5),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_175),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_118),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_12),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_17),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_41),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_25),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_162),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_172),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_170),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_93),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_106),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_91),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_90),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_45),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_167),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_169),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_37),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_37),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_128),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_97),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_89),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_114),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_10),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_13),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_36),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_142),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_87),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_156),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_168),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_9),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_5),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_63),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_44),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_42),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_95),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_94),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_150),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_42),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_178),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_208),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_179),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_0),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_184),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_183),
.B(n_0),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_4),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_205),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_180),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_210),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_219),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_272),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_185),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_207),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_183),
.B(n_4),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_217),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_187),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_219),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_187),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_214),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_220),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_227),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_248),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_221),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_229),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_181),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_182),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_227),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_203),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_242),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_218),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_248),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_257),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_264),
.B(n_7),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_228),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_249),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_249),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_230),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_288),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_257),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_235),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_236),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_246),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_250),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_253),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_269),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_262),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_191),
.B(n_7),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_263),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_191),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_193),
.B(n_8),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_265),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_288),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_194),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_271),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_186),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_266),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_254),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_298),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_194),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_188),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_277),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_215),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_278),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_197),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_198),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_215),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_283),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_196),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_199),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_285),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_290),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_195),
.B(n_9),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_202),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_211),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_291),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_212),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_222),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_224),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_192),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_366),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_366),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_300),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_308),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_301),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_303),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_192),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_317),
.B(n_189),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

NAND2x1p5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_213),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_305),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_306),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_307),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_311),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_195),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_295),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_319),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_SL g412 ( 
.A(n_355),
.B(n_189),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_387),
.Y(n_413)
);

AND2x6_ASAP7_75t_L g414 ( 
.A(n_312),
.B(n_213),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_388),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_308),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_329),
.B(n_346),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_321),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_310),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_295),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_313),
.B(n_231),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_374),
.B(n_297),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_315),
.Y(n_432)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_358),
.B(n_231),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_389),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_302),
.B(n_226),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_309),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_299),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_381),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_357),
.B(n_260),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_332),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_389),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_368),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_333),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_323),
.B(n_234),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_325),
.A2(n_190),
.B1(n_293),
.B2(n_284),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_310),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_314),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_314),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_324),
.A2(n_190),
.B1(n_284),
.B2(n_293),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_316),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_316),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_378),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_326),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_326),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_337),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_335),
.B(n_297),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_337),
.B(n_237),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_391),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_419),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_390),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_318),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_419),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_325),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_427),
.C(n_435),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_439),
.B(n_425),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_433),
.A2(n_279),
.B1(n_213),
.B2(n_275),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_403),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_433),
.A2(n_279),
.B1(n_213),
.B2(n_275),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_391),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_447),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_427),
.B(n_341),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

OR2x6_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_455),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_391),
.Y(n_483)
);

AO22x1_ASAP7_75t_L g484 ( 
.A1(n_414),
.A2(n_255),
.B1(n_238),
.B2(n_239),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_425),
.B(n_379),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_421),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_341),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_407),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_394),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_438),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_390),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_398),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_414),
.A2(n_275),
.B1(n_279),
.B2(n_282),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_450),
.B(n_344),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_427),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_427),
.B(n_344),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_447),
.B(n_328),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_435),
.B(n_347),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_395),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_448),
.B(n_347),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_349),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_452),
.B(n_349),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_405),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_450),
.B(n_441),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_395),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_450),
.B(n_350),
.Y(n_516)
);

INVx6_ASAP7_75t_L g517 ( 
.A(n_427),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_405),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_392),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_412),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_405),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_427),
.B(n_350),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_392),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_424),
.B(n_351),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_435),
.B(n_351),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_405),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_450),
.B(n_352),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_424),
.B(n_352),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_R g530 ( 
.A(n_393),
.B(n_354),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_497),
.B(n_454),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_468),
.B(n_441),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_465),
.B(n_450),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_487),
.B(n_450),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_462),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_504),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_504),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_478),
.B(n_441),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_471),
.B(n_441),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_504),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_517),
.Y(n_541)
);

AO21x2_ASAP7_75t_L g542 ( 
.A1(n_467),
.A2(n_455),
.B(n_449),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_489),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_505),
.B(n_441),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_530),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_461),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_473),
.B(n_441),
.Y(n_547)
);

NOR2xp67_ASAP7_75t_L g548 ( 
.A(n_467),
.B(n_434),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_503),
.B(n_445),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_523),
.B(n_445),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_461),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_464),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_489),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_503),
.B(n_445),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_517),
.B(n_445),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_490),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_464),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_466),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_517),
.B(n_445),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_491),
.B(n_434),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_476),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_476),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_507),
.B(n_443),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_490),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_517),
.B(n_445),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_482),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_509),
.B(n_434),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_493),
.B(n_449),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_492),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_493),
.B(n_455),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_496),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_463),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_480),
.A2(n_442),
.B1(n_434),
.B2(n_456),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_480),
.A2(n_456),
.B1(n_457),
.B2(n_453),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_494),
.B(n_456),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_L g577 ( 
.A(n_500),
.B(n_414),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_480),
.A2(n_442),
.B1(n_457),
.B2(n_453),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_510),
.B(n_442),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_492),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_511),
.B(n_442),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_480),
.A2(n_414),
.B1(n_446),
.B2(n_459),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_507),
.B(n_453),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_482),
.Y(n_584)
);

O2A1O1Ixp5_ASAP7_75t_L g585 ( 
.A1(n_484),
.A2(n_513),
.B(n_494),
.C(n_499),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_495),
.B(n_499),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_525),
.B(n_457),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_495),
.B(n_429),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_529),
.B(n_429),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_480),
.B(n_414),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_526),
.B(n_453),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_526),
.B(n_443),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_469),
.B(n_414),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_521),
.A2(n_446),
.B1(n_459),
.B2(n_414),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_469),
.B(n_443),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_488),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_502),
.B(n_393),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_479),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_342),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_516),
.B(n_459),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_469),
.B(n_459),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_469),
.B(n_431),
.Y(n_604)
);

A2O1A1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_488),
.A2(n_446),
.B(n_444),
.C(n_440),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_481),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_521),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_519),
.B(n_254),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_496),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_528),
.B(n_431),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_506),
.Y(n_612)
);

OAI221xp5_ASAP7_75t_L g613 ( 
.A1(n_481),
.A2(n_396),
.B1(n_406),
.B2(n_420),
.C(n_423),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_484),
.A2(n_446),
.B1(n_444),
.B2(n_413),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_501),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_475),
.B(n_422),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_498),
.B(n_440),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g618 ( 
.A(n_506),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_498),
.B(n_426),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_498),
.B(n_426),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_498),
.B(n_437),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_470),
.B(n_422),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_520),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_512),
.B(n_437),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_519),
.B(n_428),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_512),
.B(n_405),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_527),
.B(n_416),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_527),
.B(n_416),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_514),
.B(n_416),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_519),
.B(n_428),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_587),
.A2(n_343),
.B1(n_345),
.B2(n_334),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_564),
.B(n_432),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_532),
.A2(n_519),
.B(n_486),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_590),
.B(n_458),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_560),
.B(n_458),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_604),
.A2(n_519),
.B(n_486),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_539),
.A2(n_361),
.B1(n_519),
.B2(n_399),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_577),
.A2(n_547),
.B(n_617),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_546),
.Y(n_641)
);

O2A1O1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_594),
.A2(n_396),
.B(n_406),
.C(n_399),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_577),
.A2(n_486),
.B(n_470),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_568),
.B(n_514),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_585),
.A2(n_522),
.B(n_518),
.Y(n_645)
);

BUFx12f_ASAP7_75t_L g646 ( 
.A(n_545),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_573),
.B(n_397),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_548),
.A2(n_522),
.B(n_518),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_579),
.B(n_581),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_549),
.A2(n_486),
.B(n_470),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_534),
.A2(n_470),
.B1(n_413),
.B2(n_520),
.Y(n_651)
);

O2A1O1Ixp5_ASAP7_75t_L g652 ( 
.A1(n_533),
.A2(n_524),
.B(n_404),
.C(n_413),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_548),
.A2(n_399),
.B1(n_524),
.B2(n_268),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_538),
.A2(n_485),
.B(n_483),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_544),
.A2(n_485),
.B(n_483),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_545),
.B(n_397),
.Y(n_656)
);

AO21x1_ASAP7_75t_L g657 ( 
.A1(n_575),
.A2(n_399),
.B(n_270),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_554),
.A2(n_477),
.B(n_462),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_541),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_564),
.B(n_420),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_608),
.B(n_354),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_550),
.A2(n_474),
.B(n_460),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_603),
.A2(n_477),
.B(n_462),
.Y(n_663)
);

NOR2xp67_ASAP7_75t_L g664 ( 
.A(n_599),
.B(n_613),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_589),
.B(n_432),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_583),
.A2(n_413),
.B1(n_356),
.B2(n_385),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_622),
.B(n_432),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_592),
.B(n_362),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_616),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_569),
.B(n_462),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_578),
.B(n_574),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_611),
.B(n_369),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_591),
.A2(n_474),
.B(n_460),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_541),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_571),
.B(n_462),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_610),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_555),
.A2(n_566),
.B(n_559),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_601),
.B(n_356),
.Y(n_678)
);

AOI21x1_ASAP7_75t_L g679 ( 
.A1(n_595),
.A2(n_474),
.B(n_460),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_535),
.A2(n_477),
.B(n_462),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_582),
.B(n_360),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_576),
.A2(n_477),
.B(n_508),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_586),
.B(n_477),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_546),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_535),
.A2(n_477),
.B(n_508),
.Y(n_685)
);

OR2x6_ASAP7_75t_L g686 ( 
.A(n_601),
.B(n_451),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_602),
.B(n_531),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_605),
.B(n_360),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_535),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_597),
.B(n_365),
.Y(n_690)
);

O2A1O1Ixp5_ASAP7_75t_L g691 ( 
.A1(n_621),
.A2(n_404),
.B(n_280),
.C(n_296),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_536),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_537),
.A2(n_287),
.B(n_245),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_535),
.A2(n_515),
.B(n_508),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_542),
.B(n_365),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_537),
.A2(n_423),
.B(n_404),
.Y(n_696)
);

AND2x2_ASAP7_75t_SL g697 ( 
.A(n_612),
.B(n_451),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_542),
.B(n_371),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_614),
.B(n_371),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_610),
.Y(n_700)
);

OR2x2_ASAP7_75t_SL g701 ( 
.A(n_618),
.B(n_372),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_542),
.B(n_373),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_624),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_551),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_614),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_625),
.B(n_373),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_540),
.B(n_377),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_596),
.A2(n_430),
.B(n_404),
.C(n_377),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_624),
.Y(n_709)
);

AO21x1_ASAP7_75t_L g710 ( 
.A1(n_551),
.A2(n_430),
.B(n_409),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_619),
.A2(n_515),
.B(n_508),
.Y(n_711)
);

AND2x4_ASAP7_75t_SL g712 ( 
.A(n_596),
.B(n_376),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_620),
.A2(n_515),
.B(n_508),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_626),
.B(n_380),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_540),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_615),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_552),
.B(n_380),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_552),
.B(n_385),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_557),
.B(n_430),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_631),
.B(n_436),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_557),
.A2(n_430),
.B1(n_200),
.B2(n_267),
.Y(n_721)
);

OR2x6_ASAP7_75t_SL g722 ( 
.A(n_615),
.B(n_201),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_558),
.B(n_416),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_627),
.A2(n_515),
.B(n_508),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_623),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_628),
.A2(n_515),
.B(n_416),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_572),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_572),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_558),
.B(n_416),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_629),
.A2(n_515),
.B(n_418),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_561),
.B(n_436),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_561),
.B(n_408),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_703),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_SL g734 ( 
.A(n_646),
.B(n_535),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_649),
.A2(n_562),
.B1(n_563),
.B2(n_567),
.Y(n_735)
);

BUFx8_ASAP7_75t_L g736 ( 
.A(n_661),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_664),
.A2(n_562),
.B1(n_563),
.B2(n_567),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_635),
.A2(n_598),
.B(n_584),
.C(n_572),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_703),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_660),
.B(n_623),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_703),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_669),
.B(n_636),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_641),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_642),
.A2(n_598),
.B(n_584),
.C(n_565),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_647),
.B(n_543),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_687),
.A2(n_556),
.B(n_543),
.C(n_580),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_632),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_722),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_633),
.B(n_408),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_705),
.A2(n_553),
.B1(n_556),
.B2(n_565),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_720),
.A2(n_570),
.B(n_553),
.C(n_580),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_684),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_695),
.A2(n_570),
.B(n_607),
.C(n_606),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_732),
.B(n_606),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_648),
.A2(n_630),
.B(n_609),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_704),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_714),
.A2(n_607),
.B1(n_609),
.B2(n_204),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_671),
.A2(n_535),
.B(n_600),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_659),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_706),
.B(n_588),
.Y(n_760)
);

BUFx12f_ASAP7_75t_L g761 ( 
.A(n_701),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_715),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_665),
.B(n_588),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_640),
.A2(n_600),
.B(n_593),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_717),
.B(n_718),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_660),
.B(n_593),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_707),
.B(n_690),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_698),
.A2(n_410),
.B(n_417),
.C(n_415),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_700),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_656),
.B(n_409),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_668),
.B(n_410),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_725),
.B(n_418),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_731),
.B(n_418),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_659),
.B(n_411),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_678),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_SL g776 ( 
.A(n_697),
.B(n_260),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_SL g777 ( 
.A(n_676),
.B(n_275),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_SL g778 ( 
.A(n_672),
.B(n_260),
.Y(n_778)
);

O2A1O1Ixp5_ASAP7_75t_L g779 ( 
.A1(n_657),
.A2(n_417),
.B(n_415),
.C(n_411),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_640),
.A2(n_279),
.B(n_401),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_708),
.A2(n_252),
.B(n_209),
.C(n_216),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_639),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_683),
.A2(n_402),
.B(n_401),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_709),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_692),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_712),
.B(n_286),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_699),
.B(n_206),
.C(n_223),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_702),
.A2(n_258),
.B(n_232),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_676),
.B(n_225),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_681),
.A2(n_254),
.B1(n_286),
.B2(n_233),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_686),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_667),
.B(n_240),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_643),
.A2(n_402),
.B(n_401),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_644),
.A2(n_273),
.B1(n_243),
.B2(n_244),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_666),
.B(n_286),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_688),
.A2(n_276),
.B1(n_247),
.B2(n_251),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_643),
.A2(n_289),
.B(n_256),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_670),
.A2(n_402),
.B(n_401),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_SL g799 ( 
.A1(n_781),
.A2(n_693),
.B(n_638),
.C(n_716),
.Y(n_799)
);

OAI21x1_ASAP7_75t_L g800 ( 
.A1(n_764),
.A2(n_677),
.B(n_679),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_761),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_743),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_736),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_733),
.Y(n_804)
);

NOR2xp67_ASAP7_75t_L g805 ( 
.A(n_775),
.B(n_674),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_778),
.A2(n_686),
.B(n_721),
.C(n_719),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_774),
.B(n_741),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_764),
.A2(n_663),
.B(n_662),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_770),
.B(n_674),
.Y(n_809)
);

BUFx12f_ASAP7_75t_L g810 ( 
.A(n_736),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_759),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_752),
.Y(n_812)
);

OA21x2_ASAP7_75t_L g813 ( 
.A1(n_779),
.A2(n_710),
.B(n_645),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_755),
.A2(n_691),
.B(n_673),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_742),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_754),
.A2(n_686),
.B1(n_696),
.B2(n_651),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_755),
.A2(n_675),
.B(n_634),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_760),
.B(n_727),
.Y(n_818)
);

AO32x2_ASAP7_75t_L g819 ( 
.A1(n_750),
.A2(n_653),
.A3(n_652),
.B1(n_730),
.B2(n_682),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_756),
.Y(n_820)
);

AO31x2_ASAP7_75t_L g821 ( 
.A1(n_744),
.A2(n_682),
.A3(n_711),
.B(n_713),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_771),
.B(n_727),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_793),
.A2(n_724),
.B(n_654),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_747),
.B(n_728),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_765),
.B(n_728),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_745),
.B(n_241),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_767),
.A2(n_634),
.B(n_650),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_758),
.A2(n_689),
.B(n_637),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_780),
.A2(n_730),
.B(n_655),
.Y(n_829)
);

OAI21x1_ASAP7_75t_L g830 ( 
.A1(n_798),
.A2(n_658),
.B(n_713),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_776),
.B(n_689),
.Y(n_831)
);

AO31x2_ASAP7_75t_L g832 ( 
.A1(n_738),
.A2(n_711),
.A3(n_726),
.B(n_723),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_733),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_749),
.B(n_729),
.Y(n_834)
);

NAND2x1p5_ASAP7_75t_L g835 ( 
.A(n_741),
.B(n_726),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_798),
.A2(n_637),
.B(n_680),
.Y(n_836)
);

NOR4xp25_ASAP7_75t_L g837 ( 
.A(n_768),
.B(n_10),
.C(n_11),
.D(n_13),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_786),
.B(n_261),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_795),
.A2(n_694),
.B(n_685),
.C(n_281),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_748),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_780),
.A2(n_292),
.B(n_254),
.Y(n_841)
);

INVx6_ASAP7_75t_L g842 ( 
.A(n_733),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_785),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_773),
.A2(n_402),
.B(n_401),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_SL g845 ( 
.A(n_788),
.B(n_254),
.C(n_14),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_783),
.A2(n_254),
.B(n_96),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_768),
.A2(n_254),
.B(n_401),
.C(n_400),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_753),
.A2(n_751),
.B(n_735),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_791),
.A2(n_402),
.B1(n_400),
.B2(n_395),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_769),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_783),
.A2(n_92),
.B(n_174),
.Y(n_851)
);

OAI21x1_ASAP7_75t_L g852 ( 
.A1(n_753),
.A2(n_86),
.B(n_173),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_804),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_SL g854 ( 
.A1(n_826),
.A2(n_797),
.B1(n_774),
.B2(n_792),
.Y(n_854)
);

OAI22xp33_ASAP7_75t_L g855 ( 
.A1(n_815),
.A2(n_772),
.B1(n_762),
.B2(n_766),
.Y(n_855)
);

CKINVDCx6p67_ASAP7_75t_R g856 ( 
.A(n_810),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_824),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_822),
.B(n_740),
.Y(n_858)
);

BUFx8_ASAP7_75t_L g859 ( 
.A(n_803),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_842),
.Y(n_860)
);

INVx6_ASAP7_75t_L g861 ( 
.A(n_811),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_802),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_812),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_842),
.Y(n_864)
);

BUFx10_ASAP7_75t_L g865 ( 
.A(n_801),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_806),
.B(n_737),
.Y(n_866)
);

CKINVDCx6p67_ASAP7_75t_R g867 ( 
.A(n_833),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_833),
.Y(n_868)
);

BUFx4f_ASAP7_75t_SL g869 ( 
.A(n_840),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_820),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_838),
.B(n_740),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_845),
.A2(n_787),
.B1(n_790),
.B2(n_784),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_833),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_821),
.Y(n_874)
);

AOI22x1_ASAP7_75t_SL g875 ( 
.A1(n_811),
.A2(n_782),
.B1(n_734),
.B2(n_16),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_843),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_825),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_840),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_850),
.Y(n_879)
);

INVx6_ASAP7_75t_L g880 ( 
.A(n_807),
.Y(n_880)
);

BUFx2_ASAP7_75t_R g881 ( 
.A(n_831),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_818),
.Y(n_882)
);

BUFx12f_ASAP7_75t_L g883 ( 
.A(n_807),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_809),
.B(n_794),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_817),
.A2(n_746),
.B(n_757),
.Y(n_885)
);

BUFx4f_ASAP7_75t_SL g886 ( 
.A(n_805),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_816),
.A2(n_763),
.B1(n_796),
.B2(n_789),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_816),
.A2(n_759),
.B1(n_739),
.B2(n_777),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_821),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_821),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_834),
.B(n_739),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_834),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_818),
.Y(n_893)
);

OAI21xp33_ASAP7_75t_L g894 ( 
.A1(n_837),
.A2(n_759),
.B(n_739),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_835),
.Y(n_895)
);

INVx6_ASAP7_75t_L g896 ( 
.A(n_835),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_851),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_849),
.A2(n_402),
.B1(n_400),
.B2(n_395),
.Y(n_898)
);

BUFx4f_ASAP7_75t_SL g899 ( 
.A(n_837),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_841),
.B(n_11),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_848),
.A2(n_400),
.B1(n_395),
.B2(n_18),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_SL g902 ( 
.A1(n_848),
.A2(n_14),
.B(n_16),
.Y(n_902)
);

CKINVDCx6p67_ASAP7_75t_R g903 ( 
.A(n_839),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_813),
.Y(n_904)
);

BUFx12f_ASAP7_75t_L g905 ( 
.A(n_799),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_827),
.B(n_19),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_846),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_814),
.A2(n_813),
.B1(n_829),
.B2(n_852),
.Y(n_908)
);

BUFx4f_ASAP7_75t_SL g909 ( 
.A(n_847),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_814),
.A2(n_400),
.B1(n_20),
.B2(n_21),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_827),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_874),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_889),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_878),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_874),
.B(n_817),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_885),
.A2(n_836),
.B(n_830),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_889),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_877),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_890),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_890),
.B(n_829),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_907),
.Y(n_921)
);

OAI21x1_ASAP7_75t_L g922 ( 
.A1(n_908),
.A2(n_800),
.B(n_823),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_882),
.B(n_832),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_863),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_863),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_904),
.B(n_832),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_870),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_908),
.B(n_893),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_906),
.A2(n_828),
.B(n_808),
.Y(n_929)
);

AO21x2_ASAP7_75t_L g930 ( 
.A1(n_900),
.A2(n_844),
.B(n_819),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_870),
.Y(n_931)
);

INVx5_ASAP7_75t_SL g932 ( 
.A(n_903),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_862),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_876),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_897),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_897),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_895),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_897),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_897),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_894),
.B(n_832),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_899),
.Y(n_941)
);

BUFx2_ASAP7_75t_SL g942 ( 
.A(n_888),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_896),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_887),
.A2(n_819),
.B(n_100),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_896),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_896),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_899),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_910),
.B(n_819),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_905),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_944),
.A2(n_866),
.B(n_902),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_947),
.A2(n_866),
.B(n_911),
.C(n_910),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_926),
.B(n_887),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_926),
.B(n_857),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_926),
.B(n_901),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_920),
.B(n_901),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_915),
.B(n_891),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_921),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_938),
.B(n_868),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_933),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_938),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_943),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_921),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_924),
.B(n_855),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_938),
.B(n_935),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_941),
.A2(n_892),
.B1(n_854),
.B2(n_872),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_920),
.B(n_879),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_924),
.B(n_855),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_938),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_921),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_920),
.B(n_884),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_941),
.A2(n_909),
.B1(n_871),
.B2(n_872),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_940),
.B(n_853),
.Y(n_972)
);

AO32x2_ASAP7_75t_L g973 ( 
.A1(n_943),
.A2(n_898),
.A3(n_873),
.B1(n_864),
.B2(n_909),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_915),
.B(n_858),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_928),
.B(n_881),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_933),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_940),
.B(n_22),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_940),
.B(n_22),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_914),
.B(n_860),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_915),
.B(n_873),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_914),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_928),
.B(n_23),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_935),
.B(n_57),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_935),
.B(n_58),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_918),
.Y(n_985)
);

NAND2xp33_ASAP7_75t_R g986 ( 
.A(n_941),
.B(n_875),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_918),
.Y(n_987)
);

AO21x2_ASAP7_75t_L g988 ( 
.A1(n_922),
.A2(n_867),
.B(n_24),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_933),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_934),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_970),
.B(n_928),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_960),
.B(n_936),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_960),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_960),
.B(n_919),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_970),
.B(n_923),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_962),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_960),
.B(n_919),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_964),
.B(n_936),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_962),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_964),
.B(n_936),
.Y(n_1000)
);

AOI222xp33_ASAP7_75t_SL g1001 ( 
.A1(n_950),
.A2(n_947),
.B1(n_934),
.B2(n_27),
.C1(n_28),
.C2(n_29),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_964),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_962),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_970),
.B(n_923),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_961),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_964),
.B(n_919),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_965),
.A2(n_947),
.B1(n_948),
.B2(n_942),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_964),
.B(n_968),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_987),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_969),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_969),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_969),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_990),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_957),
.Y(n_1014)
);

OAI222xp33_ASAP7_75t_L g1015 ( 
.A1(n_965),
.A2(n_947),
.B1(n_948),
.B2(n_934),
.C1(n_925),
.C2(n_927),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_968),
.B(n_912),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_1009),
.B(n_981),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_1016),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1002),
.B(n_972),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_1009),
.B(n_985),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_996),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_1005),
.B(n_950),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_996),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_991),
.B(n_995),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1014),
.Y(n_1025)
);

OAI33xp33_ASAP7_75t_L g1026 ( 
.A1(n_1001),
.A2(n_959),
.A3(n_989),
.B1(n_976),
.B2(n_990),
.B3(n_974),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_996),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_991),
.B(n_966),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_996),
.Y(n_1029)
);

NOR2x1_ASAP7_75t_L g1030 ( 
.A(n_1005),
.B(n_988),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1014),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1002),
.B(n_972),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1002),
.B(n_972),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_995),
.B(n_974),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1007),
.A2(n_954),
.B1(n_952),
.B2(n_971),
.Y(n_1035)
);

AOI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_1015),
.A2(n_951),
.B1(n_952),
.B2(n_982),
.C(n_966),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1008),
.B(n_953),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1014),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_1031),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1024),
.B(n_953),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_1018),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1025),
.Y(n_1042)
);

AND2x2_ASAP7_75t_SL g1043 ( 
.A(n_1036),
.B(n_1001),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_1030),
.B(n_992),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1034),
.B(n_1004),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1026),
.A2(n_986),
.B1(n_1007),
.B2(n_954),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1019),
.B(n_1008),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1021),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_1030),
.B(n_992),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1025),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_1045),
.B(n_1034),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1042),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1042),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1050),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1050),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1045),
.B(n_1024),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_1039),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1052),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1053),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_L g1060 ( 
.A(n_1054),
.B(n_1044),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1056),
.B(n_1043),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_1061),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_1060),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1058),
.B(n_1051),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1059),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_1061),
.A2(n_1043),
.B1(n_1046),
.B2(n_1022),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_1061),
.B(n_1040),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_1061),
.A2(n_1043),
.B(n_1022),
.C(n_1057),
.Y(n_1068)
);

AOI221xp5_ASAP7_75t_L g1069 ( 
.A1(n_1061),
.A2(n_1046),
.B1(n_1055),
.B2(n_1049),
.C(n_1044),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1061),
.B(n_1047),
.Y(n_1070)
);

OAI322xp33_ASAP7_75t_L g1071 ( 
.A1(n_1061),
.A2(n_1057),
.A3(n_1041),
.B1(n_1017),
.B2(n_1020),
.C1(n_978),
.C2(n_977),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_L g1072 ( 
.A(n_1061),
.B(n_1044),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1066),
.A2(n_1022),
.B1(n_1035),
.B2(n_975),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1065),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1064),
.Y(n_1075)
);

OAI32xp33_ASAP7_75t_L g1076 ( 
.A1(n_1063),
.A2(n_977),
.A3(n_978),
.B1(n_975),
.B2(n_982),
.Y(n_1076)
);

OAI31xp33_ASAP7_75t_L g1077 ( 
.A1(n_1068),
.A2(n_1049),
.A3(n_1044),
.B(n_1015),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_1062),
.B(n_1028),
.Y(n_1078)
);

OAI21xp33_ASAP7_75t_SL g1079 ( 
.A1(n_1069),
.A2(n_1047),
.B(n_1022),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1071),
.A2(n_1049),
.B(n_979),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1070),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1072),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1072),
.A2(n_1022),
.B1(n_1049),
.B2(n_982),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1067),
.B(n_1039),
.Y(n_1084)
);

OAI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_1069),
.A2(n_951),
.B1(n_1028),
.B2(n_953),
.C(n_1048),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1070),
.B(n_856),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1065),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_1069),
.A2(n_952),
.B(n_978),
.C(n_977),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1075),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1086),
.B(n_865),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1081),
.B(n_1039),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1074),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1087),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1082),
.B(n_865),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1080),
.B(n_1037),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_1084),
.B(n_1048),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1078),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1083),
.B(n_1037),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1088),
.B(n_1019),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_SL g1100 ( 
.A1(n_1077),
.A2(n_869),
.B(n_954),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_SL g1101 ( 
.A1(n_1073),
.A2(n_1085),
.B1(n_1079),
.B2(n_1076),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1073),
.B(n_869),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1084),
.B(n_1032),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1075),
.B(n_1032),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1075),
.Y(n_1105)
);

XNOR2xp5_ASAP7_75t_L g1106 ( 
.A(n_1086),
.B(n_966),
.Y(n_1106)
);

XNOR2x1_ASAP7_75t_L g1107 ( 
.A(n_1073),
.B(n_23),
.Y(n_1107)
);

NAND2x1_ASAP7_75t_L g1108 ( 
.A(n_1097),
.B(n_1094),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1090),
.Y(n_1109)
);

AOI221xp5_ASAP7_75t_SL g1110 ( 
.A1(n_1102),
.A2(n_1033),
.B1(n_949),
.B2(n_942),
.C(n_1038),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_1107),
.B(n_859),
.C(n_983),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1097),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1089),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_1107),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1102),
.A2(n_988),
.B(n_984),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1105),
.Y(n_1116)
);

NAND4xp25_ASAP7_75t_L g1117 ( 
.A(n_1101),
.B(n_859),
.C(n_983),
.D(n_984),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_L g1118 ( 
.A(n_1100),
.B(n_984),
.C(n_983),
.Y(n_1118)
);

NOR2x1_ASAP7_75t_L g1119 ( 
.A(n_1092),
.B(n_988),
.Y(n_1119)
);

NOR2x1_ASAP7_75t_SL g1120 ( 
.A(n_1093),
.B(n_949),
.Y(n_1120)
);

BUFx8_ASAP7_75t_SL g1121 ( 
.A(n_1104),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1095),
.B(n_1033),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_SL g1123 ( 
.A(n_1101),
.B(n_1091),
.C(n_1099),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1098),
.A2(n_932),
.B1(n_988),
.B2(n_942),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_1112),
.A2(n_1103),
.B(n_1106),
.C(n_1096),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1114),
.A2(n_1096),
.B(n_984),
.Y(n_1126)
);

OAI211xp5_ASAP7_75t_SL g1127 ( 
.A1(n_1109),
.A2(n_1096),
.B(n_28),
.C(n_29),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1113),
.Y(n_1128)
);

OA211x2_ASAP7_75t_L g1129 ( 
.A1(n_1108),
.A2(n_886),
.B(n_932),
.C(n_31),
.Y(n_1129)
);

AND4x1_ASAP7_75t_L g1130 ( 
.A(n_1111),
.B(n_886),
.C(n_30),
.D(n_32),
.Y(n_1130)
);

AOI211xp5_ASAP7_75t_L g1131 ( 
.A1(n_1117),
.A2(n_983),
.B(n_984),
.C(n_949),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1117),
.A2(n_983),
.B1(n_1038),
.B2(n_948),
.C(n_946),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_1121),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1120),
.A2(n_1116),
.B(n_1123),
.Y(n_1134)
);

OAI211xp5_ASAP7_75t_SL g1135 ( 
.A1(n_1122),
.A2(n_26),
.B(n_30),
.C(n_33),
.Y(n_1135)
);

NOR2x1_ASAP7_75t_L g1136 ( 
.A(n_1119),
.B(n_26),
.Y(n_1136)
);

AOI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1115),
.A2(n_1110),
.B1(n_1124),
.B2(n_1118),
.C(n_946),
.Y(n_1137)
);

AOI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_1114),
.A2(n_33),
.B(n_34),
.Y(n_1138)
);

AOI211xp5_ASAP7_75t_L g1139 ( 
.A1(n_1117),
.A2(n_949),
.B(n_35),
.C(n_36),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1114),
.A2(n_1021),
.B(n_1029),
.Y(n_1140)
);

AOI211xp5_ASAP7_75t_L g1141 ( 
.A1(n_1117),
.A2(n_949),
.B(n_38),
.C(n_39),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1114),
.A2(n_944),
.B(n_949),
.C(n_1005),
.Y(n_1142)
);

OAI321xp33_ASAP7_75t_L g1143 ( 
.A1(n_1117),
.A2(n_949),
.A3(n_946),
.B1(n_945),
.B2(n_967),
.C(n_963),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1114),
.A2(n_932),
.B1(n_949),
.B2(n_998),
.Y(n_1144)
);

AOI221xp5_ASAP7_75t_L g1145 ( 
.A1(n_1117),
.A2(n_945),
.B1(n_1031),
.B2(n_949),
.C(n_1023),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_R g1146 ( 
.A(n_1112),
.B(n_34),
.Y(n_1146)
);

OAI31xp33_ASAP7_75t_L g1147 ( 
.A1(n_1117),
.A2(n_1005),
.A3(n_932),
.B(n_961),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1114),
.A2(n_932),
.B1(n_1027),
.B2(n_1023),
.Y(n_1148)
);

O2A1O1Ixp5_ASAP7_75t_SL g1149 ( 
.A1(n_1128),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1136),
.Y(n_1150)
);

AOI222xp33_ASAP7_75t_L g1151 ( 
.A1(n_1126),
.A2(n_932),
.B1(n_955),
.B2(n_944),
.C1(n_44),
.C2(n_45),
.Y(n_1151)
);

AOI221x1_ASAP7_75t_L g1152 ( 
.A1(n_1134),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.C(n_46),
.Y(n_1152)
);

NOR2x1_ASAP7_75t_L g1153 ( 
.A(n_1127),
.B(n_47),
.Y(n_1153)
);

OAI211xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1133),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1125),
.A2(n_48),
.B(n_51),
.C(n_52),
.Y(n_1155)
);

AOI222xp33_ASAP7_75t_L g1156 ( 
.A1(n_1137),
.A2(n_932),
.B1(n_955),
.B2(n_944),
.C1(n_52),
.C2(n_967),
.Y(n_1156)
);

NAND4xp25_ASAP7_75t_L g1157 ( 
.A(n_1139),
.B(n_1004),
.C(n_980),
.D(n_956),
.Y(n_1157)
);

AOI211xp5_ASAP7_75t_SL g1158 ( 
.A1(n_1138),
.A2(n_945),
.B(n_963),
.C(n_959),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1135),
.A2(n_943),
.B(n_1027),
.C(n_1029),
.Y(n_1159)
);

AOI211xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1141),
.A2(n_1016),
.B(n_980),
.C(n_939),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_1146),
.Y(n_1161)
);

AOI21xp33_ASAP7_75t_SL g1162 ( 
.A1(n_1147),
.A2(n_61),
.B(n_64),
.Y(n_1162)
);

OAI221xp5_ASAP7_75t_L g1163 ( 
.A1(n_1131),
.A2(n_880),
.B1(n_861),
.B2(n_943),
.C(n_961),
.Y(n_1163)
);

AOI211xp5_ASAP7_75t_L g1164 ( 
.A1(n_1148),
.A2(n_956),
.B(n_939),
.C(n_955),
.Y(n_1164)
);

AOI211xp5_ASAP7_75t_L g1165 ( 
.A1(n_1145),
.A2(n_939),
.B(n_958),
.C(n_1016),
.Y(n_1165)
);

AOI222xp33_ASAP7_75t_L g1166 ( 
.A1(n_1132),
.A2(n_993),
.B1(n_1008),
.B2(n_998),
.C1(n_1000),
.C2(n_883),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1143),
.A2(n_1142),
.B1(n_1140),
.B2(n_1144),
.C(n_1129),
.Y(n_1167)
);

AOI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1130),
.A2(n_958),
.B1(n_998),
.B2(n_1000),
.C(n_1008),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1133),
.A2(n_998),
.B1(n_1000),
.B2(n_861),
.Y(n_1169)
);

AOI211xp5_ASAP7_75t_L g1170 ( 
.A1(n_1134),
.A2(n_958),
.B(n_1000),
.C(n_998),
.Y(n_1170)
);

AOI221x1_ASAP7_75t_L g1171 ( 
.A1(n_1134),
.A2(n_1013),
.B1(n_1012),
.B2(n_1010),
.C(n_999),
.Y(n_1171)
);

AOI222xp33_ASAP7_75t_L g1172 ( 
.A1(n_1126),
.A2(n_993),
.B1(n_1008),
.B2(n_1000),
.C1(n_1013),
.C2(n_1012),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1161),
.B(n_1150),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_SL g1174 ( 
.A1(n_1153),
.A2(n_861),
.B1(n_880),
.B2(n_993),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1160),
.B(n_1170),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1163),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1152),
.B(n_958),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1171),
.Y(n_1178)
);

NAND2xp33_ASAP7_75t_L g1179 ( 
.A(n_1167),
.B(n_1003),
.Y(n_1179)
);

XNOR2xp5_ASAP7_75t_L g1180 ( 
.A(n_1157),
.B(n_67),
.Y(n_1180)
);

NOR2x1_ASAP7_75t_L g1181 ( 
.A(n_1154),
.B(n_976),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1155),
.B(n_1003),
.Y(n_1182)
);

XNOR2x1_ASAP7_75t_L g1183 ( 
.A(n_1169),
.B(n_70),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_L g1184 ( 
.A(n_1159),
.B(n_989),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1156),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1158),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_L g1187 ( 
.A(n_1149),
.B(n_999),
.Y(n_1187)
);

NAND4xp75_ASAP7_75t_L g1188 ( 
.A(n_1168),
.B(n_968),
.C(n_1010),
.D(n_997),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1162),
.B(n_958),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1151),
.Y(n_1190)
);

XOR2xp5_ASAP7_75t_L g1191 ( 
.A(n_1166),
.B(n_72),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1164),
.Y(n_1192)
);

NOR2x1_ASAP7_75t_L g1193 ( 
.A(n_1165),
.B(n_957),
.Y(n_1193)
);

INVxp33_ASAP7_75t_SL g1194 ( 
.A(n_1172),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1177),
.B(n_1011),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1177),
.B(n_1011),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1173),
.B(n_1006),
.Y(n_1197)
);

AOI21xp33_ASAP7_75t_SL g1198 ( 
.A1(n_1174),
.A2(n_73),
.B(n_79),
.Y(n_1198)
);

AOI21xp33_ASAP7_75t_L g1199 ( 
.A1(n_1179),
.A2(n_80),
.B(n_82),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1182),
.B(n_1006),
.Y(n_1200)
);

NOR3xp33_ASAP7_75t_L g1201 ( 
.A(n_1185),
.B(n_1190),
.C(n_1176),
.Y(n_1201)
);

NOR4xp25_ASAP7_75t_L g1202 ( 
.A(n_1192),
.B(n_927),
.C(n_925),
.D(n_1006),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1175),
.B(n_997),
.Y(n_1203)
);

AOI21xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1194),
.A2(n_83),
.B(n_84),
.Y(n_1204)
);

OA22x2_ASAP7_75t_L g1205 ( 
.A1(n_1191),
.A2(n_937),
.B1(n_994),
.B2(n_997),
.Y(n_1205)
);

AOI211x1_ASAP7_75t_L g1206 ( 
.A1(n_1187),
.A2(n_1183),
.B(n_1181),
.C(n_1189),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1178),
.A2(n_937),
.B(n_929),
.C(n_925),
.Y(n_1207)
);

NOR3xp33_ASAP7_75t_SL g1208 ( 
.A(n_1180),
.B(n_98),
.C(n_102),
.Y(n_1208)
);

NOR3xp33_ASAP7_75t_L g1209 ( 
.A(n_1186),
.B(n_929),
.C(n_916),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1206),
.B(n_1178),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_L g1211 ( 
.A1(n_1199),
.A2(n_1188),
.B1(n_1184),
.B2(n_1193),
.C(n_937),
.Y(n_1211)
);

XNOR2x1_ASAP7_75t_L g1212 ( 
.A(n_1205),
.B(n_104),
.Y(n_1212)
);

XOR2xp5_ASAP7_75t_L g1213 ( 
.A(n_1197),
.B(n_107),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1201),
.A2(n_880),
.B1(n_994),
.B2(n_930),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1196),
.B(n_927),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_SL g1216 ( 
.A(n_1204),
.B(n_109),
.C(n_111),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1208),
.B(n_931),
.Y(n_1217)
);

XOR2xp5_ASAP7_75t_L g1218 ( 
.A(n_1203),
.B(n_112),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1198),
.A2(n_930),
.B1(n_994),
.B2(n_931),
.C(n_924),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1195),
.A2(n_930),
.B1(n_912),
.B2(n_931),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1200),
.Y(n_1221)
);

OAI211xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1207),
.A2(n_113),
.B(n_115),
.C(n_117),
.Y(n_1222)
);

XNOR2x1_ASAP7_75t_L g1223 ( 
.A(n_1209),
.B(n_120),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1202),
.A2(n_924),
.B1(n_931),
.B2(n_913),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1218),
.A2(n_930),
.B1(n_913),
.B2(n_917),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1221),
.A2(n_930),
.B1(n_913),
.B2(n_917),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1210),
.Y(n_1227)
);

AOI22x1_ASAP7_75t_L g1228 ( 
.A1(n_1213),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1212),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1215),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1216),
.A2(n_917),
.B1(n_929),
.B2(n_919),
.Y(n_1231)
);

AOI211xp5_ASAP7_75t_L g1232 ( 
.A1(n_1222),
.A2(n_1211),
.B(n_1217),
.C(n_1219),
.Y(n_1232)
);

OA22x2_ASAP7_75t_L g1233 ( 
.A1(n_1214),
.A2(n_929),
.B1(n_916),
.B2(n_922),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1223),
.A2(n_973),
.B1(n_125),
.B2(n_126),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1227),
.B(n_1220),
.Y(n_1235)
);

XNOR2xp5_ASAP7_75t_L g1236 ( 
.A(n_1229),
.B(n_1224),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1228),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1230),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1231),
.B(n_124),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1234),
.B(n_127),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1238),
.Y(n_1241)
);

XNOR2x2_ASAP7_75t_L g1242 ( 
.A(n_1236),
.B(n_1232),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1240),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1237),
.A2(n_1235),
.B1(n_1239),
.B2(n_1225),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1241),
.A2(n_1233),
.B1(n_1226),
.B2(n_135),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1245),
.A2(n_1244),
.B(n_1243),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1246),
.A2(n_1242),
.B(n_916),
.Y(n_1247)
);

XOR2xp5_ASAP7_75t_L g1248 ( 
.A(n_1247),
.B(n_131),
.Y(n_1248)
);

OAI221xp5_ASAP7_75t_R g1249 ( 
.A1(n_1248),
.A2(n_132),
.B1(n_137),
.B2(n_141),
.C(n_147),
.Y(n_1249)
);

AOI211xp5_ASAP7_75t_L g1250 ( 
.A1(n_1249),
.A2(n_149),
.B(n_151),
.C(n_153),
.Y(n_1250)
);


endmodule