module real_jpeg_1666_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_0),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_37),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_2),
.A2(n_26),
.B1(n_74),
.B2(n_77),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_3),
.A2(n_32),
.B1(n_37),
.B2(n_64),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_64),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_3),
.A2(n_64),
.B1(n_74),
.B2(n_77),
.Y(n_179)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_5),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_155),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_5),
.A2(n_32),
.B1(n_37),
.B2(n_155),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_5),
.A2(n_74),
.B1(n_77),
.B2(n_155),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_6),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_6),
.A2(n_32),
.B1(n_37),
.B2(n_88),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_88),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_6),
.A2(n_74),
.B1(n_77),
.B2(n_88),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_7),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_7),
.A2(n_32),
.B1(n_37),
.B2(n_96),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_96),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_7),
.A2(n_74),
.B1(n_77),
.B2(n_96),
.Y(n_200)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_8),
.Y(n_346)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_10),
.A2(n_32),
.B1(n_37),
.B2(n_186),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_186),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_10),
.A2(n_74),
.B1(n_77),
.B2(n_186),
.Y(n_271)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_13),
.B(n_41),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_13),
.B(n_53),
.C(n_55),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_13),
.B(n_52),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_13),
.B(n_71),
.C(n_74),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_221),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_13),
.B(n_123),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_13),
.B(n_78),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_13),
.A2(n_32),
.B1(n_37),
.B2(n_221),
.Y(n_286)
);

BUFx6f_ASAP7_75t_SL g344 ( 
.A(n_14),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_14),
.B(n_346),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_15),
.A2(n_27),
.B1(n_29),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_15),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_15),
.A2(n_32),
.B1(n_37),
.B2(n_133),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_15),
.A2(n_54),
.B1(n_55),
.B2(n_133),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_15),
.A2(n_74),
.B1(n_77),
.B2(n_133),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_16),
.A2(n_27),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_16),
.A2(n_32),
.B1(n_37),
.B2(n_40),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_16),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_16),
.A2(n_40),
.B1(n_74),
.B2(n_77),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_344),
.B(n_345),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_45),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_23),
.B(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_24),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_24),
.B(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_39),
.B2(n_41),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_30),
.B1(n_41),
.B2(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_27),
.A2(n_86),
.B(n_221),
.C(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_27),
.B(n_221),
.Y(n_222)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_27),
.A2(n_34),
.A3(n_37),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_39),
.B(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_30),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_30),
.A2(n_41),
.B1(n_154),
.B2(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_38),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_31),
.A2(n_63),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_31),
.A2(n_86),
.B1(n_87),
.B2(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_31),
.A2(n_95),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_31),
.B(n_132),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_31),
.A2(n_130),
.B(n_307),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_37),
.B1(n_53),
.B2(n_57),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_32),
.B(n_211),
.Y(n_210)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_32),
.B(n_35),
.Y(n_235)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI21x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_339),
.B(n_341),
.Y(n_45)
);

AOI21x1_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_101),
.B(n_338),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_89),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_48),
.B(n_89),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_67),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_59),
.Y(n_50)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_51),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_52),
.B(n_183),
.Y(n_287)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_52)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_55),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_55),
.B(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_61),
.B(n_65),
.C(n_67),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_81),
.C(n_85),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_81),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_94),
.C(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_93),
.B1(n_98),
.B2(n_99),
.Y(n_113)
);

OAI21x1_ASAP7_75t_R g68 ( 
.A1(n_69),
.A2(n_78),
.B(n_79),
.Y(n_68)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_69),
.A2(n_78),
.B1(n_128),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_69),
.A2(n_78),
.B1(n_149),
.B2(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_69),
.A2(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_69),
.B(n_207),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_80),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_73),
.A2(n_109),
.B1(n_110),
.B2(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_73),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_73),
.A2(n_228),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_73),
.A2(n_109),
.B1(n_204),
.B2(n_254),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_74),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_74),
.B(n_267),
.Y(n_266)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_78),
.B(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_84),
.B1(n_100),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_82),
.A2(n_84),
.B1(n_107),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_82),
.A2(n_84),
.B1(n_194),
.B2(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_82),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_82),
.A2(n_225),
.B(n_287),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_84),
.A2(n_151),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_84),
.A2(n_182),
.B(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_86),
.A2(n_153),
.B(n_156),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.C(n_97),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_90),
.A2(n_94),
.B1(n_112),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_97),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_162),
.B(n_335),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_158),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_134),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_104),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_104),
.B(n_134),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_104),
.B(n_159),
.Y(n_337)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_111),
.CI(n_115),
.CON(n_104),
.SN(n_104)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_106),
.B(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_109),
.A2(n_206),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_119),
.B(n_129),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_117),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_126),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_119),
.B1(n_129),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_118),
.A2(n_119),
.B1(n_126),
.B2(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_123),
.B(n_124),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_120),
.A2(n_123),
.B1(n_146),
.B2(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_120),
.A2(n_221),
.B(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_121),
.A2(n_122),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_121),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_121),
.A2(n_122),
.B1(n_201),
.B2(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_121),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_121),
.A2(n_122),
.B1(n_246),
.B2(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_122),
.A2(n_200),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_122),
.B(n_215),
.Y(n_248)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_123),
.A2(n_214),
.B(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.C(n_141),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_150),
.C(n_152),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_143),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_144),
.A2(n_147),
.B1(n_148),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_144),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_150),
.B(n_152),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_157),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_158),
.A2(n_336),
.B(n_337),
.Y(n_335)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_187),
.B(n_334),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_164),
.B(n_167),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.C(n_173),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_168),
.B(n_171),
.Y(n_332)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_173),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_180),
.C(n_184),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_174),
.A2(n_175),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_176),
.B(n_178),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_177),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_184),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_185),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_329),
.B(n_333),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_298),
.B(n_326),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_240),
.B(n_297),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_216),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_191),
.B(n_216),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_202),
.C(n_208),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_192),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_196),
.C(n_199),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_202),
.B(n_208),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_212),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_230),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_217),
.B(n_231),
.C(n_239),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_223),
.B2(n_229),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_218),
.B(n_224),
.C(n_226),
.Y(n_311)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_239),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_232),
.B(n_237),
.Y(n_302)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_292),
.B(n_296),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_281),
.B(n_291),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_263),
.B(n_280),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_257),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_257),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_249),
.B1(n_255),
.B2(n_256),
.Y(n_244)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_252),
.C(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_274),
.B(n_279),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_269),
.B(n_273),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_272),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_277),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_283),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_288),
.C(n_289),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_295),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_313),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_312),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_312),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_309),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_310),
.C(n_311),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_304),
.C(n_308),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_308),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_325),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_325),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_319),
.C(n_321),
.Y(n_330)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_321),
.Y(n_318)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_331),
.Y(n_333)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_340),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);


endmodule