module real_jpeg_5957_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_1),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_1),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_1),
.A2(n_141),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_1),
.A2(n_141),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_1),
.A2(n_141),
.B1(n_362),
.B2(n_365),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_2),
.A2(n_45),
.B1(n_68),
.B2(n_169),
.Y(n_215)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_60),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_4),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_4),
.A2(n_79),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_4),
.A2(n_79),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_5),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_5),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_5),
.A2(n_80),
.B1(n_109),
.B2(n_169),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_5),
.A2(n_109),
.B1(n_142),
.B2(n_225),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_5),
.A2(n_35),
.B1(n_109),
.B2(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_6),
.A2(n_142),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_6),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_6),
.A2(n_188),
.B1(n_298),
.B2(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_6),
.A2(n_188),
.B1(n_260),
.B2(n_338),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_6),
.A2(n_188),
.B1(n_383),
.B2(n_401),
.Y(n_400)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_7),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_8),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_8),
.Y(n_263)
);

INVx8_ASAP7_75t_L g350 ( 
.A(n_8),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_9),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_9),
.A2(n_252),
.B1(n_284),
.B2(n_287),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_9),
.B(n_300),
.C(n_304),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_9),
.B(n_99),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_9),
.B(n_43),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_9),
.B(n_81),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_9),
.B(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_12),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_12),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_12),
.Y(n_140)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_12),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_12),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_12),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_12),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_13),
.A2(n_37),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_14),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_14),
.A2(n_59),
.B1(n_116),
.B2(n_120),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_14),
.A2(n_59),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_15),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_16),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_16),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_16),
.A2(n_148),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_16),
.A2(n_148),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_16),
.A2(n_148),
.B1(n_177),
.B2(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_229),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_228),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_197),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_20),
.B(n_197),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_152),
.C(n_164),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_21),
.B(n_152),
.CI(n_164),
.CON(n_273),
.SN(n_273)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_22),
.B(n_83),
.C(n_121),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_23),
.B(n_51),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_34),
.B1(n_41),
.B2(n_44),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_24),
.A2(n_44),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_24),
.A2(n_255),
.B1(n_261),
.B2(n_264),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_24),
.A2(n_309),
.B(n_314),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_24),
.A2(n_252),
.B(n_314),
.Y(n_334)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_25),
.A2(n_174),
.B1(n_181),
.B2(n_182),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_25),
.B(n_315),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_25),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_25),
.A2(n_256),
.B1(n_375),
.B2(n_407),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_32),
.Y(n_257)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_32),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_34),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_36),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_36),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g377 ( 
.A(n_36),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_40),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_43),
.Y(n_182)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_47),
.Y(n_177)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_47),
.Y(n_306)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_50),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_64),
.B1(n_78),
.B2(n_81),
.Y(n_51)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_52),
.Y(n_172)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_56),
.Y(n_170)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_57),
.Y(n_365)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_58),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_58),
.Y(n_298)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AO22x2_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_100),
.B1(n_103),
.B2(n_104),
.Y(n_99)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_63),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_63),
.Y(n_323)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_63),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_64),
.A2(n_78),
.B1(n_81),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_64),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_64),
.A2(n_81),
.B1(n_155),
.B2(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_64),
.B(n_291),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_70),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_66),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_70),
.A2(n_320),
.B(n_324),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_76),
.Y(n_332)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_81),
.B(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_121),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_105),
.B1(n_114),
.B2(n_115),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_84),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_84),
.A2(n_114),
.B1(n_267),
.B2(n_400),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_99),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_90),
.Y(n_371)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_93),
.Y(n_208)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_94),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_94),
.Y(n_271)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_98),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_99),
.Y(n_114)
);

AOI22x1_ASAP7_75t_L g189 ( 
.A1(n_99),
.A2(n_190),
.B1(n_191),
.B2(n_196),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_99),
.A2(n_190),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g386 ( 
.A(n_101),
.Y(n_386)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_103),
.Y(n_294)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_113),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_114),
.B(n_192),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_114),
.A2(n_400),
.B(n_403),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_119),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_137),
.B(n_146),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_122),
.A2(n_131),
.B1(n_137),
.B2(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_123),
.B(n_147),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_123),
.A2(n_422),
.B(n_423),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_126),
.Y(n_248)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_131),
.B(n_252),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_131)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_132),
.Y(n_250)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_139),
.B(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_140),
.Y(n_247)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_146),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_151),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_151),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_160),
.B2(n_163),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_154),
.B(n_160),
.Y(n_219)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_156),
.Y(n_384)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_157),
.Y(n_292)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_163),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_161),
.A2(n_337),
.B(n_340),
.Y(n_336)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_161),
.Y(n_407)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_183),
.C(n_189),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_165),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_166),
.B(n_173),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_167),
.A2(n_283),
.B(n_290),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_167),
.A2(n_171),
.B1(n_320),
.B2(n_361),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_167),
.A2(n_290),
.B(n_361),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_168),
.A2(n_171),
.B(n_324),
.Y(n_426)
);

INVx5_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_174),
.Y(n_264)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_183),
.A2(n_184),
.B1(n_189),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_185),
.A2(n_227),
.B(n_241),
.Y(n_240)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_189),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_190),
.A2(n_266),
.B(n_272),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_190),
.A2(n_272),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_190),
.B(n_191),
.Y(n_403)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_193),
.B(n_250),
.Y(n_249)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_217),
.B2(n_218),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_212),
.B(n_216),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_213),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_244),
.A3(n_248),
.B1(n_249),
.B2(n_251),
.Y(n_243)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_274),
.B(n_451),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_273),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_232),
.B(n_273),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.C(n_238),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_237),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_238),
.B(n_441),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.C(n_265),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_239),
.A2(n_240),
.B1(n_265),
.B2(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_242),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_253),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_243),
.A2(n_253),
.B1(n_254),
.B2(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_243),
.Y(n_415)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_SL g422 ( 
.A1(n_245),
.A2(n_251),
.B(n_252),
.Y(n_422)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_SL g368 ( 
.A1(n_252),
.A2(n_270),
.B(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_265),
.Y(n_436)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx6_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g453 ( 
.A(n_273),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_429),
.B(n_448),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_410),
.B(n_428),
.Y(n_276)
);

AO21x1_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_391),
.B(n_409),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_355),
.B(n_390),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_327),
.B(n_354),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_307),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_281),
.B(n_307),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_295),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_282),
.A2(n_295),
.B1(n_296),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_282),
.Y(n_352)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_318),
.C(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_309),
.Y(n_346)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_325),
.B2(n_326),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_343),
.B(n_353),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_335),
.B(n_342),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_334),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_341),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_337),
.Y(n_345)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_340),
.A2(n_374),
.B(n_378),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_351),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_351),
.Y(n_353)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx8_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_357),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_372),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_366),
.B2(n_367),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_366),
.C(n_372),
.Y(n_392)
);

INVx3_ASAP7_75t_SL g362 ( 
.A(n_363),
.Y(n_362)
);

INVx8_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AOI32xp33_ASAP7_75t_L g381 ( 
.A1(n_370),
.A2(n_382),
.A3(n_384),
.B1(n_385),
.B2(n_387),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_381),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_381),
.Y(n_397)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx5_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp33_ASAP7_75t_SL g387 ( 
.A(n_386),
.B(n_388),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_392),
.B(n_393),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_395),
.B1(n_398),
.B2(n_408),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_397),
.C(n_408),
.Y(n_411)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_398),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_405),
.C(n_406),
.Y(n_416)
);

INVx8_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_411),
.B(n_412),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_419),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.Y(n_413)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_414),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_416),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_417),
.C(n_419),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_424),
.B2(n_427),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_425),
.C(n_426),
.Y(n_439)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_424),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_443),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_432),
.A2(n_449),
.B(n_450),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_440),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_440),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.C(n_439),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_446),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_437),
.A2(n_438),
.B1(n_439),
.B2(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_439),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_444),
.B(n_445),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);


endmodule