module fake_jpeg_4778_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_21),
.B(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_45),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_36),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_65),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_49),
.B(n_62),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_26),
.B1(n_29),
.B2(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_53),
.B1(n_18),
.B2(n_17),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_16),
.B1(n_30),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_31),
.B1(n_22),
.B2(n_24),
.Y(n_83)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_30),
.B1(n_29),
.B2(n_32),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_30),
.B1(n_20),
.B2(n_33),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_40),
.Y(n_93)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_71),
.Y(n_114)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_78),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_97),
.B1(n_25),
.B2(n_22),
.Y(n_104)
);

NAND2x1_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_39),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_49),
.B(n_54),
.C(n_56),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_81),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_46),
.C(n_41),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_80),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_87),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_94),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_36),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_34),
.Y(n_126)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_98),
.Y(n_105)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_18),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_48),
.A2(n_28),
.B1(n_17),
.B2(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_28),
.B1(n_21),
.B2(n_31),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_27),
.B1(n_24),
.B2(n_33),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_127),
.B(n_123),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_54),
.B(n_49),
.C(n_32),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_77),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_123),
.B1(n_71),
.B2(n_90),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_37),
.A3(n_39),
.B1(n_40),
.B2(n_66),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_124),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_63),
.C(n_61),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_120),
.C(n_76),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_119),
.B1(n_80),
.B2(n_88),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_66),
.B1(n_52),
.B2(n_69),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_61),
.C(n_63),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_126),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_37),
.A3(n_66),
.B1(n_42),
.B2(n_58),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_129),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_130),
.B(n_132),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_123),
.A2(n_87),
.B1(n_82),
.B2(n_73),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_103),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_142),
.B1(n_144),
.B2(n_147),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_156),
.B1(n_113),
.B2(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_139),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_137),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_86),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_99),
.B(n_25),
.Y(n_177)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_91),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_76),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_75),
.B1(n_72),
.B2(n_27),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_112),
.B1(n_32),
.B2(n_70),
.Y(n_184)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g148 ( 
.A(n_125),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_148),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_155),
.A2(n_108),
.B(n_124),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_100),
.A2(n_75),
.B1(n_27),
.B2(n_31),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_116),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_126),
.C(n_121),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_169),
.C(n_173),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_161),
.A2(n_182),
.B1(n_0),
.B2(n_1),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_162),
.A2(n_167),
.B(n_177),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_107),
.B1(n_118),
.B2(n_103),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_164),
.A2(n_13),
.B1(n_12),
.B2(n_2),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_189),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_117),
.B(n_99),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_34),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_183),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_91),
.C(n_58),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_188),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_112),
.B(n_68),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_185),
.B1(n_134),
.B2(n_156),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_131),
.A2(n_70),
.B1(n_68),
.B2(n_34),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_187),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_34),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_34),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_157),
.A2(n_34),
.B(n_91),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_19),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_175),
.B1(n_164),
.B2(n_161),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_133),
.B1(n_153),
.B2(n_152),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_200),
.A2(n_213),
.B1(n_217),
.B2(n_171),
.Y(n_233)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_202),
.B(n_203),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_179),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_135),
.Y(n_204)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_138),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_212),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_144),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_138),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_130),
.B1(n_147),
.B2(n_151),
.Y(n_213)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_168),
.A2(n_150),
.A3(n_138),
.B1(n_146),
.B2(n_137),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_129),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_173),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_174),
.A2(n_68),
.B1(n_19),
.B2(n_2),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_184),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_235),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_SL g269 ( 
.A(n_223),
.B(n_236),
.C(n_1),
.Y(n_269)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_240),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_231),
.B1(n_236),
.B2(n_239),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_169),
.C(n_181),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_229),
.C(n_246),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_174),
.C(n_165),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_168),
.B1(n_171),
.B2(n_182),
.Y(n_231)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_177),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_193),
.B1(n_194),
.B2(n_218),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_200),
.B1(n_178),
.B2(n_215),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_207),
.C(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_237),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_198),
.B1(n_204),
.B2(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_232),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_264),
.B(n_268),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_217),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_255),
.B(n_259),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_197),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_263),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_208),
.B1(n_162),
.B2(n_167),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_191),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_265),
.B(n_266),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_216),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_232),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_0),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_234),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_233),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_246),
.C(n_228),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_229),
.C(n_234),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_222),
.C(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_224),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_257),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_248),
.B(n_251),
.C(n_269),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_283),
.A2(n_13),
.B1(n_12),
.B2(n_7),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_225),
.C(n_244),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_273),
.C(n_282),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_3),
.B(n_5),
.Y(n_286)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_254),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_296),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_257),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_295),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_252),
.C(n_263),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_262),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_272),
.B1(n_271),
.B2(n_280),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_12),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_299),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_11),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_5),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_286),
.Y(n_302)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_278),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_298),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_305),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_283),
.B1(n_275),
.B2(n_284),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_306),
.A2(n_307),
.B(n_294),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_277),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_277),
.B1(n_6),
.B2(n_7),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_311),
.C(n_291),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_5),
.C(n_6),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_6),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_312),
.A2(n_7),
.B(n_8),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_317),
.C(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_322),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_323),
.B1(n_311),
.B2(n_312),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_291),
.C(n_304),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_8),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_325),
.B(n_330),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_327),
.A2(n_319),
.B(n_314),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_304),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_314),
.C(n_323),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_302),
.Y(n_330)
);

AO221x1_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_332),
.B1(n_328),
.B2(n_329),
.C(n_327),
.Y(n_334)
);

OAI321xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_333),
.A3(n_324),
.B1(n_326),
.B2(n_10),
.C(n_11),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_9),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_9),
.B(n_11),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_337),
.Y(n_338)
);


endmodule