module real_jpeg_2668_n_16 (n_5, n_4, n_8, n_0, n_12, n_409, n_410, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_409;
input n_410;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_1),
.B(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_1),
.B(n_39),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_1),
.B(n_53),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_1),
.B(n_105),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_1),
.B(n_146),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_2),
.B(n_32),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_2),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_2),
.B(n_43),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_2),
.B(n_39),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_2),
.B(n_53),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_2),
.B(n_105),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_2),
.B(n_146),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_2),
.B(n_187),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_4),
.B(n_34),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_4),
.B(n_39),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_4),
.B(n_53),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_4),
.B(n_105),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_4),
.B(n_146),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_6),
.Y(n_188)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_7),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_7),
.B(n_146),
.Y(n_145)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_9),
.B(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_9),
.B(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_9),
.B(n_105),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_146),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_9),
.B(n_187),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_10),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_10),
.B(n_53),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_12),
.B(n_32),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_12),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_12),
.B(n_43),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_12),
.B(n_39),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_12),
.B(n_53),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_12),
.B(n_105),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_12),
.B(n_187),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_13),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_14),
.B(n_32),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_14),
.B(n_34),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_14),
.B(n_43),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_14),
.B(n_39),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_14),
.B(n_53),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_14),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_14),
.B(n_146),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_14),
.B(n_187),
.Y(n_374)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_301),
.B(n_403),
.C(n_407),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_396),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_378),
.B(n_395),
.Y(n_19)
);

OAI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_337),
.A3(n_360),
.B1(n_376),
.B2(n_377),
.C(n_409),
.Y(n_20)
);

AOI321xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_261),
.A3(n_326),
.B1(n_331),
.B2(n_336),
.C(n_410),
.Y(n_21)
);

NOR3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_190),
.C(n_257),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_151),
.B(n_189),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_116),
.B(n_150),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_88),
.B(n_115),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_65),
.B(n_87),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_44),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_28),
.B(n_44),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.C(n_42),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_29),
.A2(n_30),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_30),
.A2(n_31),
.B(n_33),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_36),
.A2(n_37),
.B1(n_42),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_38),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_41),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_41),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_41),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_54),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_55),
.C(n_59),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_50),
.C(n_51),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_52),
.B(n_100),
.Y(n_124)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_60),
.A2(n_61),
.B1(n_133),
.B2(n_135),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_60),
.A2(n_61),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_61),
.B(n_62),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_61),
.B(n_133),
.C(n_232),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_61),
.B(n_181),
.C(n_292),
.Y(n_317)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_78),
.B(n_86),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_71),
.B(n_77),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_69),
.B(n_112),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_73),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_73),
.B(n_186),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_112),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_76),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_90),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_102),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_101),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_101),
.C(n_102),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_99),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_98),
.C(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_95),
.B(n_186),
.Y(n_292)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_107),
.C(n_114),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_108),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_108),
.A2(n_113),
.B1(n_280),
.B2(n_285),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_108),
.A2(n_113),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_108),
.B(n_281),
.C(n_284),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_108),
.B(n_128),
.C(n_300),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_113),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_110),
.A2(n_111),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_111),
.B(n_199),
.C(n_201),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_112),
.B(n_186),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_118),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_137),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_138),
.C(n_139),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_129),
.B2(n_130),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_131),
.C(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_127),
.B2(n_128),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_125),
.C(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_126),
.B(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_127),
.A2(n_128),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_127),
.A2(n_128),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_128),
.B(n_174),
.C(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_133),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_134),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_149),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_148),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_148),
.C(n_149),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_145),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_153),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_170),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_168),
.B2(n_169),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_156),
.B(n_169),
.C(n_170),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_166),
.C(n_167),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_162),
.C(n_164),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_159),
.B(n_224),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_174),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_174),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_174),
.A2(n_198),
.B1(n_199),
.B2(n_342),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_174),
.B(n_198),
.C(n_282),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_175),
.B(n_207),
.C(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_177),
.C(n_179),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_184),
.C(n_185),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_181),
.A2(n_182),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g332 ( 
.A1(n_191),
.A2(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_226),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_192),
.B(n_226),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_211),
.C(n_212),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_193),
.B(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_194),
.B(n_196),
.C(n_205),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_204),
.B2(n_205),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_203),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_198),
.A2(n_199),
.B1(n_237),
.B2(n_238),
.Y(n_386)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_199),
.B(n_237),
.C(n_310),
.Y(n_399)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_209),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_212),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_225),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_217),
.C(n_225),
.Y(n_246)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_220),
.A2(n_221),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_220),
.B(n_308),
.C(n_310),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_256),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_245),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_228),
.B(n_245),
.C(n_256),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_235),
.C(n_236),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_232),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_232),
.A2(n_233),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_233),
.B(n_354),
.C(n_356),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_237),
.A2(n_238),
.B1(n_271),
.B2(n_272),
.Y(n_402)
);

NOR3xp33_ASAP7_75t_L g407 ( 
.A(n_237),
.B(n_272),
.C(n_345),
.Y(n_407)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_242),
.C(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_241),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_246),
.B(n_248),
.C(n_249),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_255),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_253),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_258),
.B(n_259),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_294),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_262),
.B(n_294),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_276),
.C(n_293),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_263),
.B(n_276),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_264),
.B(n_268),
.C(n_269),
.Y(n_323)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_275),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_271),
.A2(n_272),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_273),
.C(n_275),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_272),
.B(n_317),
.C(n_320),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_273),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_288),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_286),
.B2(n_287),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_287),
.C(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_281),
.A2(n_282),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_294)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_295),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_311),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_311),
.C(n_325),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_297),
.B(n_303),
.C(n_304),
.Y(n_358)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_309),
.B2(n_310),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_307),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_309),
.A2(n_310),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_322),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_315),
.C(n_316),
.Y(n_359)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_327),
.A2(n_332),
.B(n_335),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_328),
.B(n_329),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_338),
.B(n_339),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_361),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_350),
.CI(n_359),
.CON(n_339),
.SN(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_347),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_348),
.C(n_349),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_345),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_345),
.A2(n_346),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_358),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_353),
.C(n_358),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_356),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_375),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_364),
.C(n_375),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_370),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_367),
.C(n_370),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_369),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_373),
.C(n_374),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_394),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_394),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_382),
.C(n_383),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_387),
.B1(n_392),
.B2(n_393),
.Y(n_383)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_384),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_387),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_388),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_389),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_389),
.B(n_390),
.C(n_392),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_406),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_405),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_400),
.B1(n_403),
.B2(n_404),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_399),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_400),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_402),
.Y(n_401)
);


endmodule