module fake_jpeg_10058_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_28),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_59),
.Y(n_86)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_61),
.Y(n_70)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_76),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_51),
.B1(n_46),
.B2(n_52),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_79),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_46),
.B1(n_50),
.B2(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_75),
.Y(n_97)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_43),
.B1(n_48),
.B2(n_45),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_53),
.B1(n_44),
.B2(n_4),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_2),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_83),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_3),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_98),
.Y(n_109)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NAND2x1_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_3),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_108),
.B(n_87),
.C(n_7),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_47),
.B1(n_25),
.B2(n_26),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_86),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_69),
.B1(n_80),
.B2(n_83),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_96),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_111),
.B1(n_105),
.B2(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_97),
.B1(n_100),
.B2(n_104),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_109),
.B1(n_93),
.B2(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_94),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_93),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_98),
.B1(n_102),
.B2(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_10),
.B(n_11),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

AOI221xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_12),
.B1(n_14),
.B2(n_19),
.C(n_20),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_23),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_67),
.C(n_24),
.Y(n_127)
);


endmodule