module fake_netlist_6_1612_n_2465 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_385, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2465);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_385;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2465;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_798;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_544;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_1815;
wire n_659;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_1655;
wire n_1801;
wire n_835;
wire n_1214;
wire n_928;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1317;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_627;
wire n_1767;
wire n_595;
wire n_1779;
wire n_1465;
wire n_524;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_1932;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_1817;
wire n_926;
wire n_2449;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_2460;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1774;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1048;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_1207;
wire n_811;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_1837;
wire n_831;
wire n_964;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_1459;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_1617;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_1390;
wire n_906;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_1601;
wire n_609;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_1456;
wire n_394;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_1548;
wire n_799;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_786;
wire n_1962;
wire n_1236;
wire n_706;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1741;
wire n_1002;
wire n_1325;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_2062;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1882;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_400;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2284;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_1303;
wire n_761;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1737;
wire n_1464;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_472;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_1973;
wire n_708;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1821;
wire n_1537;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_31),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_133),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_258),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_222),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_137),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_371),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_88),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_317),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_24),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_121),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_234),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_283),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_251),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_261),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_233),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_296),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_144),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_271),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_45),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_57),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_0),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_165),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_235),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_358),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_114),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_231),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_380),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_85),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_121),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_290),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_85),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_74),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_243),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_259),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_140),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_340),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_347),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_207),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_200),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_247),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_309),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_324),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_156),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_146),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_386),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_291),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_24),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_172),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_153),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_343),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_232),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_350),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_17),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_377),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_315),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_263),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_304),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_354),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_328),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_35),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_8),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_116),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_268),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_167),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_357),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_72),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_185),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_65),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_82),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_252),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_42),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_361),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_331),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_299),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_335),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_97),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_130),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_132),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_62),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_65),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_260),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_37),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_61),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_154),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_191),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_32),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_73),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_302),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_228),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_381),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_180),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_70),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_32),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_305),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_366),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_39),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_93),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_168),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_367),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_58),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_38),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_89),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_212),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_190),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_79),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_295),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_237),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_16),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_119),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_9),
.Y(n_502)
);

BUFx5_ASAP7_75t_L g503 ( 
.A(n_140),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_274),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_98),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_348),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_39),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_294),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_155),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_161),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_341),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_30),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_284),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_308),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_147),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_314),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_293),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_113),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_246),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_47),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_334),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_215),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_6),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_170),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_248),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_118),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_135),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_316),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_250),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_79),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_286),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_375),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_300),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_95),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_226),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_197),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_28),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_387),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_31),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_12),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_5),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_269),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_139),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_204),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_142),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_195),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_55),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_182),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_72),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_359),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_43),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_365),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_102),
.Y(n_553)
);

INVxp33_ASAP7_75t_R g554 ( 
.A(n_42),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_187),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_112),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_363),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_106),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_313),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_27),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_14),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_22),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_132),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_141),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_123),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_23),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_28),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_276),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_95),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_319),
.Y(n_570)
);

CKINVDCx14_ASAP7_75t_R g571 ( 
.A(n_362),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_173),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_325),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_76),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_66),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_322),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_383),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_75),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_179),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_41),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_298),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_378),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_229),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_175),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_93),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_171),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_333),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_336),
.Y(n_588)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_289),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_157),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_288),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_46),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_41),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_267),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_385),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_255),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_35),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_162),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_2),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_306),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_312),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_46),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_68),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_55),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_372),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_320),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_224),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_106),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_0),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_379),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_209),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_199),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_210),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_90),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_12),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_113),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_326),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_330),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_227),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_339),
.Y(n_620)
);

CKINVDCx16_ASAP7_75t_R g621 ( 
.A(n_115),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_277),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_279),
.Y(n_623)
);

BUFx5_ASAP7_75t_L g624 ( 
.A(n_3),
.Y(n_624)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_285),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_307),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_166),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_74),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_356),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_376),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_58),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_52),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_8),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_5),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_329),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_270),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_220),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_344),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_280),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_145),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_98),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_117),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_257),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_364),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_287),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_198),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_217),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_25),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_321),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_360),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_40),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_311),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_245),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_254),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_112),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_128),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_338),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_342),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_310),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_384),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_275),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_90),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_49),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_13),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_169),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_240),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_281),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_69),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_99),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_164),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_355),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_137),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_345),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_211),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_67),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_181),
.Y(n_676)
);

BUFx2_ASAP7_75t_SL g677 ( 
.A(n_216),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_111),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_52),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_37),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_105),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_122),
.Y(n_682)
);

INVxp33_ASAP7_75t_L g683 ( 
.A(n_382),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_256),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_108),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_176),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_332),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_221),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_43),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_81),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_318),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_301),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_11),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_273),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_102),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_138),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_323),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_346),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_17),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_303),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_76),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_158),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_105),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_349),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_9),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_292),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_38),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_351),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_337),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_53),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_278),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_370),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_241),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_214),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_129),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_13),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_272),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_373),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_297),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_186),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_49),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_101),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_151),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_282),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_352),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_22),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_414),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_503),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_503),
.Y(n_729)
);

INVxp33_ASAP7_75t_L g730 ( 
.A(n_599),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_611),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_503),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_520),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_393),
.Y(n_734)
);

INVxp33_ASAP7_75t_L g735 ( 
.A(n_389),
.Y(n_735)
);

INVxp33_ASAP7_75t_SL g736 ( 
.A(n_388),
.Y(n_736)
);

INVxp33_ASAP7_75t_L g737 ( 
.A(n_389),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_624),
.Y(n_738)
);

INVxp33_ASAP7_75t_L g739 ( 
.A(n_453),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_396),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_624),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_656),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_624),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_624),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_624),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_624),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_624),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_520),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_540),
.Y(n_749)
);

INVxp33_ASAP7_75t_L g750 ( 
.A(n_453),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_540),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_567),
.Y(n_752)
);

CKINVDCx16_ASAP7_75t_R g753 ( 
.A(n_621),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_567),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_701),
.Y(n_755)
);

INVxp33_ASAP7_75t_SL g756 ( 
.A(n_398),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_391),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_410),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_549),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_549),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_656),
.Y(n_761)
);

BUFx5_ASAP7_75t_L g762 ( 
.A(n_394),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_549),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_701),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_549),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_395),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_672),
.B(n_1),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_404),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_391),
.Y(n_769)
);

INVxp33_ASAP7_75t_SL g770 ( 
.A(n_418),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_397),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_556),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_408),
.Y(n_773)
);

CKINVDCx16_ASAP7_75t_R g774 ( 
.A(n_632),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_409),
.Y(n_775)
);

INVxp33_ASAP7_75t_L g776 ( 
.A(n_556),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_417),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_683),
.B(n_1),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_451),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_458),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_471),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_472),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_474),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_656),
.Y(n_784)
);

INVxp33_ASAP7_75t_L g785 ( 
.A(n_560),
.Y(n_785)
);

INVxp33_ASAP7_75t_L g786 ( 
.A(n_560),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_479),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_484),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_485),
.Y(n_789)
);

INVxp33_ASAP7_75t_SL g790 ( 
.A(n_420),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_488),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_494),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_497),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_672),
.B(n_2),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_501),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_530),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_537),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_541),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_551),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_553),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_561),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_562),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_563),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_569),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_400),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_414),
.Y(n_806)
);

INVxp33_ASAP7_75t_L g807 ( 
.A(n_585),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_575),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_578),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_603),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_614),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_628),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_631),
.Y(n_813)
);

INVxp33_ASAP7_75t_SL g814 ( 
.A(n_421),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_642),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_404),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_648),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_403),
.Y(n_818)
);

INVxp33_ASAP7_75t_L g819 ( 
.A(n_585),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_651),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_438),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_678),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_679),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_411),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_716),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_716),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_407),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_413),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_406),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_438),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_693),
.Y(n_831)
);

INVxp67_ASAP7_75t_SL g832 ( 
.A(n_406),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_696),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_699),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_707),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_710),
.Y(n_836)
);

CKINVDCx16_ASAP7_75t_R g837 ( 
.A(n_498),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_480),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_480),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_552),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_415),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_411),
.Y(n_842)
);

INVxp33_ASAP7_75t_L g843 ( 
.A(n_683),
.Y(n_843)
);

CKINVDCx14_ASAP7_75t_R g844 ( 
.A(n_496),
.Y(n_844)
);

INVxp33_ASAP7_75t_SL g845 ( 
.A(n_425),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_552),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_623),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_623),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_401),
.Y(n_849)
);

INVxp33_ASAP7_75t_SL g850 ( 
.A(n_444),
.Y(n_850)
);

INVxp33_ASAP7_75t_L g851 ( 
.A(n_554),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_441),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_416),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_477),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_402),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_412),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_422),
.Y(n_857)
);

INVxp33_ASAP7_75t_SL g858 ( 
.A(n_452),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_419),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_426),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_427),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_424),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_428),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_429),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_430),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_431),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_432),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_433),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_390),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_434),
.Y(n_870)
);

INVxp33_ASAP7_75t_L g871 ( 
.A(n_423),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_437),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_405),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_439),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_390),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_446),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_477),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_454),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_459),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_465),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_466),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_456),
.Y(n_882)
);

CKINVDCx14_ASAP7_75t_R g883 ( 
.A(n_496),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_482),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_487),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_495),
.Y(n_886)
);

CKINVDCx14_ASAP7_75t_R g887 ( 
.A(n_571),
.Y(n_887)
);

CKINVDCx16_ASAP7_75t_R g888 ( 
.A(n_587),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_519),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_522),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_435),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_506),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_392),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_705),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_506),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_460),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_436),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_529),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_441),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_461),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_531),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_545),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_573),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_577),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_581),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_582),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_468),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_469),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_584),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_475),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_596),
.Y(n_911)
);

INVxp33_ASAP7_75t_L g912 ( 
.A(n_423),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_600),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_601),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_612),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_613),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_618),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_622),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_440),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_478),
.Y(n_920)
);

CKINVDCx16_ASAP7_75t_R g921 ( 
.A(n_589),
.Y(n_921)
);

INVxp33_ASAP7_75t_L g922 ( 
.A(n_483),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_442),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_630),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_636),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_638),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_489),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_640),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_513),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_390),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_645),
.Y(n_931)
);

INVxp33_ASAP7_75t_SL g932 ( 
.A(n_492),
.Y(n_932)
);

INVxp67_ASAP7_75t_SL g933 ( 
.A(n_647),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_493),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_665),
.Y(n_935)
);

INVxp67_ASAP7_75t_SL g936 ( 
.A(n_666),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_443),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_445),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_502),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_674),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_505),
.B(n_3),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_676),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_390),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_513),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_455),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_687),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_688),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_694),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_697),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_709),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_719),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_441),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_723),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_725),
.Y(n_954)
);

BUFx5_ASAP7_75t_L g955 ( 
.A(n_591),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_483),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_586),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_447),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_586),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_590),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_512),
.Y(n_961)
);

INVxp33_ASAP7_75t_SL g962 ( 
.A(n_518),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_590),
.Y(n_963)
);

CKINVDCx14_ASAP7_75t_R g964 ( 
.A(n_571),
.Y(n_964)
);

INVxp33_ASAP7_75t_L g965 ( 
.A(n_627),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_627),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_449),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_717),
.Y(n_968)
);

INVxp33_ASAP7_75t_L g969 ( 
.A(n_717),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_455),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_514),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_523),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_399),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_399),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_450),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_455),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_481),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_481),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_637),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_455),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_463),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_457),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_463),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_538),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_462),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_526),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_637),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_658),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_658),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_538),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_538),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_591),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_538),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_605),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_605),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_605),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_605),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_626),
.Y(n_998)
);

INVxp33_ASAP7_75t_SL g999 ( 
.A(n_527),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_626),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_626),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_626),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_714),
.Y(n_1003)
);

BUFx2_ASAP7_75t_SL g1004 ( 
.A(n_514),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_714),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_875),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_765),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_875),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_875),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_852),
.B(n_448),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_759),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_976),
.Y(n_1012)
);

AOI22x1_ASAP7_75t_SL g1013 ( 
.A1(n_727),
.A2(n_500),
.B1(n_507),
.B2(n_470),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_976),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_968),
.B(n_625),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_759),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_760),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_760),
.Y(n_1018)
);

BUFx12f_ASAP7_75t_L g1019 ( 
.A(n_758),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_757),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_763),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_843),
.A2(n_535),
.B1(n_559),
.B2(n_555),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_763),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_869),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_843),
.B(n_591),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_869),
.Y(n_1026)
);

BUFx12f_ASAP7_75t_L g1027 ( 
.A(n_758),
.Y(n_1027)
);

BUFx8_ASAP7_75t_SL g1028 ( 
.A(n_727),
.Y(n_1028)
);

AOI22x1_ASAP7_75t_SL g1029 ( 
.A1(n_981),
.A2(n_500),
.B1(n_507),
.B2(n_470),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_849),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_930),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_852),
.B(n_546),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_837),
.A2(n_535),
.B1(n_559),
.B2(n_555),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_871),
.B(n_568),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_976),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_894),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_976),
.Y(n_1037)
);

INVx6_ASAP7_75t_L g1038 ( 
.A(n_757),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_R g1039 ( 
.A1(n_981),
.A2(n_539),
.B1(n_543),
.B2(n_534),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_855),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_838),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_856),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_943),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_886),
.B(n_464),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_L g1045 ( 
.A(n_734),
.Y(n_1045)
);

BUFx8_ASAP7_75t_SL g1046 ( 
.A(n_768),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_945),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_772),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_839),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_945),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_772),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_970),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_740),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_1004),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_857),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_920),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_970),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_920),
.Y(n_1058)
);

BUFx8_ASAP7_75t_SL g1059 ( 
.A(n_816),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_931),
.B(n_467),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_824),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_840),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_927),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_933),
.B(n_473),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_805),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_888),
.A2(n_606),
.B1(n_649),
.B2(n_564),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_844),
.B(n_629),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_818),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_980),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_827),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_862),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_825),
.Y(n_1072)
);

CKINVDCx6p67_ASAP7_75t_R g1073 ( 
.A(n_753),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_899),
.B(n_579),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_828),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_863),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_778),
.B(n_574),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_927),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_984),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_936),
.B(n_476),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_984),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_994),
.Y(n_1082)
);

NOR2x1_ASAP7_75t_L g1083 ( 
.A(n_899),
.B(n_677),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_939),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_842),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_864),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_994),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_844),
.B(n_629),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_865),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_825),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_1003),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1003),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_939),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_745),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_867),
.Y(n_1095)
);

BUFx12f_ASAP7_75t_L g1096 ( 
.A(n_841),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_730),
.A2(n_574),
.B1(n_675),
.B2(n_602),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_831),
.Y(n_1098)
);

BUFx8_ASAP7_75t_SL g1099 ( 
.A(n_854),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_730),
.A2(n_602),
.B1(n_685),
.B2(n_675),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_853),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_831),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_990),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_728),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_952),
.B(n_588),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_991),
.Y(n_1106)
);

OA22x2_ASAP7_75t_SL g1107 ( 
.A1(n_731),
.A2(n_689),
.B1(n_721),
.B2(n_685),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_972),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_952),
.B(n_686),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_993),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_995),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_868),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_859),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_883),
.B(n_629),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_846),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_729),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_870),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_972),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_996),
.Y(n_1119)
);

BUFx8_ASAP7_75t_L g1120 ( 
.A(n_955),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_997),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_998),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_733),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_SL g1124 ( 
.A(n_778),
.B(n_689),
.Y(n_1124)
);

BUFx8_ASAP7_75t_SL g1125 ( 
.A(n_877),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_732),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_900),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1000),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1001),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1002),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_860),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1005),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_738),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_741),
.Y(n_1134)
);

BUFx8_ASAP7_75t_SL g1135 ( 
.A(n_892),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_992),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_872),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_861),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_743),
.Y(n_1139)
);

INVx5_ASAP7_75t_L g1140 ( 
.A(n_992),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_874),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_744),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_951),
.B(n_486),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_907),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_876),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_746),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_910),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_878),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_747),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_934),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_866),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_921),
.A2(n_606),
.B1(n_649),
.B2(n_564),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_961),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_956),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_766),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_847),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_771),
.Y(n_1157)
);

AND2x6_ASAP7_75t_L g1158 ( 
.A(n_957),
.B(n_714),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_871),
.A2(n_558),
.B1(n_565),
.B2(n_547),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_773),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_912),
.B(n_490),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_891),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_897),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_794),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_L g1165 ( 
.A(n_959),
.B(n_714),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_919),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_769),
.B(n_491),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_829),
.B(n_499),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_762),
.Y(n_1169)
);

INVx5_ASAP7_75t_L g1170 ( 
.A(n_883),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_762),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_775),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_923),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_937),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_938),
.Y(n_1175)
);

INVx5_ASAP7_75t_L g1176 ( 
.A(n_887),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_912),
.B(n_566),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_762),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_958),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_960),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_963),
.A2(n_508),
.B(n_504),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_832),
.B(n_509),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_826),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1030),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1040),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1036),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1006),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1047),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1006),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1006),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1047),
.Y(n_1191)
);

INVx6_ASAP7_75t_L g1192 ( 
.A(n_1170),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1047),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1042),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1052),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1052),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_1034),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1046),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1134),
.B(n_762),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1055),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1038),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1071),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1134),
.B(n_762),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1076),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1086),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1077),
.A2(n_1124),
.B1(n_1159),
.B2(n_1034),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1089),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1052),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1183),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1008),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1095),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1069),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1069),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1112),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1117),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1137),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1141),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1142),
.B(n_762),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1069),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1022),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1079),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1038),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1020),
.B(n_748),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1145),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1183),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1020),
.B(n_749),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1142),
.B(n_922),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1079),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1148),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1133),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1079),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1133),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1025),
.B(n_896),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1133),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1104),
.B(n_922),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1139),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1008),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1139),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1041),
.B(n_751),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1012),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1012),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1170),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1041),
.B(n_752),
.Y(n_1243)
);

INVxp67_ASAP7_75t_L g1244 ( 
.A(n_1177),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1012),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1087),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1014),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1146),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1149),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1149),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1131),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1177),
.B(n_1123),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1149),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1014),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1116),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1126),
.B(n_965),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1155),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1155),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1094),
.B(n_965),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1087),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1155),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1094),
.A2(n_966),
.B(n_880),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1164),
.B(n_908),
.Y(n_1263)
);

CKINVDCx16_ASAP7_75t_R g1264 ( 
.A(n_1061),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1024),
.B(n_969),
.Y(n_1265)
);

XNOR2x2_ASAP7_75t_R g1266 ( 
.A(n_1033),
.B(n_1066),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1087),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1157),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1164),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1091),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1044),
.A2(n_881),
.B(n_879),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1091),
.Y(n_1272)
);

AND2x6_ASAP7_75t_L g1273 ( 
.A(n_1067),
.B(n_848),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1024),
.B(n_969),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1157),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1014),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1037),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1037),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1157),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1037),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1091),
.Y(n_1281)
);

INVxp67_ASAP7_75t_L g1282 ( 
.A(n_1015),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1160),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1026),
.B(n_955),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1009),
.Y(n_1285)
);

NAND2xp33_ASAP7_75t_L g1286 ( 
.A(n_1015),
.B(n_955),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1160),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1103),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1010),
.B(n_955),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1152),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1160),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1026),
.B(n_955),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1031),
.B(n_955),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1049),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1009),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1035),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1103),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1031),
.B(n_884),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1061),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1010),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1103),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1049),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1062),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1106),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1106),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1050),
.B(n_885),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1050),
.B(n_889),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1106),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1161),
.B(n_806),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1057),
.B(n_890),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1044),
.A2(n_901),
.B(n_898),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1161),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1058),
.B(n_986),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1062),
.Y(n_1314)
);

AND2x6_ASAP7_75t_L g1315 ( 
.A(n_1088),
.B(n_902),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1115),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1115),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1110),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1110),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1110),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1156),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1111),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1032),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1056),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1111),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1084),
.B(n_873),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1111),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1156),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1056),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1077),
.A2(n_657),
.B1(n_721),
.B2(n_882),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1119),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1119),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1032),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1119),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1057),
.B(n_903),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1007),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1083),
.B(n_754),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1092),
.B(n_904),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1201),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1312),
.B(n_1060),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1312),
.B(n_1060),
.Y(n_1341)
);

OA22x2_ASAP7_75t_L g1342 ( 
.A1(n_1206),
.A2(n_1078),
.B1(n_1093),
.B2(n_1063),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1262),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1282),
.B(n_1144),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1206),
.A2(n_1124),
.B1(n_767),
.B2(n_1181),
.Y(n_1345)
);

BUFx10_ASAP7_75t_L g1346 ( 
.A(n_1198),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1184),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_SL g1348 ( 
.A(n_1251),
.B(n_1019),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1282),
.B(n_1144),
.Y(n_1349)
);

NAND2xp33_ASAP7_75t_SL g1350 ( 
.A(n_1300),
.B(n_1054),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1244),
.B(n_1144),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1187),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1262),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1185),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1186),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1296),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1194),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1244),
.B(n_1064),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1323),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1295),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1187),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1333),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1295),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1299),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1200),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1289),
.B(n_1144),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1298),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1202),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1289),
.B(n_1252),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1197),
.B(n_1074),
.Y(n_1370)
);

AND3x1_ASAP7_75t_L g1371 ( 
.A(n_1330),
.B(n_1159),
.C(n_1153),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1281),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1271),
.A2(n_1311),
.B1(n_1197),
.B2(n_1286),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1298),
.Y(n_1374)
);

INVx8_ASAP7_75t_L g1375 ( 
.A(n_1273),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1306),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1306),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1307),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1233),
.B(n_1147),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1204),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1307),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1310),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1192),
.Y(n_1383)
);

AND2x6_ASAP7_75t_L g1384 ( 
.A(n_1326),
.B(n_1114),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1209),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1205),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1223),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1281),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1207),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_SL g1390 ( 
.A(n_1329),
.B(n_1027),
.Y(n_1390)
);

AND2x6_ASAP7_75t_L g1391 ( 
.A(n_1263),
.B(n_1074),
.Y(n_1391)
);

BUFx16f_ASAP7_75t_R g1392 ( 
.A(n_1266),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1211),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1309),
.B(n_1147),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1313),
.B(n_1127),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1259),
.B(n_1064),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1198),
.Y(n_1397)
);

AND2x6_ASAP7_75t_L g1398 ( 
.A(n_1294),
.B(n_1105),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1269),
.B(n_1127),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1222),
.B(n_1136),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1255),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1281),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1336),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1214),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1310),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1335),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1215),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1216),
.Y(n_1408)
);

NAND2xp33_ASAP7_75t_L g1409 ( 
.A(n_1315),
.B(n_1054),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1335),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1271),
.A2(n_1181),
.B1(n_735),
.B2(n_739),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1259),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1338),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1338),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1311),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1227),
.B(n_1080),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1285),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1217),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1223),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1188),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1191),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1224),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1193),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1195),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1196),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1208),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1229),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1239),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1239),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1212),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1213),
.Y(n_1431)
);

NAND2xp33_ASAP7_75t_R g1432 ( 
.A(n_1220),
.B(n_1013),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1243),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1243),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1227),
.B(n_1235),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1219),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1235),
.B(n_1080),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1256),
.B(n_1143),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_R g1439 ( 
.A(n_1264),
.B(n_1131),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1226),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1221),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1226),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1256),
.B(n_1143),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1302),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1303),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1228),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1314),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1286),
.B(n_1167),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1231),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1299),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1316),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1187),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1246),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1317),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1269),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1330),
.A2(n_735),
.B1(n_739),
.B2(n_737),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1265),
.B(n_1167),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1321),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1260),
.Y(n_1459)
);

INVx6_ASAP7_75t_L g1460 ( 
.A(n_1192),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1337),
.B(n_1147),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1267),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1265),
.B(n_1168),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1328),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1290),
.B(n_1045),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1270),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1272),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1284),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1274),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1274),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1209),
.Y(n_1471)
);

AND2x6_ASAP7_75t_L g1472 ( 
.A(n_1337),
.B(n_1105),
.Y(n_1472)
);

AO22x2_ASAP7_75t_L g1473 ( 
.A1(n_1266),
.A2(n_1097),
.B1(n_1100),
.B2(n_1029),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1278),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1292),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1315),
.A2(n_737),
.B1(n_776),
.B2(n_750),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1292),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1293),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1315),
.B(n_1273),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1315),
.B(n_1168),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1293),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1324),
.B(n_1150),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1278),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1280),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1199),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1280),
.Y(n_1486)
);

INVx5_ASAP7_75t_L g1487 ( 
.A(n_1192),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1412),
.B(n_1273),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1358),
.B(n_895),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1360),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1412),
.A2(n_1324),
.B1(n_929),
.B2(n_971),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1352),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1343),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1352),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1419),
.B(n_1257),
.Y(n_1495)
);

NOR2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1340),
.B(n_1073),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1341),
.B(n_944),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1419),
.B(n_1258),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1476),
.B(n_1147),
.Y(n_1499)
);

AO22x2_ASAP7_75t_L g1500 ( 
.A1(n_1473),
.A2(n_1100),
.B1(n_1097),
.B2(n_1107),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1396),
.B(n_1273),
.Y(n_1501)
);

INVx4_ASAP7_75t_L g1502 ( 
.A(n_1352),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1339),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1356),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1370),
.B(n_1225),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1352),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1385),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1395),
.B(n_1138),
.Y(n_1508)
);

AND2x6_ASAP7_75t_L g1509 ( 
.A(n_1415),
.B(n_1109),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1356),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1417),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1395),
.B(n_1225),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1343),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1355),
.Y(n_1514)
);

INVx6_ASAP7_75t_L g1515 ( 
.A(n_1346),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1385),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1361),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1471),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1450),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1353),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1455),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1369),
.A2(n_1315),
.B1(n_1230),
.B2(n_1234),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1363),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1361),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1476),
.B(n_1138),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1439),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1472),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1353),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1456),
.B(n_1329),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_SL g1530 ( 
.A(n_1397),
.B(n_1070),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1339),
.B(n_1261),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1363),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1403),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1361),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1415),
.A2(n_1203),
.B(n_1199),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1421),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1474),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1369),
.A2(n_1232),
.B1(n_1238),
.B2(n_1236),
.Y(n_1538)
);

INVx5_ASAP7_75t_L g1539 ( 
.A(n_1472),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1408),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1437),
.B(n_1162),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1347),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1354),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1438),
.B(n_1162),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1421),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1387),
.B(n_1268),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1357),
.Y(n_1547)
);

AO22x2_ASAP7_75t_L g1548 ( 
.A1(n_1473),
.A2(n_1107),
.B1(n_830),
.B2(n_983),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1423),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1456),
.B(n_1063),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1423),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1359),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1424),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1474),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1345),
.A2(n_1150),
.B1(n_1078),
.B2(n_1118),
.C(n_1108),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1424),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1443),
.B(n_1416),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1425),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1365),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1483),
.Y(n_1560)
);

AO22x2_ASAP7_75t_L g1561 ( 
.A1(n_1473),
.A2(n_821),
.B1(n_1039),
.B2(n_941),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1454),
.B(n_1275),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1364),
.Y(n_1563)
);

CKINVDCx16_ASAP7_75t_R g1564 ( 
.A(n_1439),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1482),
.B(n_1399),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1482),
.B(n_1093),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1362),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1361),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1435),
.B(n_1182),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1368),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1400),
.B(n_1305),
.Y(n_1571)
);

NAND2x1p5_ASAP7_75t_L g1572 ( 
.A(n_1400),
.B(n_1305),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1346),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1452),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1469),
.B(n_1182),
.Y(n_1575)
);

AND2x6_ASAP7_75t_L g1576 ( 
.A(n_1479),
.B(n_1109),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1454),
.B(n_1279),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1380),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1483),
.Y(n_1579)
);

INVxp33_ASAP7_75t_L g1580 ( 
.A(n_1399),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1386),
.Y(n_1581)
);

NAND2x1_ASAP7_75t_L g1582 ( 
.A(n_1452),
.B(n_1297),
.Y(n_1582)
);

AND2x6_ASAP7_75t_L g1583 ( 
.A(n_1478),
.B(n_1218),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1470),
.B(n_1108),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1452),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1430),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1367),
.B(n_1053),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1367),
.B(n_1053),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1374),
.B(n_1163),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1457),
.B(n_1118),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1463),
.B(n_1065),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1389),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1431),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1393),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1342),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1374),
.B(n_1376),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1491),
.B(n_1068),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1557),
.B(n_1376),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1514),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1536),
.Y(n_1600)
);

O2A1O1Ixp5_ASAP7_75t_L g1601 ( 
.A1(n_1499),
.A2(n_1448),
.B(n_1366),
.C(n_1351),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1536),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1541),
.B(n_1544),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1565),
.B(n_1377),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1569),
.B(n_1377),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1590),
.B(n_1378),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1580),
.B(n_1101),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1497),
.B(n_1151),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1545),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1545),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1549),
.Y(n_1611)
);

AO22x1_ASAP7_75t_L g1612 ( 
.A1(n_1508),
.A2(n_1472),
.B1(n_1391),
.B2(n_851),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1591),
.B(n_1378),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1549),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1500),
.A2(n_1345),
.B1(n_1382),
.B2(n_1381),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1587),
.B(n_1371),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1566),
.B(n_1342),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1500),
.A2(n_1550),
.B1(n_1561),
.B2(n_1548),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1588),
.B(n_1381),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1489),
.B(n_1173),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1589),
.B(n_1382),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1531),
.B(n_1428),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1512),
.B(n_1175),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1561),
.A2(n_1405),
.B1(n_1410),
.B2(n_1406),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1531),
.B(n_1503),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1555),
.B(n_1163),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1525),
.A2(n_1394),
.B(n_1351),
.C(n_1349),
.Y(n_1627)
);

NAND2xp33_ASAP7_75t_L g1628 ( 
.A(n_1509),
.B(n_1384),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1501),
.A2(n_1373),
.B1(n_1406),
.B2(n_1405),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1551),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1575),
.B(n_1410),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1584),
.B(n_1413),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1596),
.B(n_1413),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1529),
.B(n_1414),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1551),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1553),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1539),
.B(n_1414),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1505),
.B(n_1344),
.Y(n_1638)
);

AOI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1548),
.A2(n_893),
.B1(n_770),
.B2(n_790),
.C(n_756),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1542),
.B(n_1391),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1595),
.A2(n_1485),
.B1(n_1475),
.B2(n_1477),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1543),
.B(n_1391),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1547),
.B(n_1391),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1553),
.Y(n_1644)
);

OAI21xp33_ASAP7_75t_L g1645 ( 
.A1(n_1518),
.A2(n_851),
.B(n_814),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1559),
.B(n_1391),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1556),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1556),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1507),
.B(n_1344),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1492),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1558),
.Y(n_1651)
);

OR2x6_ASAP7_75t_L g1652 ( 
.A(n_1515),
.B(n_1465),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1558),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1515),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1509),
.A2(n_1485),
.B1(n_1481),
.B2(n_1477),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1570),
.B(n_1472),
.Y(n_1656)
);

INVx8_ASAP7_75t_L g1657 ( 
.A(n_1492),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1578),
.B(n_1472),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1516),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1488),
.A2(n_1373),
.B(n_1468),
.Y(n_1660)
);

O2A1O1Ixp5_ASAP7_75t_L g1661 ( 
.A1(n_1582),
.A2(n_1366),
.B(n_1349),
.C(n_1379),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1581),
.B(n_1384),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1592),
.B(n_1384),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1594),
.B(n_1384),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1608),
.A2(n_1521),
.B1(n_1350),
.B2(n_1432),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1603),
.B(n_1085),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1602),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1611),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1599),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1626),
.A2(n_1384),
.B1(n_1509),
.B2(n_1398),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1654),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1654),
.Y(n_1672)
);

OR2x6_ASAP7_75t_L g1673 ( 
.A(n_1657),
.B(n_1465),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1657),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1659),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1626),
.A2(n_1509),
.B1(n_1398),
.B2(n_1433),
.Y(n_1676)
);

NOR2xp67_ASAP7_75t_L g1677 ( 
.A(n_1607),
.B(n_1552),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1608),
.B(n_1085),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1620),
.A2(n_1432),
.B1(n_1530),
.B2(n_1563),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1634),
.B(n_1468),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1625),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1620),
.A2(n_1398),
.B1(n_1434),
.B2(n_1429),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1632),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1644),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1623),
.B(n_1028),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1600),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1647),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1657),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1623),
.B(n_1028),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1609),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1625),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1622),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1622),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1610),
.Y(n_1694)
);

INVx5_ASAP7_75t_L g1695 ( 
.A(n_1652),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1617),
.B(n_1495),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1607),
.B(n_1046),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1634),
.B(n_1475),
.Y(n_1698)
);

AND2x6_ASAP7_75t_L g1699 ( 
.A(n_1651),
.B(n_1493),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1652),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1614),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1653),
.Y(n_1702)
);

INVx4_ASAP7_75t_L g1703 ( 
.A(n_1652),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1604),
.B(n_1481),
.Y(n_1704)
);

OR2x4_ASAP7_75t_L g1705 ( 
.A(n_1597),
.B(n_1392),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1630),
.Y(n_1706)
);

NAND2x1p5_ASAP7_75t_L g1707 ( 
.A(n_1637),
.B(n_1539),
.Y(n_1707)
);

NOR2xp67_ASAP7_75t_L g1708 ( 
.A(n_1649),
.B(n_1075),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1613),
.B(n_1616),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1635),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1683),
.B(n_1606),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1671),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1683),
.A2(n_1618),
.B1(n_1615),
.B2(n_1624),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1677),
.B(n_1638),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1686),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1678),
.A2(n_1624),
.B1(n_1618),
.B2(n_1615),
.Y(n_1716)
);

BUFx8_ASAP7_75t_L g1717 ( 
.A(n_1671),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1674),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1680),
.A2(n_1598),
.B(n_1628),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1669),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1680),
.A2(n_1598),
.B(n_1605),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1666),
.B(n_1059),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1685),
.A2(n_1645),
.B1(n_1564),
.B2(n_1390),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1709),
.B(n_1059),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1671),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1698),
.A2(n_1641),
.B1(n_1655),
.B2(n_1638),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1689),
.B(n_1099),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1679),
.B(n_1708),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1697),
.B(n_1099),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1696),
.B(n_1631),
.Y(n_1730)
);

NOR2xp67_ASAP7_75t_L g1731 ( 
.A(n_1669),
.B(n_1526),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1665),
.A2(n_1696),
.B1(n_1113),
.B2(n_1166),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1693),
.B(n_1649),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1698),
.A2(n_1660),
.B(n_1621),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1695),
.B(n_1639),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1705),
.A2(n_1174),
.B1(n_1179),
.B2(n_1096),
.Y(n_1736)
);

NOR2x1_ASAP7_75t_R g1737 ( 
.A(n_1695),
.B(n_1519),
.Y(n_1737)
);

NOR2xp67_ASAP7_75t_L g1738 ( 
.A(n_1692),
.B(n_1573),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1704),
.A2(n_1619),
.B(n_1629),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1674),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1706),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1690),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1690),
.B(n_1701),
.Y(n_1743)
);

A2O1A1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1676),
.A2(n_1627),
.B(n_1601),
.C(n_1661),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1674),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1672),
.Y(n_1746)
);

A2O1A1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1682),
.A2(n_1394),
.B(n_1379),
.C(n_1662),
.Y(n_1747)
);

AND3x2_ASAP7_75t_L g1748 ( 
.A(n_1700),
.B(n_1348),
.C(n_761),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1701),
.Y(n_1749)
);

A2O1A1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1670),
.A2(n_1664),
.B(n_1663),
.C(n_1658),
.Y(n_1750)
);

O2A1O1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1675),
.A2(n_1461),
.B(n_1465),
.C(n_1637),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1704),
.A2(n_1655),
.B(n_1522),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1688),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1672),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1672),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1692),
.B(n_1567),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1712),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1743),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1742),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1716),
.A2(n_1695),
.B1(n_1641),
.B2(n_1705),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1754),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1755),
.B(n_1695),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1711),
.B(n_1667),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1735),
.A2(n_657),
.B1(n_1612),
.B2(n_1703),
.Y(n_1764)
);

BUFx8_ASAP7_75t_SL g1765 ( 
.A(n_1725),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1749),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1715),
.Y(n_1767)
);

AND2x6_ASAP7_75t_L g1768 ( 
.A(n_1730),
.B(n_1668),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1746),
.B(n_1703),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1712),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1713),
.B(n_1684),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1728),
.B(n_1710),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1741),
.Y(n_1773)
);

INVx4_ASAP7_75t_L g1774 ( 
.A(n_1712),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_R g1775 ( 
.A(n_1717),
.B(n_1688),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1713),
.B(n_1687),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1751),
.B(n_974),
.C(n_973),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1718),
.Y(n_1778)
);

CKINVDCx8_ASAP7_75t_R g1779 ( 
.A(n_1724),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1720),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1745),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1733),
.Y(n_1782)
);

OR2x2_ASAP7_75t_SL g1783 ( 
.A(n_1756),
.B(n_774),
.Y(n_1783)
);

BUFx10_ASAP7_75t_L g1784 ( 
.A(n_1748),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1718),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1740),
.B(n_1681),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1714),
.Y(n_1787)
);

BUFx2_ASAP7_75t_L g1788 ( 
.A(n_1737),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1753),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1717),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1732),
.B(n_1694),
.Y(n_1791)
);

INVxp67_ASAP7_75t_SL g1792 ( 
.A(n_1719),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1722),
.A2(n_1576),
.B1(n_1723),
.B2(n_1398),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1753),
.B(n_1691),
.Y(n_1794)
);

OAI222xp33_ASAP7_75t_L g1795 ( 
.A1(n_1726),
.A2(n_1673),
.B1(n_680),
.B2(n_634),
.C1(n_663),
.C2(n_609),
.Y(n_1795)
);

HAxp5_ASAP7_75t_L g1796 ( 
.A(n_1736),
.B(n_1496),
.CON(n_1796),
.SN(n_1796)
);

INVx4_ASAP7_75t_L g1797 ( 
.A(n_1738),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1726),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1721),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1727),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1734),
.B(n_1702),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1744),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1729),
.A2(n_1576),
.B1(n_1398),
.B2(n_724),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1752),
.Y(n_1804)
);

AOI21xp33_ASAP7_75t_L g1805 ( 
.A1(n_1752),
.A2(n_1642),
.B(n_1640),
.Y(n_1805)
);

BUFx2_ASAP7_75t_R g1806 ( 
.A(n_1731),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1739),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1747),
.A2(n_1409),
.B(n_1646),
.C(n_1643),
.Y(n_1808)
);

OAI21x1_ASAP7_75t_L g1809 ( 
.A1(n_1799),
.A2(n_1707),
.B(n_1656),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1765),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1795),
.A2(n_1750),
.B(n_1576),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_SL g1812 ( 
.A1(n_1760),
.A2(n_1576),
.B1(n_724),
.B2(n_1673),
.Y(n_1812)
);

AO31x2_ASAP7_75t_L g1813 ( 
.A1(n_1807),
.A2(n_1527),
.A3(n_1648),
.B(n_1636),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1759),
.Y(n_1814)
);

OAI21x1_ASAP7_75t_L g1815 ( 
.A1(n_1801),
.A2(n_1707),
.B(n_1535),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1758),
.B(n_1673),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1764),
.A2(n_1498),
.B1(n_1495),
.B2(n_779),
.Y(n_1817)
);

INVx4_ASAP7_75t_L g1818 ( 
.A(n_1757),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1792),
.A2(n_1538),
.B(n_1694),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1802),
.A2(n_1539),
.B(n_1375),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1766),
.Y(n_1821)
);

A2O1A1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1764),
.A2(n_978),
.B(n_979),
.C(n_977),
.Y(n_1822)
);

BUFx8_ASAP7_75t_L g1823 ( 
.A(n_1788),
.Y(n_1823)
);

AO31x2_ASAP7_75t_L g1824 ( 
.A1(n_1808),
.A2(n_1502),
.A3(n_1513),
.B(n_1493),
.Y(n_1824)
);

INVx4_ASAP7_75t_L g1825 ( 
.A(n_1757),
.Y(n_1825)
);

OAI21x1_ASAP7_75t_L g1826 ( 
.A1(n_1771),
.A2(n_1633),
.B(n_1490),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1767),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1782),
.B(n_1710),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1760),
.A2(n_1498),
.B1(n_780),
.B2(n_781),
.Y(n_1829)
);

CKINVDCx14_ASAP7_75t_R g1830 ( 
.A(n_1775),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1787),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1777),
.A2(n_1461),
.B(n_845),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1777),
.A2(n_850),
.B(n_736),
.Y(n_1833)
);

OAI21x1_ASAP7_75t_SL g1834 ( 
.A1(n_1771),
.A2(n_1480),
.B(n_1533),
.Y(n_1834)
);

A2O1A1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1793),
.A2(n_988),
.B(n_989),
.C(n_987),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1791),
.B(n_1710),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1804),
.A2(n_1375),
.B(n_1411),
.Y(n_1837)
);

A2O1A1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1803),
.A2(n_784),
.B(n_742),
.C(n_776),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_SL g1839 ( 
.A1(n_1776),
.A2(n_1540),
.B(n_1401),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1773),
.Y(n_1840)
);

A2O1A1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1798),
.A2(n_785),
.B(n_786),
.C(n_750),
.Y(n_1841)
);

O2A1O1Ixp33_ASAP7_75t_SL g1842 ( 
.A1(n_1772),
.A2(n_809),
.B(n_826),
.C(n_858),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1763),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1763),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1805),
.A2(n_1375),
.B(n_1411),
.Y(n_1845)
);

CKINVDCx14_ASAP7_75t_R g1846 ( 
.A(n_1790),
.Y(n_1846)
);

AO21x1_ASAP7_75t_L g1847 ( 
.A1(n_1776),
.A2(n_782),
.B(n_777),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1783),
.A2(n_1650),
.B1(n_1577),
.B2(n_1562),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1800),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1768),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1768),
.A2(n_724),
.B1(n_1135),
.B2(n_1125),
.Y(n_1851)
);

BUFx3_ASAP7_75t_L g1852 ( 
.A(n_1761),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1768),
.A2(n_1800),
.B1(n_1784),
.B2(n_1797),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1780),
.B(n_1688),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1768),
.A2(n_1135),
.B1(n_1125),
.B2(n_787),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1779),
.B(n_967),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1770),
.Y(n_1857)
);

NOR2xp67_ASAP7_75t_SL g1858 ( 
.A(n_1800),
.B(n_1136),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1805),
.A2(n_1528),
.B(n_1520),
.Y(n_1859)
);

O2A1O1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1796),
.A2(n_788),
.B(n_789),
.C(n_783),
.Y(n_1860)
);

INVx3_ASAP7_75t_L g1861 ( 
.A(n_1774),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1770),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1757),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1778),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_1778),
.Y(n_1865)
);

O2A1O1Ixp33_ASAP7_75t_SL g1866 ( 
.A1(n_1806),
.A2(n_962),
.B(n_999),
.C(n_932),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1778),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1785),
.Y(n_1868)
);

O2A1O1Ixp33_ASAP7_75t_SL g1869 ( 
.A1(n_1784),
.A2(n_786),
.B(n_807),
.C(n_785),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1762),
.A2(n_1528),
.B(n_1494),
.Y(n_1870)
);

OA21x2_ASAP7_75t_L g1871 ( 
.A1(n_1769),
.A2(n_792),
.B(n_791),
.Y(n_1871)
);

NAND2x1p5_ASAP7_75t_L g1872 ( 
.A(n_1762),
.B(n_1492),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1785),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1769),
.A2(n_1506),
.B(n_1494),
.Y(n_1874)
);

O2A1O1Ixp33_ASAP7_75t_SL g1875 ( 
.A1(n_1781),
.A2(n_819),
.B(n_807),
.C(n_795),
.Y(n_1875)
);

O2A1O1Ixp33_ASAP7_75t_L g1876 ( 
.A1(n_1794),
.A2(n_796),
.B(n_797),
.C(n_793),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1785),
.Y(n_1877)
);

O2A1O1Ixp33_ASAP7_75t_SL g1878 ( 
.A1(n_1789),
.A2(n_819),
.B(n_799),
.C(n_800),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1814),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1812),
.A2(n_1794),
.B1(n_1786),
.B2(n_801),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1821),
.Y(n_1881)
);

CKINVDCx9p33_ASAP7_75t_R g1882 ( 
.A(n_1830),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1849),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1817),
.A2(n_1786),
.B1(n_592),
.B2(n_593),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1829),
.A2(n_1789),
.B1(n_1699),
.B2(n_802),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1811),
.A2(n_597),
.B1(n_604),
.B2(n_580),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1831),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1840),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1843),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1833),
.A2(n_615),
.B1(n_616),
.B2(n_608),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1852),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1844),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1836),
.B(n_1789),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1848),
.A2(n_641),
.B1(n_655),
.B2(n_633),
.Y(n_1894)
);

OAI21x1_ASAP7_75t_SL g1895 ( 
.A1(n_1847),
.A2(n_764),
.B(n_755),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1856),
.B(n_975),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1827),
.Y(n_1897)
);

AOI221xp5_ASAP7_75t_L g1898 ( 
.A1(n_1869),
.A2(n_668),
.B1(n_669),
.B2(n_664),
.C(n_662),
.Y(n_1898)
);

OAI21x1_ASAP7_75t_L g1899 ( 
.A1(n_1834),
.A2(n_1593),
.B(n_1586),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1810),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1816),
.B(n_798),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1851),
.A2(n_804),
.B1(n_808),
.B2(n_803),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1850),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1865),
.Y(n_1904)
);

INVx2_ASAP7_75t_SL g1905 ( 
.A(n_1865),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1832),
.A2(n_1855),
.B1(n_1823),
.B2(n_1828),
.Y(n_1906)
);

AOI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1842),
.A2(n_690),
.B1(n_695),
.B2(n_682),
.C(n_681),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1841),
.A2(n_1853),
.B1(n_1846),
.B2(n_1838),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1862),
.Y(n_1909)
);

NAND3xp33_ASAP7_75t_L g1910 ( 
.A(n_1822),
.B(n_811),
.C(n_810),
.Y(n_1910)
);

NAND2x1p5_ASAP7_75t_L g1911 ( 
.A(n_1871),
.B(n_1494),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1813),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1865),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1813),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1857),
.Y(n_1915)
);

OAI222xp33_ASAP7_75t_L g1916 ( 
.A1(n_1858),
.A2(n_726),
.B1(n_715),
.B2(n_722),
.C1(n_703),
.C2(n_1444),
.Y(n_1916)
);

BUFx2_ASAP7_75t_L g1917 ( 
.A(n_1863),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1854),
.B(n_982),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1813),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1864),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1826),
.Y(n_1921)
);

INVx4_ASAP7_75t_L g1922 ( 
.A(n_1868),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1823),
.A2(n_813),
.B1(n_815),
.B2(n_812),
.Y(n_1923)
);

INVx4_ASAP7_75t_L g1924 ( 
.A(n_1868),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1868),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1867),
.B(n_1824),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1877),
.B(n_1154),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_1818),
.Y(n_1928)
);

BUFx2_ASAP7_75t_R g1929 ( 
.A(n_1861),
.Y(n_1929)
);

INVx6_ASAP7_75t_SL g1930 ( 
.A(n_1854),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1926),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1881),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1917),
.B(n_1824),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1887),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1879),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1908),
.B(n_1873),
.Y(n_1936)
);

OAI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1886),
.A2(n_1871),
.B1(n_1835),
.B2(n_1837),
.Y(n_1937)
);

AO21x2_ASAP7_75t_L g1938 ( 
.A1(n_1912),
.A2(n_1839),
.B(n_1820),
.Y(n_1938)
);

AO21x2_ASAP7_75t_L g1939 ( 
.A1(n_1914),
.A2(n_1859),
.B(n_1815),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1888),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1921),
.Y(n_1941)
);

INVx2_ASAP7_75t_SL g1942 ( 
.A(n_1903),
.Y(n_1942)
);

OAI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1908),
.A2(n_1886),
.B(n_1907),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_L g1944 ( 
.A1(n_1919),
.A2(n_1809),
.B(n_1819),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1928),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1915),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1897),
.Y(n_1947)
);

OAI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1885),
.A2(n_1825),
.B1(n_1818),
.B2(n_1870),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1920),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1889),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1909),
.B(n_1928),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1892),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1904),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1909),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1911),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1901),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1911),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1891),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1891),
.B(n_1824),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1899),
.Y(n_1960)
);

OAI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1943),
.A2(n_1929),
.B1(n_1906),
.B2(n_1894),
.Y(n_1961)
);

AOI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1943),
.A2(n_1898),
.B1(n_1907),
.B2(n_1894),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1936),
.A2(n_1884),
.B1(n_1898),
.B2(n_1918),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1937),
.A2(n_1890),
.B1(n_1895),
.B2(n_1906),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_SL g1965 ( 
.A1(n_1937),
.A2(n_1884),
.B1(n_1883),
.B2(n_1896),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1952),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1953),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1951),
.B(n_1893),
.Y(n_1968)
);

AOI222xp33_ASAP7_75t_L g1969 ( 
.A1(n_1956),
.A2(n_1890),
.B1(n_1916),
.B2(n_1923),
.C1(n_1902),
.C2(n_1910),
.Y(n_1969)
);

AND2x4_ASAP7_75t_SL g1970 ( 
.A(n_1956),
.B(n_1883),
.Y(n_1970)
);

BUFx4f_ASAP7_75t_SL g1971 ( 
.A(n_1953),
.Y(n_1971)
);

OAI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1948),
.A2(n_1930),
.B1(n_1924),
.B2(n_1922),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1934),
.A2(n_1880),
.B1(n_1930),
.B2(n_1923),
.Y(n_1973)
);

AOI221xp5_ASAP7_75t_L g1974 ( 
.A1(n_1932),
.A2(n_1916),
.B1(n_1860),
.B2(n_1866),
.C(n_1875),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1952),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1941),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1932),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1951),
.B(n_1925),
.Y(n_1978)
);

AOI221xp5_ASAP7_75t_L g1979 ( 
.A1(n_1931),
.A2(n_909),
.B1(n_911),
.B2(n_906),
.C(n_905),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1958),
.A2(n_1929),
.B1(n_1922),
.B2(n_1924),
.Y(n_1980)
);

BUFx4f_ASAP7_75t_SL g1981 ( 
.A(n_1953),
.Y(n_1981)
);

OAI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1953),
.A2(n_1904),
.B1(n_1913),
.B2(n_1905),
.Y(n_1982)
);

OAI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1959),
.A2(n_1957),
.B(n_1955),
.Y(n_1983)
);

BUFx12f_ASAP7_75t_L g1984 ( 
.A(n_1953),
.Y(n_1984)
);

O2A1O1Ixp5_ASAP7_75t_L g1985 ( 
.A1(n_1955),
.A2(n_1927),
.B(n_1825),
.C(n_1845),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1968),
.B(n_1951),
.Y(n_1986)
);

INVx3_ASAP7_75t_L g1987 ( 
.A(n_1967),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1977),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1975),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1984),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1978),
.B(n_1951),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1976),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1976),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1983),
.B(n_1945),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1965),
.B(n_1949),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1966),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1967),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1967),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1967),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1971),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1970),
.B(n_1945),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1985),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1981),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1982),
.B(n_1947),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1963),
.B(n_1900),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1985),
.Y(n_2006)
);

INVx3_ASAP7_75t_L g2007 ( 
.A(n_1972),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1979),
.Y(n_2008)
);

AOI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1965),
.A2(n_1938),
.B1(n_1960),
.B2(n_1958),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1980),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1961),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1962),
.B(n_817),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1973),
.B(n_1945),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1974),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1964),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1969),
.Y(n_2016)
);

AO21x2_ASAP7_75t_L g2017 ( 
.A1(n_1983),
.A2(n_1941),
.B(n_1944),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1988),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1991),
.B(n_1954),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1991),
.B(n_1954),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_2011),
.A2(n_1957),
.B1(n_1955),
.B2(n_1942),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1987),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1988),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1987),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1989),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_2016),
.A2(n_823),
.B1(n_833),
.B2(n_822),
.C(n_820),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_2016),
.A2(n_2011),
.B1(n_2014),
.B2(n_2015),
.Y(n_2027)
);

OR2x6_ASAP7_75t_L g2028 ( 
.A(n_1990),
.B(n_1882),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1989),
.Y(n_2029)
);

AOI33xp33_ASAP7_75t_L g2030 ( 
.A1(n_2016),
.A2(n_1931),
.A3(n_1947),
.B1(n_1941),
.B2(n_1942),
.B3(n_1933),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_1990),
.Y(n_2031)
);

AOI221xp5_ASAP7_75t_L g2032 ( 
.A1(n_2014),
.A2(n_2012),
.B1(n_2015),
.B2(n_2008),
.C(n_2009),
.Y(n_2032)
);

OAI211xp5_ASAP7_75t_L g2033 ( 
.A1(n_2014),
.A2(n_1878),
.B(n_1876),
.C(n_1933),
.Y(n_2033)
);

OAI33xp33_ASAP7_75t_L g2034 ( 
.A1(n_1996),
.A2(n_1931),
.A3(n_1940),
.B1(n_835),
.B2(n_836),
.B3(n_834),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1992),
.Y(n_2035)
);

INVx1_ASAP7_75t_SL g2036 ( 
.A(n_1990),
.Y(n_2036)
);

OAI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1995),
.A2(n_1953),
.B1(n_1957),
.B2(n_1942),
.Y(n_2037)
);

OAI221xp5_ASAP7_75t_SL g2038 ( 
.A1(n_2008),
.A2(n_1882),
.B1(n_1959),
.B2(n_1960),
.C(n_915),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_2010),
.B(n_2004),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2028),
.B(n_2007),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2028),
.B(n_2007),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2028),
.B(n_2007),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2018),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_2032),
.B(n_2007),
.Y(n_2044)
);

NAND2xp33_ASAP7_75t_L g2045 ( 
.A(n_2027),
.B(n_2010),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2036),
.B(n_2013),
.Y(n_2046)
);

BUFx3_ASAP7_75t_L g2047 ( 
.A(n_2031),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2019),
.B(n_1986),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2023),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2020),
.B(n_1986),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2032),
.B(n_2039),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2022),
.B(n_1997),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_2024),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2035),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_2025),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_2047),
.Y(n_2056)
);

OAI221xp5_ASAP7_75t_L g2057 ( 
.A1(n_2044),
.A2(n_2033),
.B1(n_2038),
.B2(n_2005),
.C(n_2026),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_2047),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_2040),
.B(n_2029),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2055),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_2040),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2041),
.B(n_2013),
.Y(n_2062)
);

BUFx2_ASAP7_75t_L g2063 ( 
.A(n_2041),
.Y(n_2063)
);

OAI221xp5_ASAP7_75t_L g2064 ( 
.A1(n_2051),
.A2(n_2033),
.B1(n_2038),
.B2(n_2026),
.C(n_2002),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2058),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_2063),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2062),
.B(n_2042),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2058),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2061),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2056),
.B(n_2046),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2060),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2065),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_2068),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2066),
.B(n_2045),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2067),
.B(n_2042),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2067),
.B(n_2059),
.Y(n_2076)
);

INVx2_ASAP7_75t_SL g2077 ( 
.A(n_2076),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2074),
.B(n_2070),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_2074),
.B(n_2069),
.Y(n_2079)
);

AOI21xp5_ASAP7_75t_L g2080 ( 
.A1(n_2077),
.A2(n_2045),
.B(n_2057),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2078),
.Y(n_2081)
);

AOI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2081),
.A2(n_2057),
.B1(n_2075),
.B2(n_2064),
.Y(n_2082)
);

O2A1O1Ixp33_ASAP7_75t_L g2083 ( 
.A1(n_2080),
.A2(n_2073),
.B(n_2064),
.C(n_2072),
.Y(n_2083)
);

AOI21xp33_ASAP7_75t_L g2084 ( 
.A1(n_2083),
.A2(n_2079),
.B(n_2069),
.Y(n_2084)
);

XNOR2x1_ASAP7_75t_L g2085 ( 
.A(n_2082),
.B(n_2071),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2084),
.B(n_2059),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2085),
.B(n_2054),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2085),
.Y(n_2088)
);

OAI21xp5_ASAP7_75t_SL g2089 ( 
.A1(n_2086),
.A2(n_2049),
.B(n_2043),
.Y(n_2089)
);

NOR3xp33_ASAP7_75t_L g2090 ( 
.A(n_2088),
.B(n_2055),
.C(n_2053),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2087),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2086),
.Y(n_2092)
);

AOI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_2092),
.A2(n_2053),
.B(n_2052),
.Y(n_2093)
);

OAI21xp33_ASAP7_75t_L g2094 ( 
.A1(n_2090),
.A2(n_2052),
.B(n_2030),
.Y(n_2094)
);

NOR3xp33_ASAP7_75t_L g2095 ( 
.A(n_2091),
.B(n_964),
.C(n_887),
.Y(n_2095)
);

AOI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_2093),
.A2(n_2089),
.B(n_985),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2094),
.Y(n_2097)
);

OAI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2095),
.A2(n_1999),
.B1(n_1998),
.B2(n_2021),
.Y(n_2098)
);

NOR2x1p5_ASAP7_75t_L g2099 ( 
.A(n_2093),
.B(n_1172),
.Y(n_2099)
);

AOI211xp5_ASAP7_75t_SL g2100 ( 
.A1(n_2093),
.A2(n_2037),
.B(n_1999),
.C(n_1998),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2093),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2093),
.B(n_1987),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2093),
.Y(n_2103)
);

NAND3xp33_ASAP7_75t_L g2104 ( 
.A(n_2093),
.B(n_1140),
.C(n_1136),
.Y(n_2104)
);

AOI31xp33_ASAP7_75t_L g2105 ( 
.A1(n_2093),
.A2(n_2034),
.A3(n_964),
.B(n_2006),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2093),
.Y(n_2106)
);

AOI211xp5_ASAP7_75t_L g2107 ( 
.A1(n_2093),
.A2(n_2006),
.B(n_2002),
.C(n_2003),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_SL g2108 ( 
.A(n_2093),
.B(n_2000),
.Y(n_2108)
);

NAND5xp2_ASAP7_75t_L g2109 ( 
.A(n_2108),
.B(n_2003),
.C(n_2050),
.D(n_2048),
.E(n_1418),
.Y(n_2109)
);

NOR2x1_ASAP7_75t_L g2110 ( 
.A(n_2101),
.B(n_1172),
.Y(n_2110)
);

NAND4xp25_ASAP7_75t_L g2111 ( 
.A(n_2097),
.B(n_2048),
.C(n_2050),
.D(n_2004),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_2102),
.B(n_1987),
.Y(n_2112)
);

NOR3xp33_ASAP7_75t_L g2113 ( 
.A(n_2103),
.B(n_2106),
.C(n_2096),
.Y(n_2113)
);

NOR2x1_ASAP7_75t_L g2114 ( 
.A(n_2099),
.B(n_1404),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2104),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2107),
.B(n_2002),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2100),
.B(n_1994),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2105),
.Y(n_2118)
);

AND5x1_ASAP7_75t_L g2119 ( 
.A(n_2098),
.B(n_2006),
.C(n_7),
.D(n_4),
.E(n_6),
.Y(n_2119)
);

NOR3x1_ASAP7_75t_L g2120 ( 
.A(n_2102),
.B(n_1993),
.C(n_1992),
.Y(n_2120)
);

OAI211xp5_ASAP7_75t_L g2121 ( 
.A1(n_2101),
.A2(n_1140),
.B(n_1136),
.C(n_1407),
.Y(n_2121)
);

NAND4xp75_ASAP7_75t_L g2122 ( 
.A(n_2101),
.B(n_1442),
.C(n_1440),
.D(n_1427),
.Y(n_2122)
);

NAND3xp33_ASAP7_75t_L g2123 ( 
.A(n_2108),
.B(n_1140),
.C(n_914),
.Y(n_2123)
);

NOR2x1_ASAP7_75t_L g2124 ( 
.A(n_2101),
.B(n_1422),
.Y(n_2124)
);

NAND3xp33_ASAP7_75t_L g2125 ( 
.A(n_2108),
.B(n_1140),
.C(n_916),
.Y(n_2125)
);

NOR4xp25_ASAP7_75t_L g2126 ( 
.A(n_2101),
.B(n_1993),
.C(n_917),
.D(n_918),
.Y(n_2126)
);

NOR3xp33_ASAP7_75t_L g2127 ( 
.A(n_2101),
.B(n_924),
.C(n_913),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2108),
.B(n_1994),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2102),
.Y(n_2129)
);

NOR3xp33_ASAP7_75t_L g2130 ( 
.A(n_2101),
.B(n_926),
.C(n_925),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_2102),
.B(n_2017),
.Y(n_2131)
);

NAND4xp25_ASAP7_75t_L g2132 ( 
.A(n_2108),
.B(n_935),
.C(n_940),
.D(n_928),
.Y(n_2132)
);

NOR2x1_ASAP7_75t_L g2133 ( 
.A(n_2101),
.B(n_1098),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2108),
.B(n_2001),
.Y(n_2134)
);

NAND3xp33_ASAP7_75t_L g2135 ( 
.A(n_2108),
.B(n_946),
.C(n_942),
.Y(n_2135)
);

NAND4xp25_ASAP7_75t_L g2136 ( 
.A(n_2108),
.B(n_948),
.C(n_949),
.D(n_947),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2108),
.B(n_2001),
.Y(n_2137)
);

NOR3xp33_ASAP7_75t_L g2138 ( 
.A(n_2101),
.B(n_953),
.C(n_950),
.Y(n_2138)
);

NOR3xp33_ASAP7_75t_L g2139 ( 
.A(n_2101),
.B(n_954),
.C(n_1098),
.Y(n_2139)
);

BUFx2_ASAP7_75t_L g2140 ( 
.A(n_2102),
.Y(n_2140)
);

NAND4xp25_ASAP7_75t_SL g2141 ( 
.A(n_2107),
.B(n_10),
.C(n_4),
.D(n_7),
.Y(n_2141)
);

NOR3xp33_ASAP7_75t_L g2142 ( 
.A(n_2101),
.B(n_1447),
.C(n_1445),
.Y(n_2142)
);

NAND3x1_ASAP7_75t_L g2143 ( 
.A(n_2096),
.B(n_10),
.C(n_11),
.Y(n_2143)
);

NAND4xp75_ASAP7_75t_L g2144 ( 
.A(n_2101),
.B(n_1458),
.C(n_1464),
.D(n_1451),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2108),
.B(n_2017),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2108),
.B(n_2017),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2102),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2108),
.B(n_2017),
.Y(n_2148)
);

NOR2x1_ASAP7_75t_L g2149 ( 
.A(n_2101),
.B(n_1546),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2108),
.B(n_1927),
.Y(n_2150)
);

NOR2xp67_ASAP7_75t_L g2151 ( 
.A(n_2102),
.B(n_14),
.Y(n_2151)
);

OAI211xp5_ASAP7_75t_SL g2152 ( 
.A1(n_2129),
.A2(n_1165),
.B(n_1176),
.C(n_1170),
.Y(n_2152)
);

AOI211x1_ASAP7_75t_L g2153 ( 
.A1(n_2141),
.A2(n_18),
.B(n_15),
.C(n_16),
.Y(n_2153)
);

AO21x1_ASAP7_75t_L g2154 ( 
.A1(n_2113),
.A2(n_15),
.B(n_18),
.Y(n_2154)
);

NOR2xp67_ASAP7_75t_L g2155 ( 
.A(n_2109),
.B(n_19),
.Y(n_2155)
);

AOI221xp5_ASAP7_75t_L g2156 ( 
.A1(n_2134),
.A2(n_1102),
.B1(n_515),
.B2(n_516),
.C(n_511),
.Y(n_2156)
);

AOI22xp5_ASAP7_75t_L g2157 ( 
.A1(n_2137),
.A2(n_1913),
.B1(n_1904),
.B2(n_1180),
.Y(n_2157)
);

AOI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_2128),
.A2(n_1180),
.B1(n_1154),
.B2(n_1562),
.Y(n_2158)
);

OAI211xp5_ASAP7_75t_L g2159 ( 
.A1(n_2151),
.A2(n_2140),
.B(n_2147),
.C(n_2126),
.Y(n_2159)
);

AOI221x1_ASAP7_75t_L g2160 ( 
.A1(n_2127),
.A2(n_2138),
.B1(n_2130),
.B2(n_2142),
.C(n_2139),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_2112),
.B(n_19),
.Y(n_2161)
);

AOI221xp5_ASAP7_75t_L g2162 ( 
.A1(n_2116),
.A2(n_1102),
.B1(n_521),
.B2(n_524),
.C(n_517),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_2150),
.B(n_20),
.Y(n_2163)
);

AOI21xp5_ASAP7_75t_L g2164 ( 
.A1(n_2110),
.A2(n_1176),
.B(n_1170),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2120),
.B(n_2118),
.Y(n_2165)
);

AOI21xp33_ASAP7_75t_SL g2166 ( 
.A1(n_2123),
.A2(n_20),
.B(n_21),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2111),
.B(n_21),
.Y(n_2167)
);

NOR3xp33_ASAP7_75t_SL g2168 ( 
.A(n_2121),
.B(n_525),
.C(n_510),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_2132),
.B(n_23),
.Y(n_2169)
);

AOI21xp33_ASAP7_75t_L g2170 ( 
.A1(n_2149),
.A2(n_1176),
.B(n_25),
.Y(n_2170)
);

OAI211xp5_ASAP7_75t_SL g2171 ( 
.A1(n_2115),
.A2(n_1176),
.B(n_1287),
.C(n_1283),
.Y(n_2171)
);

AOI221xp5_ASAP7_75t_SL g2172 ( 
.A1(n_2145),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.C(n_30),
.Y(n_2172)
);

NAND4xp25_ASAP7_75t_L g2173 ( 
.A(n_2125),
.B(n_33),
.C(n_26),
.D(n_29),
.Y(n_2173)
);

AOI221xp5_ASAP7_75t_L g2174 ( 
.A1(n_2148),
.A2(n_1102),
.B1(n_533),
.B2(n_536),
.C(n_532),
.Y(n_2174)
);

AOI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_2143),
.A2(n_1577),
.B1(n_542),
.B2(n_544),
.Y(n_2175)
);

OAI211xp5_ASAP7_75t_L g2176 ( 
.A1(n_2124),
.A2(n_36),
.B(n_33),
.C(n_34),
.Y(n_2176)
);

AOI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_2146),
.A2(n_548),
.B1(n_550),
.B2(n_528),
.Y(n_2177)
);

AOI211xp5_ASAP7_75t_L g2178 ( 
.A1(n_2135),
.A2(n_40),
.B(n_34),
.C(n_36),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2114),
.Y(n_2179)
);

OAI211xp5_ASAP7_75t_SL g2180 ( 
.A1(n_2133),
.A2(n_1291),
.B(n_47),
.C(n_44),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_2136),
.B(n_45),
.Y(n_2181)
);

OAI211xp5_ASAP7_75t_L g2182 ( 
.A1(n_2131),
.A2(n_51),
.B(n_48),
.C(n_50),
.Y(n_2182)
);

AOI211x1_ASAP7_75t_L g2183 ( 
.A1(n_2119),
.A2(n_51),
.B(n_48),
.C(n_50),
.Y(n_2183)
);

OAI32xp33_ASAP7_75t_L g2184 ( 
.A1(n_2122),
.A2(n_1572),
.A3(n_1571),
.B1(n_56),
.B2(n_53),
.Y(n_2184)
);

BUFx2_ASAP7_75t_L g2185 ( 
.A(n_2144),
.Y(n_2185)
);

AOI211x1_ASAP7_75t_L g2186 ( 
.A1(n_2141),
.A2(n_57),
.B(n_54),
.C(n_56),
.Y(n_2186)
);

AO22x2_ASAP7_75t_L g2187 ( 
.A1(n_2129),
.A2(n_60),
.B1(n_54),
.B2(n_59),
.Y(n_2187)
);

NOR2x1p5_ASAP7_75t_L g2188 ( 
.A(n_2134),
.B(n_557),
.Y(n_2188)
);

AOI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_2151),
.A2(n_572),
.B(n_570),
.Y(n_2189)
);

OAI21xp33_ASAP7_75t_SL g2190 ( 
.A1(n_2111),
.A2(n_59),
.B(n_60),
.Y(n_2190)
);

OAI211xp5_ASAP7_75t_SL g2191 ( 
.A1(n_2129),
.A2(n_66),
.B(n_63),
.C(n_64),
.Y(n_2191)
);

OAI32xp33_ASAP7_75t_L g2192 ( 
.A1(n_2134),
.A2(n_68),
.A3(n_64),
.B1(n_67),
.B2(n_69),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2134),
.Y(n_2193)
);

AOI22xp33_ASAP7_75t_L g2194 ( 
.A1(n_2117),
.A2(n_1950),
.B1(n_1939),
.B2(n_1960),
.Y(n_2194)
);

OAI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_2134),
.A2(n_583),
.B(n_576),
.Y(n_2195)
);

INVx1_ASAP7_75t_SL g2196 ( 
.A(n_2112),
.Y(n_2196)
);

AO32x1_ASAP7_75t_L g2197 ( 
.A1(n_2129),
.A2(n_73),
.A3(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2117),
.Y(n_2198)
);

OAI211xp5_ASAP7_75t_L g2199 ( 
.A1(n_2151),
.A2(n_78),
.B(n_71),
.C(n_77),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2134),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2117),
.B(n_77),
.Y(n_2201)
);

XNOR2xp5_ASAP7_75t_L g2202 ( 
.A(n_2143),
.B(n_78),
.Y(n_2202)
);

NAND4xp75_ASAP7_75t_L g2203 ( 
.A(n_2151),
.B(n_82),
.C(n_80),
.D(n_81),
.Y(n_2203)
);

OAI211xp5_ASAP7_75t_SL g2204 ( 
.A1(n_2129),
.A2(n_84),
.B(n_80),
.C(n_83),
.Y(n_2204)
);

OAI211xp5_ASAP7_75t_L g2205 ( 
.A1(n_2151),
.A2(n_86),
.B(n_83),
.C(n_84),
.Y(n_2205)
);

AOI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_2117),
.A2(n_595),
.B1(n_598),
.B2(n_594),
.Y(n_2206)
);

OA22x2_ASAP7_75t_L g2207 ( 
.A1(n_2134),
.A2(n_1950),
.B1(n_88),
.B2(n_86),
.Y(n_2207)
);

OAI211xp5_ASAP7_75t_L g2208 ( 
.A1(n_2151),
.A2(n_91),
.B(n_87),
.C(n_89),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_2134),
.B(n_87),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2117),
.Y(n_2210)
);

OA22x2_ASAP7_75t_L g2211 ( 
.A1(n_2134),
.A2(n_94),
.B1(n_91),
.B2(n_92),
.Y(n_2211)
);

AOI22xp5_ASAP7_75t_SL g2212 ( 
.A1(n_2109),
.A2(n_610),
.B1(n_617),
.B2(n_607),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2117),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2117),
.B(n_92),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2134),
.Y(n_2215)
);

INVxp33_ASAP7_75t_SL g2216 ( 
.A(n_2151),
.Y(n_2216)
);

AOI221xp5_ASAP7_75t_L g2217 ( 
.A1(n_2141),
.A2(n_635),
.B1(n_639),
.B2(n_620),
.C(n_619),
.Y(n_2217)
);

NOR3xp33_ASAP7_75t_L g2218 ( 
.A(n_2140),
.B(n_1242),
.C(n_1051),
.Y(n_2218)
);

AOI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_2117),
.A2(n_644),
.B1(n_646),
.B2(n_643),
.Y(n_2219)
);

OAI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2134),
.A2(n_1940),
.B1(n_1935),
.B2(n_1946),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_SL g2221 ( 
.A1(n_2183),
.A2(n_652),
.B1(n_653),
.B2(n_650),
.Y(n_2221)
);

OAI211xp5_ASAP7_75t_L g2222 ( 
.A1(n_2190),
.A2(n_97),
.B(n_94),
.C(n_96),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2198),
.B(n_1935),
.Y(n_2223)
);

AOI22xp33_ASAP7_75t_SL g2224 ( 
.A1(n_2216),
.A2(n_1120),
.B1(n_659),
.B2(n_660),
.Y(n_2224)
);

AOI21xp5_ASAP7_75t_SL g2225 ( 
.A1(n_2202),
.A2(n_661),
.B(n_654),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2187),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2161),
.B(n_96),
.Y(n_2227)
);

NOR2xp67_ASAP7_75t_L g2228 ( 
.A(n_2199),
.B(n_99),
.Y(n_2228)
);

NAND3xp33_ASAP7_75t_L g2229 ( 
.A(n_2209),
.B(n_1120),
.C(n_670),
.Y(n_2229)
);

NAND4xp25_ASAP7_75t_L g2230 ( 
.A(n_2153),
.B(n_103),
.C(n_100),
.D(n_101),
.Y(n_2230)
);

NAND5xp2_ASAP7_75t_L g2231 ( 
.A(n_2193),
.B(n_104),
.C(n_100),
.D(n_103),
.E(n_107),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2211),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_2205),
.B(n_2208),
.Y(n_2233)
);

OAI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2210),
.A2(n_1935),
.B1(n_1946),
.B2(n_671),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2154),
.Y(n_2235)
);

AND3x4_ASAP7_75t_L g2236 ( 
.A(n_2155),
.B(n_104),
.C(n_107),
.Y(n_2236)
);

INVx1_ASAP7_75t_SL g2237 ( 
.A(n_2203),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_2207),
.Y(n_2238)
);

NOR2x1_ASAP7_75t_L g2239 ( 
.A(n_2159),
.B(n_109),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2187),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2197),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_2201),
.B(n_109),
.Y(n_2242)
);

NAND3xp33_ASAP7_75t_L g2243 ( 
.A(n_2214),
.B(n_673),
.C(n_667),
.Y(n_2243)
);

NAND4xp75_ASAP7_75t_L g2244 ( 
.A(n_2165),
.B(n_114),
.C(n_110),
.D(n_111),
.Y(n_2244)
);

INVx1_ASAP7_75t_SL g2245 ( 
.A(n_2167),
.Y(n_2245)
);

NOR3xp33_ASAP7_75t_L g2246 ( 
.A(n_2213),
.B(n_1242),
.C(n_1051),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2186),
.Y(n_2247)
);

NAND3xp33_ASAP7_75t_L g2248 ( 
.A(n_2172),
.B(n_691),
.C(n_684),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2163),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2197),
.Y(n_2250)
);

BUFx2_ASAP7_75t_L g2251 ( 
.A(n_2200),
.Y(n_2251)
);

INVx1_ASAP7_75t_SL g2252 ( 
.A(n_2196),
.Y(n_2252)
);

INVx5_ASAP7_75t_L g2253 ( 
.A(n_2185),
.Y(n_2253)
);

OAI21xp33_ASAP7_75t_L g2254 ( 
.A1(n_2215),
.A2(n_698),
.B(n_692),
.Y(n_2254)
);

INVx1_ASAP7_75t_SL g2255 ( 
.A(n_2212),
.Y(n_2255)
);

AOI22x1_ASAP7_75t_L g2256 ( 
.A1(n_2188),
.A2(n_702),
.B1(n_704),
.B2(n_700),
.Y(n_2256)
);

NAND4xp75_ASAP7_75t_L g2257 ( 
.A(n_2169),
.B(n_116),
.C(n_110),
.D(n_115),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2197),
.Y(n_2258)
);

AOI21xp5_ASAP7_75t_L g2259 ( 
.A1(n_2164),
.A2(n_708),
.B(n_706),
.Y(n_2259)
);

NAND3xp33_ASAP7_75t_SL g2260 ( 
.A(n_2182),
.B(n_712),
.C(n_711),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2178),
.B(n_117),
.Y(n_2261)
);

OAI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_2173),
.A2(n_718),
.B1(n_720),
.B2(n_713),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_2176),
.Y(n_2263)
);

INVx1_ASAP7_75t_SL g2264 ( 
.A(n_2179),
.Y(n_2264)
);

NOR3xp33_ASAP7_75t_L g2265 ( 
.A(n_2152),
.B(n_1072),
.C(n_1048),
.Y(n_2265)
);

NOR3xp33_ASAP7_75t_L g2266 ( 
.A(n_2181),
.B(n_1072),
.C(n_1048),
.Y(n_2266)
);

NAND2x1p5_ASAP7_75t_L g2267 ( 
.A(n_2175),
.B(n_1090),
.Y(n_2267)
);

AOI211xp5_ASAP7_75t_L g2268 ( 
.A1(n_2166),
.A2(n_123),
.B(n_120),
.C(n_122),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2191),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2157),
.B(n_124),
.Y(n_2270)
);

INVxp67_ASAP7_75t_SL g2271 ( 
.A(n_2189),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2217),
.B(n_125),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_2160),
.B(n_2168),
.Y(n_2273)
);

NOR3x1_ASAP7_75t_L g2274 ( 
.A(n_2195),
.B(n_126),
.C(n_127),
.Y(n_2274)
);

NAND4xp25_ASAP7_75t_L g2275 ( 
.A(n_2170),
.B(n_128),
.C(n_126),
.D(n_127),
.Y(n_2275)
);

OAI322xp33_ASAP7_75t_L g2276 ( 
.A1(n_2252),
.A2(n_2219),
.A3(n_2206),
.B1(n_2177),
.B2(n_2158),
.C1(n_2171),
.C2(n_2180),
.Y(n_2276)
);

OR2x2_ASAP7_75t_L g2277 ( 
.A(n_2230),
.B(n_2275),
.Y(n_2277)
);

NAND3xp33_ASAP7_75t_SL g2278 ( 
.A(n_2236),
.B(n_2237),
.C(n_2235),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2242),
.Y(n_2279)
);

NAND3xp33_ASAP7_75t_SL g2280 ( 
.A(n_2264),
.B(n_2156),
.C(n_2162),
.Y(n_2280)
);

NAND3xp33_ASAP7_75t_SL g2281 ( 
.A(n_2268),
.B(n_2250),
.C(n_2241),
.Y(n_2281)
);

NOR2xp67_ASAP7_75t_L g2282 ( 
.A(n_2231),
.B(n_2204),
.Y(n_2282)
);

NAND5xp2_ASAP7_75t_L g2283 ( 
.A(n_2233),
.B(n_2232),
.C(n_2247),
.D(n_2269),
.E(n_2222),
.Y(n_2283)
);

NOR3xp33_ASAP7_75t_SL g2284 ( 
.A(n_2262),
.B(n_2174),
.C(n_2184),
.Y(n_2284)
);

NAND3x1_ASAP7_75t_L g2285 ( 
.A(n_2239),
.B(n_2218),
.C(n_2192),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2244),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2238),
.B(n_2194),
.Y(n_2287)
);

OAI222xp33_ASAP7_75t_L g2288 ( 
.A1(n_2251),
.A2(n_2220),
.B1(n_130),
.B2(n_131),
.C1(n_133),
.C2(n_134),
.Y(n_2288)
);

NAND3xp33_ASAP7_75t_L g2289 ( 
.A(n_2253),
.B(n_2263),
.C(n_2258),
.Y(n_2289)
);

AOI221xp5_ASAP7_75t_L g2290 ( 
.A1(n_2226),
.A2(n_2240),
.B1(n_2234),
.B2(n_2225),
.C(n_2260),
.Y(n_2290)
);

NAND3xp33_ASAP7_75t_L g2291 ( 
.A(n_2253),
.B(n_1090),
.C(n_136),
.Y(n_2291)
);

NAND3xp33_ASAP7_75t_SL g2292 ( 
.A(n_2227),
.B(n_1018),
.C(n_1011),
.Y(n_2292)
);

XNOR2xp5_ASAP7_75t_L g2293 ( 
.A(n_2257),
.B(n_143),
.Y(n_2293)
);

NAND4xp25_ASAP7_75t_L g2294 ( 
.A(n_2228),
.B(n_1128),
.C(n_1304),
.D(n_1301),
.Y(n_2294)
);

O2A1O1Ixp33_ASAP7_75t_L g2295 ( 
.A1(n_2261),
.A2(n_1372),
.B(n_1402),
.C(n_1388),
.Y(n_2295)
);

NOR3xp33_ASAP7_75t_L g2296 ( 
.A(n_2249),
.B(n_1383),
.C(n_1128),
.Y(n_2296)
);

AND5x1_ASAP7_75t_L g2297 ( 
.A(n_2259),
.B(n_1874),
.C(n_149),
.D(n_150),
.E(n_152),
.Y(n_2297)
);

NOR3xp33_ASAP7_75t_L g2298 ( 
.A(n_2221),
.B(n_1383),
.C(n_1372),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2253),
.A2(n_1939),
.B1(n_1938),
.B2(n_1517),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2223),
.Y(n_2300)
);

OAI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2245),
.A2(n_1506),
.B1(n_1524),
.B2(n_1517),
.Y(n_2301)
);

AOI32xp33_ASAP7_75t_L g2302 ( 
.A1(n_2255),
.A2(n_1523),
.A3(n_1537),
.B1(n_1579),
.B2(n_1560),
.Y(n_2302)
);

AOI22xp33_ASAP7_75t_L g2303 ( 
.A1(n_2273),
.A2(n_1939),
.B1(n_1938),
.B2(n_1534),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2274),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2272),
.B(n_148),
.Y(n_2305)
);

INVxp67_ASAP7_75t_SL g2306 ( 
.A(n_2270),
.Y(n_2306)
);

AOI221xp5_ASAP7_75t_L g2307 ( 
.A1(n_2248),
.A2(n_1534),
.B1(n_1574),
.B2(n_1568),
.C(n_1524),
.Y(n_2307)
);

AND3x1_ASAP7_75t_L g2308 ( 
.A(n_2246),
.B(n_1402),
.C(n_1388),
.Y(n_2308)
);

NAND5xp2_ASAP7_75t_L g2309 ( 
.A(n_2224),
.B(n_1872),
.C(n_160),
.D(n_163),
.E(n_174),
.Y(n_2309)
);

NOR2x1p5_ASAP7_75t_L g2310 ( 
.A(n_2271),
.B(n_1320),
.Y(n_2310)
);

OAI21xp33_ASAP7_75t_L g2311 ( 
.A1(n_2273),
.A2(n_1534),
.B(n_1524),
.Y(n_2311)
);

NAND3xp33_ASAP7_75t_L g2312 ( 
.A(n_2229),
.B(n_1452),
.C(n_1308),
.Y(n_2312)
);

INVxp33_ASAP7_75t_SL g2313 ( 
.A(n_2256),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2267),
.Y(n_2314)
);

BUFx2_ASAP7_75t_L g2315 ( 
.A(n_2243),
.Y(n_2315)
);

NOR4xp75_ASAP7_75t_L g2316 ( 
.A(n_2254),
.B(n_159),
.C(n_177),
.D(n_178),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2266),
.B(n_183),
.Y(n_2317)
);

NAND3xp33_ASAP7_75t_SL g2318 ( 
.A(n_2265),
.B(n_1325),
.C(n_1322),
.Y(n_2318)
);

OAI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2230),
.A2(n_1460),
.B1(n_1579),
.B2(n_1537),
.C(n_1554),
.Y(n_2319)
);

AOI22xp33_ASAP7_75t_SL g2320 ( 
.A1(n_2251),
.A2(n_1574),
.B1(n_1568),
.B2(n_1585),
.Y(n_2320)
);

OAI211xp5_ASAP7_75t_L g2321 ( 
.A1(n_2222),
.A2(n_1486),
.B(n_1484),
.C(n_1334),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2293),
.Y(n_2322)
);

O2A1O1Ixp33_ASAP7_75t_L g2323 ( 
.A1(n_2281),
.A2(n_1486),
.B(n_1484),
.C(n_1327),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_2286),
.B(n_184),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2282),
.B(n_188),
.Y(n_2325)
);

INVxp67_ASAP7_75t_L g2326 ( 
.A(n_2283),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2304),
.B(n_1939),
.Y(n_2327)
);

OAI211xp5_ASAP7_75t_L g2328 ( 
.A1(n_2290),
.A2(n_1331),
.B(n_1249),
.C(n_1250),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2277),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2305),
.B(n_189),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2310),
.Y(n_2331)
);

OAI22xp5_ASAP7_75t_SL g2332 ( 
.A1(n_2313),
.A2(n_1460),
.B1(n_1332),
.B2(n_1319),
.Y(n_2332)
);

AOI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2278),
.A2(n_2287),
.B1(n_2279),
.B2(n_2306),
.Y(n_2333)
);

NOR4xp25_ASAP7_75t_L g2334 ( 
.A(n_2280),
.B(n_1420),
.C(n_1426),
.D(n_1453),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2300),
.Y(n_2335)
);

NOR3xp33_ASAP7_75t_L g2336 ( 
.A(n_2294),
.B(n_1253),
.C(n_1248),
.Y(n_2336)
);

NAND2x1_ASAP7_75t_SL g2337 ( 
.A(n_2314),
.B(n_1016),
.Y(n_2337)
);

OA22x2_ASAP7_75t_L g2338 ( 
.A1(n_2311),
.A2(n_1511),
.B1(n_1504),
.B2(n_1510),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2291),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2284),
.B(n_2315),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2285),
.Y(n_2341)
);

OA22x2_ASAP7_75t_L g2342 ( 
.A1(n_2321),
.A2(n_2317),
.B1(n_2301),
.B2(n_2288),
.Y(n_2342)
);

OAI22xp5_ASAP7_75t_SL g2343 ( 
.A1(n_2320),
.A2(n_1288),
.B1(n_1308),
.B2(n_1318),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_2316),
.B(n_192),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2276),
.B(n_193),
.Y(n_2345)
);

BUFx2_ASAP7_75t_L g2346 ( 
.A(n_2308),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2319),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2295),
.Y(n_2348)
);

OAI222xp33_ASAP7_75t_L g2349 ( 
.A1(n_2302),
.A2(n_1532),
.B1(n_1560),
.B2(n_1554),
.C1(n_1467),
.C2(n_1466),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2312),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_2297),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2309),
.Y(n_2352)
);

AO22x2_ASAP7_75t_L g2353 ( 
.A1(n_2296),
.A2(n_2318),
.B1(n_2292),
.B2(n_2298),
.Y(n_2353)
);

NAND4xp75_ASAP7_75t_L g2354 ( 
.A(n_2307),
.B(n_1467),
.C(n_1466),
.D(n_1462),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2299),
.Y(n_2355)
);

INVxp33_ASAP7_75t_SL g2356 ( 
.A(n_2303),
.Y(n_2356)
);

OAI22xp5_ASAP7_75t_L g2357 ( 
.A1(n_2289),
.A2(n_1441),
.B1(n_1462),
.B2(n_1459),
.Y(n_2357)
);

AOI22xp33_ASAP7_75t_SL g2358 ( 
.A1(n_2289),
.A2(n_1332),
.B1(n_1288),
.B2(n_1318),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2293),
.Y(n_2359)
);

INVx1_ASAP7_75t_SL g2360 ( 
.A(n_2277),
.Y(n_2360)
);

BUFx2_ASAP7_75t_L g2361 ( 
.A(n_2304),
.Y(n_2361)
);

OAI22xp5_ASAP7_75t_SL g2362 ( 
.A1(n_2293),
.A2(n_1319),
.B1(n_1288),
.B2(n_1308),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_2286),
.B(n_194),
.Y(n_2363)
);

NOR2x1p5_ASAP7_75t_L g2364 ( 
.A(n_2281),
.B(n_1318),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2325),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2330),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2361),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2344),
.B(n_196),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2335),
.Y(n_2369)
);

NOR3xp33_ASAP7_75t_L g2370 ( 
.A(n_2326),
.B(n_2345),
.C(n_2329),
.Y(n_2370)
);

NOR4xp25_ASAP7_75t_L g2371 ( 
.A(n_2360),
.B(n_1017),
.C(n_1021),
.D(n_1023),
.Y(n_2371)
);

OAI22xp5_ASAP7_75t_SL g2372 ( 
.A1(n_2362),
.A2(n_1319),
.B1(n_1332),
.B2(n_1132),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2351),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2352),
.B(n_1938),
.Y(n_2374)
);

NAND5xp2_ASAP7_75t_L g2375 ( 
.A(n_2333),
.B(n_201),
.C(n_202),
.D(n_203),
.E(n_205),
.Y(n_2375)
);

OR3x2_ASAP7_75t_L g2376 ( 
.A(n_2322),
.B(n_206),
.C(n_208),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_2341),
.B(n_1121),
.Y(n_2377)
);

OAI222xp33_ASAP7_75t_L g2378 ( 
.A1(n_2342),
.A2(n_1459),
.B1(n_1449),
.B2(n_1446),
.C1(n_1441),
.C2(n_1436),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2324),
.Y(n_2379)
);

INVxp67_ASAP7_75t_L g2380 ( 
.A(n_2340),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2363),
.Y(n_2381)
);

AOI22xp33_ASAP7_75t_SL g2382 ( 
.A1(n_2327),
.A2(n_1132),
.B1(n_1121),
.B2(n_1122),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2359),
.B(n_1122),
.Y(n_2383)
);

NOR4xp25_ASAP7_75t_L g2384 ( 
.A(n_2328),
.B(n_1449),
.C(n_1446),
.D(n_1436),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2338),
.Y(n_2385)
);

AOI22xp5_ASAP7_75t_L g2386 ( 
.A1(n_2347),
.A2(n_1431),
.B1(n_1158),
.B2(n_1129),
.Y(n_2386)
);

AOI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_2356),
.A2(n_1132),
.B1(n_1130),
.B2(n_1129),
.Y(n_2387)
);

OAI222xp33_ASAP7_75t_L g2388 ( 
.A1(n_2339),
.A2(n_1082),
.B1(n_1081),
.B2(n_1043),
.C1(n_218),
.C2(n_219),
.Y(n_2388)
);

OA22x2_ASAP7_75t_L g2389 ( 
.A1(n_2355),
.A2(n_1944),
.B1(n_1092),
.B2(n_213),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_2364),
.Y(n_2390)
);

AOI22xp33_ASAP7_75t_SL g2391 ( 
.A1(n_2346),
.A2(n_1129),
.B1(n_1130),
.B2(n_1583),
.Y(n_2391)
);

AND2x4_ASAP7_75t_L g2392 ( 
.A(n_2331),
.B(n_223),
.Y(n_2392)
);

AOI22xp33_ASAP7_75t_L g2393 ( 
.A1(n_2350),
.A2(n_1130),
.B1(n_1240),
.B2(n_1189),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2337),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2376),
.Y(n_2395)
);

XNOR2xp5_ASAP7_75t_L g2396 ( 
.A(n_2373),
.B(n_2370),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2367),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_2369),
.B(n_2348),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2368),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2392),
.Y(n_2400)
);

OR2x2_ASAP7_75t_L g2401 ( 
.A(n_2375),
.B(n_2334),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2380),
.Y(n_2402)
);

AO21x2_ASAP7_75t_L g2403 ( 
.A1(n_2377),
.A2(n_2336),
.B(n_2357),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2389),
.Y(n_2404)
);

INVx3_ASAP7_75t_SL g2405 ( 
.A(n_2379),
.Y(n_2405)
);

INVx2_ASAP7_75t_SL g2406 ( 
.A(n_2381),
.Y(n_2406)
);

NOR3xp33_ASAP7_75t_L g2407 ( 
.A(n_2365),
.B(n_2323),
.C(n_2358),
.Y(n_2407)
);

AO22x2_ASAP7_75t_L g2408 ( 
.A1(n_2366),
.A2(n_2354),
.B1(n_2353),
.B2(n_2332),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2390),
.Y(n_2409)
);

XNOR2xp5_ASAP7_75t_L g2410 ( 
.A(n_2394),
.B(n_2343),
.Y(n_2410)
);

AOI22x1_ASAP7_75t_L g2411 ( 
.A1(n_2385),
.A2(n_2349),
.B1(n_1277),
.B2(n_1276),
.Y(n_2411)
);

XOR2xp5_ASAP7_75t_L g2412 ( 
.A(n_2372),
.B(n_225),
.Y(n_2412)
);

INVx1_ASAP7_75t_SL g2413 ( 
.A(n_2383),
.Y(n_2413)
);

XNOR2xp5_ASAP7_75t_L g2414 ( 
.A(n_2384),
.B(n_230),
.Y(n_2414)
);

AOI22xp33_ASAP7_75t_L g2415 ( 
.A1(n_2397),
.A2(n_2374),
.B1(n_2391),
.B2(n_2393),
.Y(n_2415)
);

NAND4xp25_ASAP7_75t_L g2416 ( 
.A(n_2402),
.B(n_2382),
.C(n_2387),
.D(n_2386),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2414),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2396),
.Y(n_2418)
);

INVx3_ASAP7_75t_SL g2419 ( 
.A(n_2405),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2400),
.Y(n_2420)
);

AOI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2406),
.A2(n_2371),
.B1(n_2388),
.B2(n_2378),
.Y(n_2421)
);

BUFx3_ASAP7_75t_L g2422 ( 
.A(n_2398),
.Y(n_2422)
);

OR3x2_ASAP7_75t_L g2423 ( 
.A(n_2409),
.B(n_236),
.C(n_238),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2401),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2395),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2399),
.Y(n_2426)
);

INVx1_ASAP7_75t_SL g2427 ( 
.A(n_2404),
.Y(n_2427)
);

AOI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_2407),
.A2(n_1241),
.B1(n_1189),
.B2(n_1190),
.Y(n_2428)
);

NAND5xp2_ASAP7_75t_L g2429 ( 
.A(n_2412),
.B(n_239),
.C(n_242),
.D(n_244),
.E(n_249),
.Y(n_2429)
);

INVxp67_ASAP7_75t_SL g2430 ( 
.A(n_2410),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2411),
.Y(n_2431)
);

OA22x2_ASAP7_75t_L g2432 ( 
.A1(n_2419),
.A2(n_2413),
.B1(n_2408),
.B2(n_2403),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2422),
.B(n_253),
.Y(n_2433)
);

NOR3xp33_ASAP7_75t_L g2434 ( 
.A(n_2418),
.B(n_1218),
.C(n_1178),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_2427),
.A2(n_1487),
.B(n_1277),
.Y(n_2435)
);

OAI22xp5_ASAP7_75t_L g2436 ( 
.A1(n_2423),
.A2(n_1241),
.B1(n_1277),
.B2(n_1276),
.Y(n_2436)
);

AND3x1_ASAP7_75t_L g2437 ( 
.A(n_2420),
.B(n_262),
.C(n_264),
.Y(n_2437)
);

XNOR2xp5_ASAP7_75t_L g2438 ( 
.A(n_2424),
.B(n_2430),
.Y(n_2438)
);

OAI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2426),
.A2(n_1240),
.B1(n_1276),
.B2(n_1254),
.Y(n_2439)
);

INVx3_ASAP7_75t_SL g2440 ( 
.A(n_2425),
.Y(n_2440)
);

OAI22xp5_ASAP7_75t_L g2441 ( 
.A1(n_2417),
.A2(n_1240),
.B1(n_1254),
.B2(n_1247),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2421),
.Y(n_2442)
);

INVx4_ASAP7_75t_L g2443 ( 
.A(n_2431),
.Y(n_2443)
);

AND3x1_ASAP7_75t_L g2444 ( 
.A(n_2442),
.B(n_2415),
.C(n_2429),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2437),
.Y(n_2445)
);

AOI22xp33_ASAP7_75t_L g2446 ( 
.A1(n_2440),
.A2(n_2416),
.B1(n_2428),
.B2(n_1237),
.Y(n_2446)
);

XNOR2xp5_ASAP7_75t_L g2447 ( 
.A(n_2438),
.B(n_265),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2433),
.Y(n_2448)
);

BUFx2_ASAP7_75t_SL g2449 ( 
.A(n_2432),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2443),
.B(n_266),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2434),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2435),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2439),
.Y(n_2453)
);

AOI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_2444),
.A2(n_2441),
.B(n_2436),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2450),
.Y(n_2455)
);

AOI222xp33_ASAP7_75t_SL g2456 ( 
.A1(n_2455),
.A2(n_2445),
.B1(n_2448),
.B2(n_2451),
.C1(n_2452),
.C2(n_2453),
.Y(n_2456)
);

AOI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2454),
.A2(n_2449),
.B1(n_2446),
.B2(n_2447),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2457),
.B(n_2456),
.Y(n_2458)
);

OAI21xp5_ASAP7_75t_SL g2459 ( 
.A1(n_2457),
.A2(n_1254),
.B(n_1247),
.Y(n_2459)
);

OAI22xp33_ASAP7_75t_L g2460 ( 
.A1(n_2458),
.A2(n_1487),
.B1(n_1247),
.B2(n_1245),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2459),
.Y(n_2461)
);

AOI21xp5_ASAP7_75t_L g2462 ( 
.A1(n_2458),
.A2(n_1171),
.B(n_1169),
.Y(n_2462)
);

OR2x6_ASAP7_75t_L g2463 ( 
.A(n_2462),
.B(n_2461),
.Y(n_2463)
);

AOI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_2463),
.A2(n_2460),
.B(n_1210),
.Y(n_2464)
);

AOI211xp5_ASAP7_75t_L g2465 ( 
.A1(n_2464),
.A2(n_1245),
.B(n_1241),
.C(n_1237),
.Y(n_2465)
);


endmodule