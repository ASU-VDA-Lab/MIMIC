module fake_netlist_1_12722_n_474 (n_117, n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_16, n_13, n_113, n_95, n_120, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_118, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_474);
input n_117;
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_16;
input n_13;
input n_113;
input n_95;
input n_120;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_118;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_474;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_133;
wire n_149;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_245;
wire n_357;
wire n_260;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_158;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g122 ( .A(n_114), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_121), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_107), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_43), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_76), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_54), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_120), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_17), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_95), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_15), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_47), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_118), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_50), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_105), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_9), .Y(n_137) );
CKINVDCx14_ASAP7_75t_R g138 ( .A(n_74), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_29), .Y(n_140) );
INVx2_ASAP7_75t_SL g141 ( .A(n_60), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_16), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_6), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_71), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_111), .Y(n_145) );
NOR2xp67_ASAP7_75t_L g146 ( .A(n_35), .B(n_14), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_51), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_22), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_32), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_93), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_37), .Y(n_151) );
BUFx10_ASAP7_75t_L g152 ( .A(n_75), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_23), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_97), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_5), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_88), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_98), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_112), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_8), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_33), .Y(n_160) );
BUFx5_ASAP7_75t_L g161 ( .A(n_18), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_61), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_48), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_21), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_62), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_56), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_110), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_26), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_31), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_104), .Y(n_170) );
NOR2xp67_ASAP7_75t_L g171 ( .A(n_13), .B(n_39), .Y(n_171) );
BUFx10_ASAP7_75t_L g172 ( .A(n_108), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_41), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_83), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_2), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_0), .Y(n_176) );
BUFx10_ASAP7_75t_L g177 ( .A(n_79), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_25), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_78), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_96), .Y(n_180) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_58), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_82), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_63), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_77), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_49), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_113), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_109), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_45), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_115), .Y(n_189) );
BUFx10_ASAP7_75t_L g190 ( .A(n_64), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_101), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_24), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_116), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_128), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_143), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_168), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_137), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_123), .Y(n_198) );
BUFx2_ASAP7_75t_L g199 ( .A(n_159), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_166), .B(n_0), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_173), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
BUFx12f_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_172), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_183), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_172), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_173), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_177), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_141), .B(n_1), .Y(n_209) );
INVx6_ASAP7_75t_L g210 ( .A(n_177), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_161), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_173), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_161), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_194), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_195), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_203), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_199), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_210), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_197), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_202), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_198), .A2(n_181), .B1(n_185), .B2(n_176), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_204), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_200), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_210), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_209), .Y(n_225) );
NOR2xp33_ASAP7_75t_R g226 ( .A(n_206), .B(n_138), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_211), .Y(n_227) );
NOR2x1p5_ASAP7_75t_L g228 ( .A(n_208), .B(n_155), .Y(n_228) );
BUFx10_ASAP7_75t_L g229 ( .A(n_205), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_213), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_230), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_229), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_227), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_225), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_228), .Y(n_235) );
BUFx6f_ASAP7_75t_SL g236 ( .A(n_218), .Y(n_236) );
NAND2xp33_ASAP7_75t_SL g237 ( .A(n_226), .B(n_130), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_217), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_221), .Y(n_239) );
BUFx6f_ASAP7_75t_SL g240 ( .A(n_219), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_220), .B(n_190), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_222), .B(n_124), .Y(n_242) );
NAND3xp33_ASAP7_75t_L g243 ( .A(n_223), .B(n_133), .C(n_125), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_224), .B(n_126), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_216), .B(n_127), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_232), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_232), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_232), .B(n_129), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_238), .B(n_215), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_233), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_234), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_239), .A2(n_131), .B1(n_148), .B2(n_132), .Y(n_252) );
INVxp67_ASAP7_75t_SL g253 ( .A(n_244), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_243), .A2(n_178), .B1(n_184), .B2(n_214), .Y(n_254) );
OR2x4_ASAP7_75t_L g255 ( .A(n_240), .B(n_175), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_242), .B(n_190), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_235), .B(n_179), .Y(n_257) );
NAND2x1p5_ASAP7_75t_L g258 ( .A(n_245), .B(n_155), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_231), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_240), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_236), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_241), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_253), .Y(n_263) );
NAND2x1_ASAP7_75t_L g264 ( .A(n_246), .B(n_193), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_259), .A2(n_136), .B(n_135), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_254), .B(n_237), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_251), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_262), .B(n_139), .Y(n_268) );
OAI22xp33_ASAP7_75t_L g269 ( .A1(n_252), .A2(n_144), .B1(n_145), .B2(n_140), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_257), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_257), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_250), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g273 ( .A(n_260), .B(n_134), .Y(n_273) );
BUFx12f_ASAP7_75t_L g274 ( .A(n_249), .Y(n_274) );
NOR2xp33_ASAP7_75t_SL g275 ( .A(n_247), .B(n_147), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_250), .B(n_153), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_258), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_256), .B(n_154), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_249), .B(n_149), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_255), .B(n_150), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_248), .A2(n_174), .B(n_158), .C(n_160), .Y(n_281) );
NAND2x1_ASAP7_75t_L g282 ( .A(n_261), .B(n_193), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_272), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_267), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_276), .Y(n_285) );
INVx6_ASAP7_75t_L g286 ( .A(n_274), .Y(n_286) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_265), .A2(n_171), .B(n_146), .Y(n_287) );
INVxp67_ASAP7_75t_SL g288 ( .A(n_272), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_272), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_273), .Y(n_290) );
BUFx4f_ASAP7_75t_L g291 ( .A(n_270), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_271), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_264), .A2(n_142), .B(n_122), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_279), .B(n_3), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_282), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_266), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_268), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_278), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_281), .A2(n_180), .B(n_170), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_269), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_280), .Y(n_302) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_275), .A2(n_186), .B(n_161), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_275), .B(n_151), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_274), .Y(n_305) );
BUFx12f_ASAP7_75t_L g306 ( .A(n_274), .Y(n_306) );
INVx6_ASAP7_75t_L g307 ( .A(n_274), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_267), .Y(n_308) );
AOI22x1_ASAP7_75t_L g309 ( .A1(n_272), .A2(n_212), .B1(n_207), .B2(n_201), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_263), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_274), .Y(n_311) );
AO21x1_ASAP7_75t_L g312 ( .A1(n_266), .A2(n_161), .B(n_4), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_274), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_267), .Y(n_314) );
AO21x1_ASAP7_75t_L g315 ( .A1(n_304), .A2(n_6), .B(n_7), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_310), .Y(n_316) );
BUFx8_ASAP7_75t_L g317 ( .A(n_306), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_308), .Y(n_318) );
INVx5_ASAP7_75t_L g319 ( .A(n_286), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_290), .B(n_311), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_305), .Y(n_321) );
INVx6_ASAP7_75t_L g322 ( .A(n_286), .Y(n_322) );
CKINVDCx11_ASAP7_75t_R g323 ( .A(n_313), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_283), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_314), .Y(n_325) );
INVx6_ASAP7_75t_L g326 ( .A(n_307), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_297), .A2(n_169), .B(n_167), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_307), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_301), .A2(n_182), .B1(n_188), .B2(n_191), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_299), .A2(n_196), .B1(n_207), .B2(n_201), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_298), .Y(n_332) );
NOR2x1_ASAP7_75t_SL g333 ( .A(n_295), .B(n_196), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_298), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_299), .A2(n_196), .B1(n_207), .B2(n_201), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_291), .B(n_212), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_292), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_293), .A2(n_212), .B(n_10), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_302), .B(n_156), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_283), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_299), .A2(n_192), .B1(n_189), .B2(n_187), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_294), .B(n_157), .Y(n_342) );
INVx4_ASAP7_75t_L g343 ( .A(n_289), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_287), .Y(n_344) );
NOR2x1_ASAP7_75t_SL g345 ( .A(n_289), .B(n_11), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_288), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_287), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_312), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_296), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_303), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_309), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_290), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_290), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_284), .Y(n_357) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_344), .A2(n_347), .B(n_349), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_327), .B(n_162), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_346), .B(n_348), .Y(n_360) );
CKINVDCx12_ASAP7_75t_R g361 ( .A(n_317), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_318), .Y(n_362) );
NAND2xp33_ASAP7_75t_R g363 ( .A(n_356), .B(n_12), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_316), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_330), .B(n_163), .Y(n_365) );
NOR3xp33_ASAP7_75t_SL g366 ( .A(n_321), .B(n_165), .C(n_164), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_323), .Y(n_367) );
NAND3xp33_ASAP7_75t_L g368 ( .A(n_329), .B(n_19), .C(n_20), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_322), .Y(n_369) );
NOR2xp33_ASAP7_75t_R g370 ( .A(n_319), .B(n_28), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_333), .B(n_30), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_355), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_354), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_343), .Y(n_374) );
OR2x6_ASAP7_75t_L g375 ( .A(n_320), .B(n_34), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_357), .B(n_36), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_325), .B(n_119), .Y(n_377) );
XOR2xp5_ASAP7_75t_L g378 ( .A(n_355), .B(n_38), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_337), .B(n_334), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_346), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_350), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_332), .Y(n_382) );
NAND2xp33_ASAP7_75t_R g383 ( .A(n_328), .B(n_40), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_315), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_326), .Y(n_385) );
NOR2xp33_ASAP7_75t_R g386 ( .A(n_324), .B(n_42), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_342), .Y(n_387) );
OR2x6_ASAP7_75t_L g388 ( .A(n_336), .B(n_44), .Y(n_388) );
OR2x6_ASAP7_75t_L g389 ( .A(n_324), .B(n_46), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_339), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_345), .A2(n_52), .B1(n_53), .B2(n_55), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_341), .B(n_57), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_340), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_340), .B(n_59), .Y(n_395) );
INVx8_ASAP7_75t_L g396 ( .A(n_331), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_335), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_360), .B(n_351), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_364), .B(n_65), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_382), .B(n_66), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_380), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_362), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_373), .B(n_338), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_374), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_379), .B(n_67), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_390), .B(n_352), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_381), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_363), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_394), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_384), .B(n_72), .Y(n_410) );
AND2x4_ASAP7_75t_SL g411 ( .A(n_375), .B(n_73), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_372), .B(n_80), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_358), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_396), .A2(n_81), .B1(n_85), .B2(n_86), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_377), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_372), .B(n_87), .Y(n_416) );
INVx3_ASAP7_75t_L g417 ( .A(n_371), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_385), .B(n_89), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_370), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_389), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_361), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_383), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_376), .B(n_94), .Y(n_423) );
INVx3_ASAP7_75t_SL g424 ( .A(n_369), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_395), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_387), .B(n_99), .Y(n_426) );
OAI222xp33_ASAP7_75t_L g427 ( .A1(n_378), .A2(n_117), .B1(n_100), .B2(n_102), .C1(n_103), .C2(n_106), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_389), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_401), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_404), .B(n_367), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_398), .B(n_391), .Y(n_431) );
AND2x4_ASAP7_75t_SL g432 ( .A(n_421), .B(n_388), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_407), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_413), .B(n_397), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_409), .B(n_386), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_406), .B(n_368), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_417), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_415), .B(n_365), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_424), .B(n_359), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_403), .B(n_392), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_417), .Y(n_443) );
BUFx3_ASAP7_75t_L g444 ( .A(n_419), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_410), .Y(n_445) );
INVx4_ASAP7_75t_SL g446 ( .A(n_444), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_429), .B(n_428), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_434), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_445), .B(n_438), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_439), .B(n_425), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_443), .B(n_399), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_433), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_431), .B(n_400), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_440), .B(n_435), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_452), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_447), .B(n_430), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_448), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_456), .A2(n_432), .B1(n_454), .B2(n_453), .Y(n_458) );
AOI21xp33_ASAP7_75t_SL g459 ( .A1(n_457), .A2(n_446), .B(n_422), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_458), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_460), .A2(n_459), .B(n_449), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_461), .A2(n_441), .B1(n_436), .B2(n_455), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_462), .A2(n_411), .B1(n_437), .B2(n_408), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_463), .Y(n_464) );
NOR2x1p5_ASAP7_75t_L g465 ( .A(n_464), .B(n_426), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_465), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_466), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_467), .B(n_451), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_468), .Y(n_469) );
OAI21x1_ASAP7_75t_L g470 ( .A1(n_469), .A2(n_418), .B(n_416), .Y(n_470) );
AOI21xp33_ASAP7_75t_L g471 ( .A1(n_470), .A2(n_366), .B(n_412), .Y(n_471) );
AOI22xp5_ASAP7_75t_SL g472 ( .A1(n_471), .A2(n_393), .B1(n_423), .B2(n_405), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_472), .B(n_414), .Y(n_473) );
AOI211xp5_ASAP7_75t_L g474 ( .A1(n_473), .A2(n_427), .B(n_450), .C(n_442), .Y(n_474) );
endmodule