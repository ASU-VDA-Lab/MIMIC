module fake_netlist_5_1163_n_2878 (n_137, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_649, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_631, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_637, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_645, n_539, n_175, n_538, n_262, n_238, n_639, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2878);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_639;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2878;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2520;
wire n_2347;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_2434;
wire n_1884;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2529;
wire n_2195;
wire n_2698;
wire n_809;
wire n_931;
wire n_870;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2491;
wire n_2177;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2314;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2457;
wire n_2346;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2521;
wire n_2111;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2424;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1534;
wire n_1354;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_968;
wire n_912;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_762;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2393;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2471;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2377;
wire n_2080;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_990;
wire n_836;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2437;
wire n_2219;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2093;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_766;
wire n_1457;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_2160;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_703;
wire n_698;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1530;
wire n_1497;
wire n_2654;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_2129;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2447;
wire n_1813;
wire n_2343;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2552;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2505;
wire n_2438;
wire n_2427;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2335;
wire n_2135;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_2044;
wire n_1990;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_525),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_106),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_341),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_482),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_310),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_55),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_101),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_421),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_453),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_285),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_314),
.Y(n_671)
);

CKINVDCx16_ASAP7_75t_R g672 ( 
.A(n_653),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_567),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_400),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_573),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_36),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_205),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_275),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_119),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_340),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_294),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_392),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_122),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_240),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_78),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_302),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_214),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_172),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_541),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_301),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_644),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_212),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_94),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_279),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_110),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_345),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_162),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_608),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_79),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_384),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_21),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_8),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_268),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_35),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_304),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_595),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_610),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_18),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_469),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_242),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_17),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_577),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_362),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_184),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_625),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_503),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_638),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_514),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_543),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_481),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_216),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_546),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_28),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_552),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_650),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_463),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_22),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_73),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_109),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_32),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_244),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_275),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_216),
.Y(n_734)
);

CKINVDCx16_ASAP7_75t_R g735 ( 
.A(n_602),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_566),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_298),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_587),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_151),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_540),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_335),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_132),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_616),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_33),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_528),
.Y(n_745)
);

CKINVDCx16_ASAP7_75t_R g746 ( 
.A(n_6),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_183),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_22),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_51),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_343),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_136),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_561),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_621),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_582),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_492),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_210),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_635),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_297),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_145),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_81),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_241),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_185),
.Y(n_762)
);

BUFx5_ASAP7_75t_L g763 ( 
.A(n_402),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_62),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_550),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_604),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_628),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_589),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_226),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_607),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_202),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_36),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_1),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_636),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_580),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_468),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_596),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_39),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_594),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_32),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_110),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_484),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_383),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_238),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_272),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_456),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_603),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_306),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_515),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_152),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_440),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_15),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_425),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_651),
.Y(n_794)
);

BUFx10_ASAP7_75t_L g795 ( 
.A(n_574),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_23),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_284),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_531),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_659),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_572),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_297),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_466),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_129),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_18),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_300),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_257),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_220),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_441),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_487),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_305),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_530),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_563),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_385),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_245),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_527),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_55),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_615),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_194),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_355),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_379),
.Y(n_820)
);

BUFx10_ASAP7_75t_L g821 ( 
.A(n_221),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_553),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_501),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_631),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_337),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_600),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_63),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_510),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_643),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_138),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_97),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_660),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_557),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_590),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_66),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_493),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_347),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_498),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_439),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_279),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_371),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_558),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_264),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_248),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_551),
.Y(n_845)
);

BUFx10_ASAP7_75t_L g846 ( 
.A(n_458),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_511),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_238),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_586),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_614),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_411),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_237),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_258),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_599),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_5),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_131),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_97),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_598),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_188),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_200),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_559),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_562),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_94),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_431),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_344),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_630),
.Y(n_866)
);

BUFx10_ASAP7_75t_L g867 ( 
.A(n_346),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_470),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_29),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_116),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_161),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_606),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_521),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_612),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_25),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_494),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_295),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_483),
.Y(n_878)
);

BUFx2_ASAP7_75t_SL g879 ( 
.A(n_443),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_560),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_332),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_231),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_432),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_331),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_301),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_132),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_477),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_278),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_262),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_123),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_149),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_565),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_165),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_126),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_584),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_58),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_575),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_433),
.Y(n_898)
);

BUFx10_ASAP7_75t_L g899 ( 
.A(n_243),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_376),
.Y(n_900)
);

BUFx5_ASAP7_75t_L g901 ( 
.A(n_363),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_143),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_356),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_214),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_556),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_167),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_294),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_524),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_212),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_490),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_348),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_479),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_259),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_312),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_475),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_228),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_336),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_449),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_153),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_281),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_583),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_576),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_168),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_426),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_381),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_307),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_143),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_320),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_508),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_622),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_641),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_47),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_613),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_45),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_544),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_35),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_442),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_178),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_293),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_326),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_223),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_290),
.Y(n_942)
);

CKINVDCx16_ASAP7_75t_R g943 ( 
.A(n_266),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_455),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_471),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_243),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_14),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_280),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_23),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_545),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_273),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_308),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_365),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_160),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_260),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_228),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_382),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_136),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_184),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_486),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_53),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_532),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_311),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_195),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_518),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_491),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_459),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_59),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_256),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_649),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_640),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_200),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_290),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_624),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_597),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_241),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_299),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_548),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_634),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_321),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_444),
.Y(n_981)
);

BUFx10_ASAP7_75t_L g982 ( 
.A(n_424),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_529),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_465),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_126),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_639),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_57),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_286),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_537),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_107),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_284),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_517),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_60),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_637),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_648),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_260),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_324),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_182),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_164),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_124),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_250),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_533),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_522),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_14),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_159),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_611),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_617),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_389),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_234),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_538),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_367),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_547),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_239),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_201),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_569),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_27),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_581),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_113),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_534),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_627),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_497),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_536),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_454),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_380),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_58),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_233),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_265),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_513),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_618),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_579),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_496),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_117),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_309),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_293),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_286),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_438),
.Y(n_1036)
);

BUFx10_ASAP7_75t_L g1037 ( 
.A(n_155),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_187),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_591),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_642),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_267),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_120),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_122),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_288),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_125),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_115),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_354),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_224),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_219),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_247),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_539),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_258),
.Y(n_1052)
);

CKINVDCx14_ASAP7_75t_R g1053 ( 
.A(n_240),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_554),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_109),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_489),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_73),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_619),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_67),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_605),
.Y(n_1060)
);

CKINVDCx14_ASAP7_75t_R g1061 ( 
.A(n_59),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_542),
.Y(n_1062)
);

CKINVDCx16_ASAP7_75t_R g1063 ( 
.A(n_163),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_209),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_570),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_40),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_592),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_207),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_127),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_193),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_265),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_632),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_124),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_63),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_395),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_645),
.Y(n_1076)
);

CKINVDCx16_ASAP7_75t_R g1077 ( 
.A(n_66),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_101),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_535),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_609),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_626),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_654),
.Y(n_1082)
);

INVxp33_ASAP7_75t_L g1083 ( 
.A(n_98),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_116),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_374),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_350),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_71),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_67),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_196),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_261),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_351),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_620),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_657),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_134),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_173),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_274),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_601),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_133),
.Y(n_1098)
);

BUFx5_ASAP7_75t_L g1099 ( 
.A(n_330),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_495),
.Y(n_1100)
);

BUFx10_ASAP7_75t_L g1101 ( 
.A(n_183),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_333),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_647),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_549),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_172),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_179),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_512),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_445),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_199),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_11),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_47),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_413),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_308),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_585),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_269),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_652),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_227),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_296),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_408),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_328),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_502),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_555),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_656),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_593),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_578),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_448),
.Y(n_1126)
);

CKINVDCx16_ASAP7_75t_R g1127 ( 
.A(n_255),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_306),
.Y(n_1128)
);

CKINVDCx16_ASAP7_75t_R g1129 ( 
.A(n_276),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_629),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_655),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_99),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_42),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_115),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_588),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_74),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_472),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_194),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_72),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_273),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_91),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_185),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_357),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_359),
.Y(n_1144)
);

INVxp67_ASAP7_75t_L g1145 ( 
.A(n_129),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_303),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_564),
.Y(n_1147)
);

CKINVDCx16_ASAP7_75t_R g1148 ( 
.A(n_153),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_161),
.Y(n_1149)
);

CKINVDCx16_ASAP7_75t_R g1150 ( 
.A(n_103),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_658),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_8),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_334),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_623),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_281),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_168),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_117),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_302),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_248),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_37),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_420),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_571),
.Y(n_1162)
);

CKINVDCx16_ASAP7_75t_R g1163 ( 
.A(n_313),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_646),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_226),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_407),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_81),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_500),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_633),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_436),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_76),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_182),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_77),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_688),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_688),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_688),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1053),
.B(n_0),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_746),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_666),
.Y(n_1179)
);

BUFx12f_ASAP7_75t_L g1180 ( 
.A(n_662),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1053),
.B(n_0),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_688),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_666),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_697),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1058),
.B(n_1),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_697),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1112),
.B(n_2),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_696),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_696),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1061),
.B(n_2),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_697),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_689),
.B(n_3),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_729),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_696),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_696),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_741),
.B(n_3),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1061),
.B(n_4),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_716),
.B(n_4),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_729),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_796),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_701),
.B(n_5),
.Y(n_1201)
);

INVx5_ASAP7_75t_L g1202 ( 
.A(n_697),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_943),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_857),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_701),
.B(n_6),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_980),
.B(n_7),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_857),
.Y(n_1207)
);

INVx5_ASAP7_75t_L g1208 ( 
.A(n_929),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1076),
.B(n_7),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_796),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_716),
.B(n_9),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1085),
.B(n_9),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1083),
.B(n_10),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1002),
.B(n_10),
.Y(n_1214)
);

INVx5_ASAP7_75t_L g1215 ( 
.A(n_929),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_857),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_857),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_727),
.B(n_11),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1103),
.B(n_12),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_727),
.B(n_12),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1116),
.B(n_776),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_802),
.B(n_13),
.Y(n_1222)
);

BUFx12f_ASAP7_75t_L g1223 ( 
.A(n_662),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_776),
.B(n_13),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_961),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_823),
.B(n_15),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1083),
.B(n_823),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_961),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_961),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_806),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_961),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1063),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_929),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_964),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_964),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_950),
.B(n_16),
.Y(n_1236)
);

XNOR2x1_ASAP7_75t_L g1237 ( 
.A(n_667),
.B(n_16),
.Y(n_1237)
);

BUFx8_ASAP7_75t_SL g1238 ( 
.A(n_860),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_950),
.B(n_17),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_970),
.B(n_19),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_970),
.B(n_19),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_981),
.B(n_20),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_802),
.B(n_20),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_932),
.B(n_21),
.Y(n_1244)
);

BUFx8_ASAP7_75t_L g1245 ( 
.A(n_985),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_964),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_981),
.B(n_24),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_806),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_827),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1024),
.B(n_24),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1024),
.B(n_25),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_SL g1252 ( 
.A(n_672),
.B(n_26),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_SL g1253 ( 
.A(n_735),
.B(n_26),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_964),
.Y(n_1254)
);

INVx5_ASAP7_75t_L g1255 ( 
.A(n_929),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1146),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1146),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_832),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1146),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_1031),
.Y(n_1260)
);

INVx5_ASAP7_75t_L g1261 ( 
.A(n_1031),
.Y(n_1261)
);

INVx5_ASAP7_75t_L g1262 ( 
.A(n_1031),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1028),
.B(n_27),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1146),
.Y(n_1264)
);

BUFx12f_ASAP7_75t_L g1265 ( 
.A(n_662),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_827),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1031),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_763),
.Y(n_1268)
);

INVx6_ASAP7_75t_L g1269 ( 
.A(n_795),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_763),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1028),
.B(n_28),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_832),
.B(n_29),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_914),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_834),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_763),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_834),
.B(n_30),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1001),
.B(n_30),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_914),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_987),
.B(n_969),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1001),
.B(n_31),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1074),
.B(n_31),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_969),
.B(n_33),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_850),
.B(n_876),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1152),
.Y(n_1284)
);

INVxp33_ASAP7_75t_SL g1285 ( 
.A(n_818),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_763),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_661),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1152),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_779),
.B(n_34),
.Y(n_1289)
);

BUFx12f_ASAP7_75t_L g1290 ( 
.A(n_685),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_850),
.B(n_34),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_876),
.B(n_37),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_997),
.Y(n_1293)
);

CKINVDCx11_ASAP7_75t_R g1294 ( 
.A(n_685),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1157),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_664),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_997),
.B(n_38),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_691),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1077),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1047),
.B(n_38),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1157),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1047),
.B(n_39),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1120),
.B(n_40),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1121),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_685),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_665),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1121),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1120),
.B(n_41),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_821),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_821),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1122),
.B(n_41),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1122),
.B(n_42),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_820),
.B(n_43),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_691),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_821),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1121),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_702),
.B(n_43),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_663),
.B(n_44),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_678),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_763),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1121),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_671),
.B(n_44),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_763),
.B(n_901),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_931),
.B(n_45),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_899),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_702),
.B(n_46),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_899),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_763),
.B(n_46),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1166),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_940),
.B(n_48),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_690),
.B(n_48),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_995),
.B(n_49),
.Y(n_1332)
);

INVx5_ASAP7_75t_L g1333 ( 
.A(n_1166),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1166),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_795),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_714),
.B(n_49),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_721),
.B(n_50),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1008),
.B(n_50),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_725),
.B(n_51),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_899),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_901),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_901),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_901),
.B(n_52),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_745),
.B(n_52),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_750),
.B(n_53),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_901),
.B(n_54),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1285),
.A2(n_975),
.B1(n_767),
.B2(n_1127),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1279),
.B(n_1163),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1175),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1176),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1174),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1185),
.A2(n_686),
.B1(n_694),
.B2(n_684),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1177),
.A2(n_1148),
.B1(n_1150),
.B2(n_1129),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1174),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1182),
.Y(n_1355)
);

AO22x2_ASAP7_75t_L g1356 ( 
.A1(n_1244),
.A2(n_891),
.B1(n_1115),
.B2(n_906),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1252),
.A2(n_1023),
.B1(n_674),
.B2(n_768),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1253),
.A2(n_1023),
.B1(n_833),
.B2(n_845),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1181),
.A2(n_998),
.B1(n_790),
.B2(n_848),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1279),
.B(n_795),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1258),
.B(n_846),
.Y(n_1361)
);

AO22x2_ASAP7_75t_L g1362 ( 
.A1(n_1244),
.A2(n_906),
.B1(n_1035),
.B2(n_705),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1182),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1197),
.A2(n_895),
.B1(n_915),
.B2(n_766),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1190),
.A2(n_882),
.B1(n_1057),
.B2(n_703),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1274),
.B(n_846),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1281),
.A2(n_1145),
.B1(n_801),
.B2(n_676),
.Y(n_1367)
);

AND2x2_ASAP7_75t_SL g1368 ( 
.A(n_1197),
.B(n_705),
.Y(n_1368)
);

AO22x2_ASAP7_75t_L g1369 ( 
.A1(n_1187),
.A2(n_1098),
.B1(n_1149),
.B2(n_1035),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1192),
.A2(n_925),
.B1(n_1056),
.B2(n_924),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1293),
.B(n_846),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1221),
.A2(n_1219),
.B1(n_1214),
.B2(n_1269),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1283),
.B(n_1287),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1296),
.B(n_867),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1335),
.B(n_1249),
.Y(n_1375)
);

AND2x2_ASAP7_75t_SL g1376 ( 
.A(n_1213),
.B(n_1098),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1196),
.A2(n_1164),
.B1(n_1065),
.B2(n_677),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1289),
.A2(n_683),
.B1(n_687),
.B2(n_670),
.Y(n_1378)
);

BUFx10_ASAP7_75t_L g1379 ( 
.A(n_1269),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1201),
.A2(n_695),
.B1(n_698),
.B2(n_693),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1188),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1194),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1178),
.B(n_1160),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1227),
.B(n_1019),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_R g1385 ( 
.A1(n_1305),
.A2(n_1171),
.B1(n_1167),
.B2(n_681),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1206),
.B(n_1067),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1205),
.A2(n_700),
.B1(n_706),
.B2(n_704),
.Y(n_1387)
);

INVx8_ASAP7_75t_L g1388 ( 
.A(n_1180),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1313),
.A2(n_711),
.B1(n_712),
.B2(n_709),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1324),
.A2(n_724),
.B1(n_732),
.B2(n_715),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1184),
.B(n_752),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1272),
.A2(n_734),
.B1(n_742),
.B2(n_733),
.Y(n_1392)
);

OAI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1292),
.A2(n_747),
.B1(n_748),
.B2(n_744),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1203),
.A2(n_751),
.B1(n_759),
.B2(n_749),
.Y(n_1394)
);

OA22x2_ASAP7_75t_L g1395 ( 
.A1(n_1179),
.A2(n_728),
.B1(n_730),
.B2(n_679),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1249),
.B(n_867),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1309),
.B(n_867),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1273),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1189),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1330),
.A2(n_764),
.B1(n_769),
.B2(n_762),
.Y(n_1400)
);

NAND3x1_ASAP7_75t_L g1401 ( 
.A(n_1213),
.B(n_737),
.C(n_731),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1302),
.A2(n_780),
.B1(n_781),
.B2(n_772),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1195),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1325),
.Y(n_1404)
);

AO22x2_ASAP7_75t_L g1405 ( 
.A1(n_1237),
.A2(n_1198),
.B1(n_1218),
.B2(n_1211),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1303),
.A2(n_785),
.B1(n_788),
.B2(n_784),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1327),
.B(n_982),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1232),
.A2(n_797),
.B1(n_803),
.B2(n_792),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1299),
.A2(n_807),
.B1(n_810),
.B2(n_804),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1305),
.B(n_982),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1332),
.A2(n_830),
.B1(n_831),
.B2(n_816),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1338),
.B(n_982),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1340),
.B(n_1119),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1340),
.B(n_1144),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1312),
.A2(n_844),
.B1(n_863),
.B2(n_843),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1273),
.B(n_1147),
.Y(n_1416)
);

NAND2xp33_ASAP7_75t_SL g1417 ( 
.A(n_1282),
.B(n_684),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1284),
.B(n_1168),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1284),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1223),
.B(n_1149),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1209),
.A2(n_1212),
.B1(n_1226),
.B2(n_1224),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1265),
.A2(n_1310),
.B1(n_1315),
.B2(n_1290),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1277),
.A2(n_871),
.B1(n_875),
.B2(n_870),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1280),
.A2(n_886),
.B1(n_888),
.B2(n_877),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1288),
.B(n_1295),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1288),
.B(n_1169),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1236),
.A2(n_694),
.B1(n_722),
.B2(n_686),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1295),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_SL g1429 ( 
.A(n_1183),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1220),
.A2(n_890),
.B1(n_893),
.B2(n_889),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1222),
.A2(n_902),
.B1(n_907),
.B2(n_894),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1301),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1204),
.Y(n_1433)
);

XNOR2xp5_ASAP7_75t_L g1434 ( 
.A(n_1282),
.B(n_1173),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1301),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1243),
.A2(n_913),
.B1(n_920),
.B2(n_909),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1242),
.A2(n_1250),
.B1(n_1263),
.B2(n_1247),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1276),
.A2(n_934),
.B1(n_936),
.B2(n_927),
.Y(n_1438)
);

AO22x2_ASAP7_75t_L g1439 ( 
.A1(n_1291),
.A2(n_1300),
.B1(n_1308),
.B2(n_1297),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1311),
.A2(n_939),
.B1(n_941),
.B2(n_938),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1328),
.A2(n_942),
.B1(n_947),
.B2(n_946),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1194),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1318),
.B(n_754),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1193),
.B(n_949),
.Y(n_1444)
);

OAI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1343),
.A2(n_952),
.B1(n_958),
.B2(n_955),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1322),
.B(n_777),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1228),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1239),
.A2(n_1241),
.B1(n_1251),
.B2(n_1240),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1346),
.A2(n_968),
.B1(n_972),
.B2(n_963),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1207),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1271),
.A2(n_988),
.B1(n_991),
.B2(n_976),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1199),
.A2(n_1004),
.B1(n_1009),
.B2(n_1000),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1331),
.A2(n_1018),
.B1(n_1026),
.B2(n_1014),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1207),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1216),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1200),
.A2(n_1032),
.B1(n_1033),
.B2(n_1027),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1184),
.B(n_783),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1210),
.B(n_1034),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1230),
.A2(n_1044),
.B1(n_1045),
.B2(n_1042),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1235),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1336),
.A2(n_1052),
.B1(n_1059),
.B2(n_1048),
.Y(n_1461)
);

INVx8_ASAP7_75t_L g1462 ( 
.A(n_1238),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1337),
.B(n_789),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1216),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1248),
.B(n_1037),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1294),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1217),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1339),
.A2(n_1071),
.B1(n_1078),
.B2(n_1064),
.Y(n_1468)
);

BUFx10_ASAP7_75t_L g1469 ( 
.A(n_1266),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1217),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1256),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1344),
.B(n_794),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1278),
.A2(n_1088),
.B1(n_1089),
.B2(n_1084),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1225),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1323),
.A2(n_1095),
.B1(n_1105),
.B2(n_1090),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1317),
.A2(n_1111),
.B1(n_1118),
.B2(n_1106),
.Y(n_1476)
);

AO22x2_ASAP7_75t_L g1477 ( 
.A1(n_1317),
.A2(n_756),
.B1(n_758),
.B2(n_739),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1345),
.A2(n_1245),
.B1(n_1133),
.B2(n_1134),
.Y(n_1478)
);

OAI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1326),
.A2(n_1136),
.B1(n_1139),
.B2(n_1128),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1306),
.A2(n_1141),
.B1(n_1142),
.B2(n_1140),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1326),
.A2(n_1159),
.B1(n_1156),
.B2(n_1172),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1319),
.A2(n_773),
.B1(n_840),
.B2(n_814),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1298),
.A2(n_954),
.B1(n_1173),
.B2(n_722),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1186),
.A2(n_859),
.B1(n_904),
.B2(n_856),
.Y(n_1484)
);

AO22x2_ASAP7_75t_L g1485 ( 
.A1(n_1298),
.A2(n_761),
.B1(n_771),
.B2(n_760),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1191),
.B(n_1037),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1259),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1225),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1229),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1260),
.A2(n_1038),
.B1(n_1069),
.B2(n_1055),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1267),
.A2(n_1094),
.B1(n_1117),
.B2(n_1110),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1268),
.A2(n_805),
.B1(n_835),
.B2(n_778),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1229),
.Y(n_1493)
);

XNOR2xp5_ASAP7_75t_L g1494 ( 
.A(n_1314),
.B(n_954),
.Y(n_1494)
);

OR2x6_ASAP7_75t_L g1495 ( 
.A(n_1314),
.B(n_852),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1231),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1270),
.A2(n_1132),
.B1(n_669),
.B2(n_673),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1231),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1342),
.A2(n_855),
.B1(n_869),
.B2(n_853),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1191),
.B(n_800),
.Y(n_1500)
);

AO22x2_ASAP7_75t_L g1501 ( 
.A1(n_1275),
.A2(n_885),
.B1(n_916),
.B2(n_896),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1234),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1202),
.B(n_1208),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1286),
.A2(n_675),
.B1(n_680),
.B2(n_668),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1202),
.B(n_1037),
.Y(n_1505)
);

AO22x2_ASAP7_75t_L g1506 ( 
.A1(n_1320),
.A2(n_919),
.B1(n_926),
.B2(n_923),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1208),
.B(n_1101),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1341),
.A2(n_692),
.B1(n_699),
.B2(n_682),
.Y(n_1508)
);

AO22x2_ASAP7_75t_L g1509 ( 
.A1(n_1234),
.A2(n_948),
.B1(n_956),
.B2(n_951),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1246),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1246),
.Y(n_1511)
);

OAI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1254),
.A2(n_1025),
.B1(n_1046),
.B2(n_996),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1254),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1257),
.A2(n_708),
.B1(n_710),
.B2(n_707),
.Y(n_1514)
);

OAI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1215),
.A2(n_973),
.B1(n_977),
.B2(n_959),
.Y(n_1515)
);

OA22x2_ASAP7_75t_L g1516 ( 
.A1(n_1257),
.A2(n_993),
.B1(n_999),
.B2(n_990),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1264),
.A2(n_717),
.B1(n_718),
.B2(n_713),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1264),
.A2(n_720),
.B1(n_723),
.B2(n_719),
.Y(n_1518)
);

OAI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1304),
.A2(n_1087),
.B1(n_1138),
.B2(n_1050),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1304),
.A2(n_736),
.B1(n_738),
.B2(n_726),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1215),
.A2(n_1013),
.B1(n_1016),
.B2(n_1005),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1233),
.B(n_1101),
.Y(n_1522)
);

OR2x6_ASAP7_75t_L g1523 ( 
.A(n_1307),
.B(n_1041),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1307),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1233),
.A2(n_1049),
.B1(n_1066),
.B2(n_1043),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1255),
.B(n_815),
.Y(n_1526)
);

NAND3x1_ASAP7_75t_L g1527 ( 
.A(n_1316),
.B(n_1070),
.C(n_1068),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1316),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1321),
.Y(n_1529)
);

INVx5_ASAP7_75t_L g1530 ( 
.A(n_1321),
.Y(n_1530)
);

AO22x2_ASAP7_75t_L g1531 ( 
.A1(n_1329),
.A2(n_1073),
.B1(n_1109),
.B2(n_1096),
.Y(n_1531)
);

AO22x2_ASAP7_75t_L g1532 ( 
.A1(n_1329),
.A2(n_1113),
.B1(n_1158),
.B2(n_1155),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1255),
.B(n_819),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1334),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1261),
.B(n_1101),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1334),
.Y(n_1536)
);

BUFx10_ASAP7_75t_L g1537 ( 
.A(n_1261),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1262),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1262),
.B(n_825),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1333),
.A2(n_743),
.B1(n_753),
.B2(n_740),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1333),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1175),
.Y(n_1542)
);

OAI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1252),
.A2(n_1165),
.B1(n_872),
.B2(n_922),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1279),
.B(n_755),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1279),
.B(n_757),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1285),
.A2(n_770),
.B1(n_774),
.B2(n_765),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1279),
.B(n_775),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1175),
.Y(n_1548)
);

OA22x2_ASAP7_75t_L g1549 ( 
.A1(n_1279),
.A2(n_829),
.B1(n_838),
.B2(n_826),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1175),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1175),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1174),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1285),
.A2(n_786),
.B1(n_787),
.B2(n_782),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1285),
.A2(n_793),
.B1(n_798),
.B2(n_791),
.Y(n_1554)
);

AOI22x1_ASAP7_75t_L g1555 ( 
.A1(n_1213),
.A2(n_808),
.B1(n_809),
.B2(n_799),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1252),
.A2(n_854),
.B1(n_858),
.B2(n_847),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1285),
.A2(n_812),
.B1(n_813),
.B2(n_811),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1174),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1285),
.A2(n_822),
.B1(n_824),
.B2(n_817),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1285),
.A2(n_836),
.B1(n_837),
.B2(n_828),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1175),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1175),
.Y(n_1562)
);

AO22x1_ASAP7_75t_SL g1563 ( 
.A1(n_1187),
.A2(n_883),
.B1(n_897),
.B2(n_864),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1273),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1285),
.A2(n_841),
.B1(n_842),
.B2(n_839),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1279),
.B(n_849),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1279),
.B(n_851),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1279),
.B(n_861),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1221),
.B(n_900),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1252),
.A2(n_918),
.B1(n_928),
.B2(n_910),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1258),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1285),
.A2(n_865),
.B1(n_866),
.B2(n_862),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1175),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_1287),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_R g1575 ( 
.A(n_1287),
.B(n_868),
.Y(n_1575)
);

OAI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1252),
.A2(n_933),
.B1(n_945),
.B2(n_930),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1279),
.B(n_873),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1252),
.A2(n_971),
.B1(n_979),
.B2(n_953),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1175),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1252),
.A2(n_984),
.B1(n_992),
.B2(n_983),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1174),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1285),
.A2(n_878),
.B1(n_880),
.B2(n_874),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_SL g1583 ( 
.A1(n_1285),
.A2(n_1020),
.B1(n_1022),
.B2(n_1007),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1252),
.A2(n_1039),
.B1(n_1051),
.B2(n_1036),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1287),
.B(n_1072),
.Y(n_1585)
);

OAI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1252),
.A2(n_1081),
.B1(n_1100),
.B2(n_1079),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1175),
.Y(n_1587)
);

XOR2xp5_ASAP7_75t_L g1588 ( 
.A(n_1237),
.B(n_881),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1175),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1285),
.A2(n_884),
.B1(n_892),
.B2(n_887),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1269),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1175),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1175),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1252),
.A2(n_1125),
.B1(n_1154),
.B2(n_1107),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1175),
.Y(n_1595)
);

AO22x2_ASAP7_75t_L g1596 ( 
.A1(n_1244),
.A2(n_879),
.B1(n_57),
.B2(n_54),
.Y(n_1596)
);

NAND3x1_ASAP7_75t_L g1597 ( 
.A(n_1185),
.B(n_56),
.C(n_60),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1175),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1175),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1174),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1285),
.A2(n_903),
.B1(n_905),
.B2(n_898),
.Y(n_1601)
);

OAI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1252),
.A2(n_911),
.B1(n_912),
.B2(n_908),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1175),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1252),
.A2(n_917),
.B1(n_935),
.B2(n_921),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1252),
.A2(n_944),
.B1(n_957),
.B2(n_937),
.Y(n_1605)
);

AO22x2_ASAP7_75t_L g1606 ( 
.A1(n_1244),
.A2(n_62),
.B1(n_56),
.B2(n_61),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1174),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1279),
.B(n_960),
.Y(n_1608)
);

OAI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1252),
.A2(n_965),
.B1(n_966),
.B2(n_962),
.Y(n_1609)
);

INVx5_ASAP7_75t_L g1610 ( 
.A(n_1269),
.Y(n_1610)
);

AO22x2_ASAP7_75t_L g1611 ( 
.A1(n_1244),
.A2(n_65),
.B1(n_61),
.B2(n_64),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1279),
.B(n_967),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1285),
.A2(n_978),
.B1(n_986),
.B2(n_974),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1175),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1252),
.A2(n_989),
.B1(n_1003),
.B2(n_994),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1279),
.B(n_1006),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1279),
.B(n_1010),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1252),
.A2(n_1011),
.B1(n_1015),
.B2(n_1012),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1279),
.B(n_1017),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1252),
.A2(n_1029),
.B1(n_1030),
.B2(n_1021),
.Y(n_1620)
);

OAI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1252),
.A2(n_1054),
.B1(n_1060),
.B2(n_1040),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1174),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1285),
.A2(n_1062),
.B1(n_1080),
.B2(n_1075),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1174),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1285),
.A2(n_1082),
.B1(n_1091),
.B2(n_1086),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1174),
.Y(n_1626)
);

AO22x2_ASAP7_75t_L g1627 ( 
.A1(n_1244),
.A2(n_68),
.B1(n_64),
.B2(n_65),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1285),
.A2(n_1092),
.B1(n_1097),
.B2(n_1093),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1285),
.A2(n_1104),
.B1(n_1108),
.B2(n_1102),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1175),
.Y(n_1630)
);

NAND3x1_ASAP7_75t_L g1631 ( 
.A(n_1185),
.B(n_68),
.C(n_69),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1269),
.Y(n_1632)
);

AO22x2_ASAP7_75t_L g1633 ( 
.A1(n_1244),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1633)
);

BUFx10_ASAP7_75t_L g1634 ( 
.A(n_1269),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1175),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1269),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1285),
.A2(n_1123),
.B1(n_1124),
.B2(n_1114),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1175),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1279),
.B(n_1126),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1285),
.A2(n_1131),
.B1(n_1135),
.B2(n_1130),
.Y(n_1640)
);

AO22x2_ASAP7_75t_L g1641 ( 
.A1(n_1244),
.A2(n_74),
.B1(n_70),
.B2(n_72),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1285),
.A2(n_1143),
.B1(n_1151),
.B2(n_1137),
.Y(n_1642)
);

AO22x2_ASAP7_75t_L g1643 ( 
.A1(n_1244),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1643)
);

NAND2xp33_ASAP7_75t_SL g1644 ( 
.A(n_1197),
.B(n_1166),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1273),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1175),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1175),
.Y(n_1647)
);

CKINVDCx6p67_ASAP7_75t_R g1648 ( 
.A(n_1294),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1252),
.A2(n_1161),
.B1(n_1162),
.B2(n_1153),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1174),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1285),
.A2(n_1170),
.B1(n_1099),
.B2(n_901),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1178),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1279),
.B(n_1099),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1285),
.A2(n_1099),
.B1(n_901),
.B2(n_79),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1279),
.B(n_1099),
.Y(n_1655)
);

AO22x2_ASAP7_75t_L g1656 ( 
.A1(n_1244),
.A2(n_80),
.B1(n_75),
.B2(n_78),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1279),
.B(n_1099),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1221),
.B(n_1099),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1174),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1279),
.B(n_1099),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1221),
.B(n_80),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1279),
.B(n_315),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1174),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_R g1664 ( 
.A1(n_1305),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1285),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1175),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1287),
.B(n_316),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1279),
.B(n_317),
.Y(n_1668)
);

OAI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1252),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1285),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1279),
.B(n_318),
.Y(n_1671)
);

OAI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1252),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1285),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1285),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1252),
.A2(n_95),
.B1(n_92),
.B2(n_93),
.Y(n_1675)
);

OA22x2_ASAP7_75t_L g1676 ( 
.A1(n_1279),
.A2(n_98),
.B1(n_95),
.B2(n_96),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1285),
.A2(n_100),
.B1(n_96),
.B2(n_99),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1285),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1252),
.A2(n_105),
.B1(n_102),
.B2(n_104),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1279),
.B(n_319),
.Y(n_1680)
);

OAI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1252),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1279),
.B(n_322),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1375),
.B(n_107),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1349),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1575),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1421),
.A2(n_325),
.B(n_323),
.Y(n_1686)
);

AND2x6_ASAP7_75t_L g1687 ( 
.A(n_1653),
.B(n_327),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1350),
.Y(n_1688)
);

XOR2xp5_ASAP7_75t_L g1689 ( 
.A(n_1574),
.B(n_1588),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1381),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1571),
.B(n_329),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1413),
.B(n_108),
.Y(n_1692)
);

XOR2x2_ASAP7_75t_L g1693 ( 
.A(n_1352),
.B(n_108),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1399),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1524),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1403),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1425),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1528),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1414),
.B(n_111),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1529),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1384),
.B(n_111),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1348),
.B(n_112),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1536),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1534),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1493),
.Y(n_1705)
);

XOR2xp5_ASAP7_75t_L g1706 ( 
.A(n_1357),
.B(n_338),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1496),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1502),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1510),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1538),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1351),
.Y(n_1711)
);

INVxp33_ASAP7_75t_L g1712 ( 
.A(n_1494),
.Y(n_1712)
);

XOR2xp5_ASAP7_75t_L g1713 ( 
.A(n_1358),
.B(n_339),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1354),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1355),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1396),
.B(n_112),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1363),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1382),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1442),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1450),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1433),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1454),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1455),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1464),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1467),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1470),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1412),
.B(n_113),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1474),
.Y(n_1728)
);

INVxp67_ASAP7_75t_SL g1729 ( 
.A(n_1398),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1513),
.Y(n_1730)
);

INVx4_ASAP7_75t_SL g1731 ( 
.A(n_1429),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1552),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1558),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1581),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1360),
.B(n_114),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1386),
.B(n_114),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1600),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1376),
.B(n_342),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1607),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1437),
.A2(n_1448),
.B(n_1368),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1622),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1543),
.B(n_118),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1624),
.Y(n_1743)
);

XNOR2xp5_ASAP7_75t_L g1744 ( 
.A(n_1370),
.B(n_1434),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1626),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1410),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1650),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1447),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1416),
.B(n_349),
.Y(n_1749)
);

INVxp67_ASAP7_75t_SL g1750 ( 
.A(n_1419),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1655),
.B(n_352),
.Y(n_1751)
);

OR2x6_ASAP7_75t_L g1752 ( 
.A(n_1462),
.B(n_118),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1663),
.Y(n_1753)
);

INVxp67_ASAP7_75t_SL g1754 ( 
.A(n_1428),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1397),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1460),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1471),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1488),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1487),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1542),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_1432),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1659),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1548),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1550),
.Y(n_1764)
);

XOR2xp5_ASAP7_75t_L g1765 ( 
.A(n_1364),
.B(n_353),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1652),
.Y(n_1766)
);

XOR2xp5_ASAP7_75t_L g1767 ( 
.A(n_1422),
.B(n_358),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1585),
.B(n_119),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1644),
.A2(n_1439),
.B(n_1443),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1657),
.B(n_360),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1602),
.B(n_120),
.Y(n_1771)
);

INVx4_ASAP7_75t_L g1772 ( 
.A(n_1530),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1551),
.Y(n_1773)
);

AOI21x1_ASAP7_75t_L g1774 ( 
.A1(n_1660),
.A2(n_364),
.B(n_361),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1407),
.B(n_121),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1561),
.Y(n_1776)
);

CKINVDCx14_ASAP7_75t_R g1777 ( 
.A(n_1648),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1662),
.A2(n_1680),
.B(n_1671),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1610),
.B(n_121),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1562),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1573),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1610),
.B(n_123),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1439),
.B(n_366),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1579),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1610),
.B(n_125),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1486),
.B(n_127),
.Y(n_1786)
);

NAND2xp33_ASAP7_75t_R g1787 ( 
.A(n_1383),
.B(n_1373),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1361),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1366),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1505),
.B(n_128),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1587),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1589),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1592),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1507),
.B(n_1522),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1535),
.B(n_128),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1593),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1595),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1605),
.B(n_130),
.Y(n_1798)
);

OR2x6_ASAP7_75t_L g1799 ( 
.A(n_1462),
.B(n_130),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1609),
.B(n_131),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1598),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1599),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1418),
.B(n_133),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1603),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1614),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1426),
.B(n_134),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1544),
.B(n_135),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1620),
.B(n_135),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1630),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1635),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1638),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1646),
.Y(n_1812)
);

INVxp33_ASAP7_75t_L g1813 ( 
.A(n_1394),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1647),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1666),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1435),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1498),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1659),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1511),
.Y(n_1819)
);

XOR2xp5_ASAP7_75t_L g1820 ( 
.A(n_1377),
.B(n_368),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1489),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1564),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1668),
.A2(n_370),
.B(n_369),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1545),
.B(n_1547),
.Y(n_1824)
);

NAND2x1p5_ASAP7_75t_L g1825 ( 
.A(n_1645),
.B(n_372),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1523),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1523),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1501),
.Y(n_1828)
);

INVx4_ASAP7_75t_L g1829 ( 
.A(n_1530),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1501),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1506),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1506),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1516),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1371),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1444),
.B(n_137),
.Y(n_1835)
);

XOR2xp5_ASAP7_75t_L g1836 ( 
.A(n_1405),
.B(n_373),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1379),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1566),
.B(n_137),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1395),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1458),
.B(n_138),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1469),
.Y(n_1841)
);

NOR2xp67_ASAP7_75t_L g1842 ( 
.A(n_1520),
.B(n_375),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1682),
.B(n_377),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1362),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1495),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1417),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1495),
.Y(n_1847)
);

NAND2xp33_ASAP7_75t_R g1848 ( 
.A(n_1374),
.B(n_139),
.Y(n_1848)
);

XNOR2xp5_ASAP7_75t_L g1849 ( 
.A(n_1347),
.B(n_139),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1567),
.B(n_140),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1391),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1634),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1530),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1568),
.B(n_140),
.Y(n_1854)
);

XOR2xp5_ASAP7_75t_L g1855 ( 
.A(n_1405),
.B(n_378),
.Y(n_1855)
);

AO21x1_ASAP7_75t_L g1856 ( 
.A1(n_1576),
.A2(n_141),
.B(n_142),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1457),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1533),
.Y(n_1858)
);

INVx8_ASAP7_75t_L g1859 ( 
.A(n_1388),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1369),
.Y(n_1860)
);

NOR2xp67_ASAP7_75t_L g1861 ( 
.A(n_1514),
.B(n_386),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1369),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1362),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1531),
.Y(n_1864)
);

XOR2xp5_ASAP7_75t_L g1865 ( 
.A(n_1484),
.B(n_387),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1577),
.B(n_141),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1531),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1532),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1463),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1446),
.A2(n_390),
.B(n_388),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1532),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1509),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1608),
.B(n_391),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1509),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1472),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1549),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1612),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1616),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1485),
.Y(n_1879)
);

CKINVDCx16_ASAP7_75t_R g1880 ( 
.A(n_1490),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1621),
.B(n_142),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1617),
.Y(n_1882)
);

INVxp33_ASAP7_75t_L g1883 ( 
.A(n_1465),
.Y(n_1883)
);

NOR2xp67_ASAP7_75t_L g1884 ( 
.A(n_1517),
.B(n_393),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1619),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1578),
.B(n_144),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1639),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1485),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1404),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1503),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1477),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1500),
.Y(n_1892)
);

XOR2x2_ASAP7_75t_L g1893 ( 
.A(n_1427),
.B(n_144),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1591),
.B(n_145),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1526),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1580),
.B(n_146),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1539),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1492),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1527),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1491),
.B(n_146),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1499),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1477),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1546),
.B(n_147),
.Y(n_1903)
);

INVxp33_ASAP7_75t_L g1904 ( 
.A(n_1482),
.Y(n_1904)
);

INVx4_ASAP7_75t_L g1905 ( 
.A(n_1541),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1518),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_1466),
.Y(n_1907)
);

CKINVDCx16_ASAP7_75t_R g1908 ( 
.A(n_1613),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1356),
.Y(n_1909)
);

CKINVDCx20_ASAP7_75t_R g1910 ( 
.A(n_1642),
.Y(n_1910)
);

INVx8_ASAP7_75t_L g1911 ( 
.A(n_1388),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1356),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1658),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1515),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1651),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1553),
.Y(n_1916)
);

BUFx2_ASAP7_75t_L g1917 ( 
.A(n_1420),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1555),
.Y(n_1918)
);

XOR2xp5_ASAP7_75t_L g1919 ( 
.A(n_1478),
.B(n_394),
.Y(n_1919)
);

NOR2xp67_ASAP7_75t_L g1920 ( 
.A(n_1557),
.B(n_396),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1661),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1676),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1372),
.Y(n_1923)
);

INVx2_ASAP7_75t_SL g1924 ( 
.A(n_1632),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1654),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1554),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1569),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1401),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1504),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1636),
.B(n_147),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1508),
.B(n_397),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1378),
.B(n_148),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1521),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1525),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1537),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1563),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1519),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1556),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1570),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1584),
.Y(n_1940)
);

XOR2xp5_ASAP7_75t_L g1941 ( 
.A(n_1559),
.B(n_398),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1586),
.Y(n_1942)
);

XOR2xp5_ASAP7_75t_L g1943 ( 
.A(n_1560),
.B(n_399),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1590),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1594),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1497),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1667),
.Y(n_1947)
);

XOR2xp5_ASAP7_75t_L g1948 ( 
.A(n_1565),
.B(n_401),
.Y(n_1948)
);

XNOR2x2_ASAP7_75t_L g1949 ( 
.A(n_1606),
.B(n_148),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1583),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1389),
.B(n_1390),
.Y(n_1951)
);

XNOR2xp5_ASAP7_75t_L g1952 ( 
.A(n_1353),
.B(n_149),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1420),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1604),
.B(n_150),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1475),
.B(n_403),
.Y(n_1955)
);

INVx8_ASAP7_75t_L g1956 ( 
.A(n_1615),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1596),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1596),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1441),
.B(n_404),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1512),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1606),
.Y(n_1961)
);

CKINVDCx20_ASAP7_75t_R g1962 ( 
.A(n_1572),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1611),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1540),
.Y(n_1964)
);

XOR2xp5_ASAP7_75t_L g1965 ( 
.A(n_1582),
.B(n_405),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1623),
.B(n_150),
.Y(n_1966)
);

XOR2x2_ASAP7_75t_L g1967 ( 
.A(n_1597),
.B(n_151),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1611),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1627),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1415),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1627),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1400),
.B(n_152),
.Y(n_1972)
);

INVx2_ASAP7_75t_SL g1973 ( 
.A(n_1601),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1633),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1633),
.Y(n_1975)
);

INVxp67_ASAP7_75t_SL g1976 ( 
.A(n_1669),
.Y(n_1976)
);

NAND2xp33_ASAP7_75t_SL g1977 ( 
.A(n_1674),
.B(n_154),
.Y(n_1977)
);

INVxp33_ASAP7_75t_SL g1978 ( 
.A(n_1625),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1618),
.B(n_154),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1641),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1649),
.B(n_155),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1641),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1643),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1643),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1367),
.B(n_156),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1656),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1411),
.B(n_156),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1656),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1672),
.Y(n_1989)
);

XOR2xp5_ASAP7_75t_L g1990 ( 
.A(n_1628),
.B(n_406),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1675),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1679),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1629),
.B(n_157),
.Y(n_1993)
);

INVxp67_ASAP7_75t_L g1994 ( 
.A(n_1451),
.Y(n_1994)
);

INVxp67_ASAP7_75t_SL g1995 ( 
.A(n_1681),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1678),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1665),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1481),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1670),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1445),
.B(n_409),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1637),
.B(n_157),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1449),
.B(n_410),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1452),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1677),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1430),
.Y(n_2005)
);

OAI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1918),
.A2(n_1436),
.B(n_1431),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1746),
.B(n_1423),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1684),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1788),
.B(n_1424),
.Y(n_2009)
);

BUFx2_ASAP7_75t_L g2010 ( 
.A(n_1766),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1684),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1913),
.B(n_1438),
.Y(n_2012)
);

INVx2_ASAP7_75t_SL g2013 ( 
.A(n_1789),
.Y(n_2013)
);

INVx3_ASAP7_75t_L g2014 ( 
.A(n_1721),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1927),
.B(n_1640),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1778),
.B(n_1440),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1883),
.B(n_1453),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1794),
.B(n_1461),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1692),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1748),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1688),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1688),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1701),
.B(n_1380),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1758),
.Y(n_2024)
);

AND2x4_ASAP7_75t_L g2025 ( 
.A(n_1697),
.B(n_1839),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1685),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1947),
.B(n_1468),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1804),
.Y(n_2028)
);

BUFx5_ASAP7_75t_L g2029 ( 
.A(n_1687),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1755),
.B(n_1921),
.Y(n_2030)
);

INVxp33_ASAP7_75t_L g2031 ( 
.A(n_1689),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1749),
.B(n_1476),
.Y(n_2032)
);

INVx4_ASAP7_75t_L g2033 ( 
.A(n_1869),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1834),
.B(n_1673),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1694),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_1699),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1690),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1875),
.B(n_412),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1690),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1749),
.B(n_1479),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1762),
.Y(n_2041)
);

INVxp67_ASAP7_75t_L g2042 ( 
.A(n_1787),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_1813),
.B(n_1408),
.Y(n_2043)
);

INVx2_ASAP7_75t_SL g2044 ( 
.A(n_1821),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1694),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1824),
.B(n_1483),
.Y(n_2046)
);

AND2x2_ASAP7_75t_SL g2047 ( 
.A(n_1727),
.B(n_1385),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1696),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1851),
.B(n_1387),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1696),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1756),
.Y(n_2051)
);

INVxp67_ASAP7_75t_L g2052 ( 
.A(n_1848),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1857),
.B(n_1392),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1892),
.B(n_1895),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1757),
.Y(n_2055)
);

INVx2_ASAP7_75t_SL g2056 ( 
.A(n_1803),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1994),
.B(n_1409),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1859),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1759),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_1859),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_1762),
.Y(n_2061)
);

AND2x6_ASAP7_75t_L g2062 ( 
.A(n_1844),
.B(n_1631),
.Y(n_2062)
);

AND2x2_ASAP7_75t_SL g2063 ( 
.A(n_1908),
.B(n_1664),
.Y(n_2063)
);

BUFx3_ASAP7_75t_L g2064 ( 
.A(n_1762),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1760),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1763),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1869),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1764),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1773),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1858),
.B(n_1393),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1915),
.B(n_1402),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1776),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1806),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_1923),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1897),
.B(n_158),
.Y(n_2075)
);

OAI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1751),
.A2(n_1770),
.B(n_1738),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1877),
.B(n_158),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1716),
.B(n_1406),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1780),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1878),
.B(n_159),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_1929),
.B(n_1456),
.Y(n_2081)
);

BUFx3_ASAP7_75t_L g2082 ( 
.A(n_1911),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1781),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1784),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1775),
.B(n_1473),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1791),
.Y(n_2086)
);

BUFx3_ASAP7_75t_L g2087 ( 
.A(n_1911),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1792),
.Y(n_2088)
);

AND2x2_ASAP7_75t_SL g2089 ( 
.A(n_1880),
.B(n_1359),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1793),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1882),
.B(n_160),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1833),
.B(n_414),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1796),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1797),
.Y(n_2094)
);

INVx3_ASAP7_75t_L g2095 ( 
.A(n_1695),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1885),
.B(n_162),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1887),
.B(n_1904),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1801),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1802),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_1729),
.B(n_415),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1805),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1740),
.B(n_1459),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1809),
.Y(n_2103)
);

AND2x6_ASAP7_75t_L g2104 ( 
.A(n_1844),
.B(n_1480),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1691),
.B(n_1365),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1869),
.Y(n_2106)
);

INVxp67_ASAP7_75t_L g2107 ( 
.A(n_1736),
.Y(n_2107)
);

INVx4_ASAP7_75t_L g2108 ( 
.A(n_1687),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_1774),
.A2(n_417),
.B(n_416),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1810),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1691),
.B(n_418),
.Y(n_2111)
);

HB1xp67_ASAP7_75t_L g2112 ( 
.A(n_1938),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1811),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1812),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1702),
.B(n_163),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1818),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1814),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1815),
.Y(n_2118)
);

INVxp67_ASAP7_75t_L g2119 ( 
.A(n_1903),
.Y(n_2119)
);

OAI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_1843),
.A2(n_1769),
.B(n_1823),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_1907),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1700),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1939),
.B(n_419),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1841),
.B(n_164),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1698),
.Y(n_2125)
);

INVx4_ASAP7_75t_L g2126 ( 
.A(n_1687),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1940),
.B(n_422),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1890),
.B(n_165),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_1687),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1942),
.B(n_423),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1735),
.B(n_166),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1924),
.B(n_166),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1889),
.B(n_167),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1683),
.B(n_169),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1905),
.B(n_169),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_1750),
.B(n_427),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1945),
.B(n_428),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1863),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1946),
.B(n_429),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1860),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1822),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_1905),
.B(n_1932),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_1978),
.B(n_170),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1703),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1972),
.B(n_170),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1862),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1705),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1951),
.B(n_430),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1768),
.B(n_434),
.Y(n_2149)
);

INVx2_ASAP7_75t_SL g2150 ( 
.A(n_1956),
.Y(n_2150)
);

INVx1_ASAP7_75t_SL g2151 ( 
.A(n_1837),
.Y(n_2151)
);

BUFx3_ASAP7_75t_L g2152 ( 
.A(n_1826),
.Y(n_2152)
);

AND2x4_ASAP7_75t_L g2153 ( 
.A(n_1754),
.B(n_435),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1970),
.B(n_437),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1707),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_1987),
.B(n_171),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1708),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1761),
.B(n_171),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1709),
.Y(n_2159)
);

OAI21xp5_ASAP7_75t_L g2160 ( 
.A1(n_1876),
.A2(n_447),
.B(n_446),
.Y(n_2160)
);

INVx2_ASAP7_75t_SL g2161 ( 
.A(n_1956),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1828),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_1976),
.B(n_173),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1704),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1711),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_1966),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1786),
.B(n_450),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_SL g2168 ( 
.A(n_1852),
.B(n_174),
.Y(n_2168)
);

INVx2_ASAP7_75t_SL g2169 ( 
.A(n_1894),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_1928),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_1830),
.B(n_451),
.Y(n_2171)
);

INVx4_ASAP7_75t_L g2172 ( 
.A(n_1772),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_1827),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_1995),
.B(n_1930),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1998),
.B(n_174),
.Y(n_2175)
);

INVx1_ASAP7_75t_SL g2176 ( 
.A(n_1835),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1790),
.B(n_452),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1795),
.B(n_457),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_1973),
.A2(n_461),
.B1(n_462),
.B2(n_460),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_1816),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1714),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1807),
.B(n_175),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1906),
.B(n_464),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1838),
.B(n_1850),
.Y(n_2184)
);

OAI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_1873),
.A2(n_473),
.B(n_467),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1854),
.B(n_175),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1866),
.B(n_1914),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1715),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1717),
.Y(n_2189)
);

BUFx8_ASAP7_75t_L g2190 ( 
.A(n_1917),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_1845),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_1909),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1831),
.Y(n_2193)
);

INVxp67_ASAP7_75t_L g2194 ( 
.A(n_1993),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_1731),
.B(n_176),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1718),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1719),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_1777),
.Y(n_2198)
);

BUFx3_ASAP7_75t_L g2199 ( 
.A(n_1847),
.Y(n_2199)
);

BUFx2_ASAP7_75t_L g2200 ( 
.A(n_1846),
.Y(n_2200)
);

BUFx3_ASAP7_75t_L g2201 ( 
.A(n_1853),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2005),
.B(n_474),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1720),
.Y(n_2203)
);

AND2x2_ASAP7_75t_SL g2204 ( 
.A(n_1771),
.B(n_176),
.Y(n_2204)
);

INVxp67_ASAP7_75t_SL g2205 ( 
.A(n_1722),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_1916),
.B(n_177),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_1731),
.B(n_177),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_1891),
.B(n_178),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_1879),
.B(n_179),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_1832),
.B(n_476),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1898),
.B(n_478),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1723),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1926),
.B(n_480),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1912),
.B(n_485),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_1864),
.B(n_488),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_1922),
.B(n_180),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1724),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_R g2218 ( 
.A(n_1944),
.B(n_499),
.Y(n_2218)
);

INVx3_ASAP7_75t_L g2219 ( 
.A(n_1725),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_1925),
.B(n_180),
.Y(n_2220)
);

AND2x4_ASAP7_75t_SL g2221 ( 
.A(n_2003),
.B(n_504),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_1902),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_1950),
.B(n_181),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1840),
.B(n_181),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2001),
.B(n_186),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1996),
.B(n_186),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1686),
.B(n_505),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1726),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1920),
.B(n_506),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1728),
.Y(n_2230)
);

OAI21xp5_ASAP7_75t_L g2231 ( 
.A1(n_1870),
.A2(n_509),
.B(n_507),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1931),
.B(n_516),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1798),
.B(n_519),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1800),
.B(n_1808),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1730),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1881),
.B(n_520),
.Y(n_2236)
);

AND2x2_ASAP7_75t_SL g2237 ( 
.A(n_1900),
.B(n_187),
.Y(n_2237)
);

INVx1_ASAP7_75t_SL g2238 ( 
.A(n_1849),
.Y(n_2238)
);

BUFx3_ASAP7_75t_L g2239 ( 
.A(n_1817),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1732),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_1964),
.B(n_188),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_1996),
.B(n_189),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1997),
.B(n_189),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1997),
.B(n_190),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1710),
.B(n_523),
.Y(n_2245)
);

BUFx3_ASAP7_75t_L g2246 ( 
.A(n_1819),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1888),
.B(n_526),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1733),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_1867),
.Y(n_2249)
);

BUFx3_ASAP7_75t_L g2250 ( 
.A(n_1935),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1999),
.B(n_190),
.Y(n_2251)
);

NAND2x2_ASAP7_75t_L g2252 ( 
.A(n_2082),
.B(n_1953),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2174),
.B(n_1999),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_2026),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2107),
.B(n_1989),
.Y(n_2255)
);

INVx4_ASAP7_75t_L g2256 ( 
.A(n_2067),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_2041),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2184),
.B(n_1989),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2234),
.B(n_2030),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2187),
.B(n_1991),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2048),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2097),
.B(n_2004),
.Y(n_2262)
);

BUFx12f_ASAP7_75t_L g2263 ( 
.A(n_2058),
.Y(n_2263)
);

CKINVDCx20_ASAP7_75t_R g2264 ( 
.A(n_2198),
.Y(n_2264)
);

BUFx2_ASAP7_75t_L g2265 ( 
.A(n_2010),
.Y(n_2265)
);

CKINVDCx20_ASAP7_75t_R g2266 ( 
.A(n_2024),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_2087),
.B(n_1868),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_2013),
.B(n_2004),
.Y(n_2268)
);

BUFx4f_ASAP7_75t_L g2269 ( 
.A(n_2067),
.Y(n_2269)
);

HB1xp67_ASAP7_75t_L g2270 ( 
.A(n_2074),
.Y(n_2270)
);

INVx3_ASAP7_75t_L g2271 ( 
.A(n_2067),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_2033),
.B(n_1871),
.Y(n_2272)
);

BUFx12f_ASAP7_75t_L g2273 ( 
.A(n_2060),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_2194),
.B(n_1712),
.Y(n_2274)
);

INVx3_ASAP7_75t_L g2275 ( 
.A(n_2106),
.Y(n_2275)
);

NAND2x1p5_ASAP7_75t_L g2276 ( 
.A(n_2033),
.B(n_1899),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2016),
.B(n_1991),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2012),
.B(n_1992),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2106),
.B(n_1872),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_SL g2280 ( 
.A(n_2121),
.B(n_1910),
.Y(n_2280)
);

BUFx4f_ASAP7_75t_L g2281 ( 
.A(n_2106),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2008),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2015),
.B(n_1992),
.Y(n_2283)
);

INVx3_ASAP7_75t_L g2284 ( 
.A(n_2061),
.Y(n_2284)
);

NAND2x1p5_ASAP7_75t_L g2285 ( 
.A(n_2041),
.B(n_1899),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2054),
.B(n_1901),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2008),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_2064),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2011),
.Y(n_2289)
);

BUFx8_ASAP7_75t_L g2290 ( 
.A(n_2200),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2046),
.B(n_1874),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2042),
.B(n_2003),
.Y(n_2292)
);

AND2x4_ASAP7_75t_L g2293 ( 
.A(n_2025),
.B(n_1783),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_2119),
.B(n_1957),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2056),
.B(n_1958),
.Y(n_2295)
);

AND2x6_ASAP7_75t_L g2296 ( 
.A(n_2129),
.B(n_1986),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2052),
.B(n_1936),
.Y(n_2297)
);

INVx3_ASAP7_75t_L g2298 ( 
.A(n_2041),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2073),
.B(n_2019),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_2141),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2007),
.B(n_2036),
.Y(n_2301)
);

BUFx3_ASAP7_75t_L g2302 ( 
.A(n_2191),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2011),
.B(n_1986),
.Y(n_2303)
);

NAND2x1p5_ASAP7_75t_L g2304 ( 
.A(n_2108),
.B(n_1734),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2021),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2021),
.B(n_1988),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2022),
.B(n_1988),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_L g2308 ( 
.A(n_2166),
.B(n_1744),
.Y(n_2308)
);

AND2x2_ASAP7_75t_SL g2309 ( 
.A(n_2204),
.B(n_1886),
.Y(n_2309)
);

HB1xp67_ASAP7_75t_L g2310 ( 
.A(n_2222),
.Y(n_2310)
);

INVx4_ASAP7_75t_L g2311 ( 
.A(n_2250),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2022),
.Y(n_2312)
);

OR2x6_ASAP7_75t_L g2313 ( 
.A(n_2150),
.B(n_1752),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2035),
.Y(n_2314)
);

BUFx2_ASAP7_75t_L g2315 ( 
.A(n_2062),
.Y(n_2315)
);

INVxp67_ASAP7_75t_SL g2316 ( 
.A(n_2215),
.Y(n_2316)
);

BUFx5_ASAP7_75t_L g2317 ( 
.A(n_2035),
.Y(n_2317)
);

AND2x4_ASAP7_75t_L g2318 ( 
.A(n_2025),
.B(n_1937),
.Y(n_2318)
);

NOR2x1_ASAP7_75t_L g2319 ( 
.A(n_2148),
.B(n_1941),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2043),
.B(n_1961),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2009),
.B(n_1960),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_2218),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2045),
.Y(n_2323)
);

INVx8_ASAP7_75t_L g2324 ( 
.A(n_2104),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2045),
.B(n_1963),
.Y(n_2325)
);

BUFx3_ASAP7_75t_L g2326 ( 
.A(n_2199),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2050),
.B(n_1968),
.Y(n_2327)
);

INVx4_ASAP7_75t_L g2328 ( 
.A(n_2100),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2142),
.B(n_1975),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2050),
.B(n_1969),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2228),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2228),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2176),
.B(n_1980),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2027),
.B(n_1971),
.Y(n_2334)
);

INVx2_ASAP7_75t_SL g2335 ( 
.A(n_2044),
.Y(n_2335)
);

OR2x6_ASAP7_75t_L g2336 ( 
.A(n_2161),
.B(n_1752),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2017),
.B(n_1933),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_2057),
.B(n_1974),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2102),
.B(n_1982),
.Y(n_2339)
);

OR2x6_ASAP7_75t_L g2340 ( 
.A(n_2092),
.B(n_1799),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2248),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2170),
.B(n_1934),
.Y(n_2342)
);

NOR2xp67_ASAP7_75t_L g2343 ( 
.A(n_2169),
.B(n_1955),
.Y(n_2343)
);

BUFx2_ASAP7_75t_L g2344 ( 
.A(n_2062),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2248),
.Y(n_2345)
);

BUFx2_ASAP7_75t_L g2346 ( 
.A(n_2062),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_2062),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_2152),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2051),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2134),
.B(n_1983),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2051),
.Y(n_2351)
);

INVx1_ASAP7_75t_SL g2352 ( 
.A(n_2151),
.Y(n_2352)
);

INVxp67_ASAP7_75t_L g2353 ( 
.A(n_2192),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_2081),
.B(n_1984),
.Y(n_2354)
);

AND2x6_ASAP7_75t_L g2355 ( 
.A(n_2129),
.B(n_2003),
.Y(n_2355)
);

INVxp67_ASAP7_75t_L g2356 ( 
.A(n_2112),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_2173),
.Y(n_2357)
);

OR2x2_ASAP7_75t_L g2358 ( 
.A(n_2238),
.B(n_1949),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2215),
.B(n_2002),
.Y(n_2359)
);

AND2x4_ASAP7_75t_L g2360 ( 
.A(n_2038),
.B(n_2092),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2055),
.Y(n_2361)
);

INVx2_ASAP7_75t_SL g2362 ( 
.A(n_2132),
.Y(n_2362)
);

INVx4_ASAP7_75t_L g2363 ( 
.A(n_2100),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2055),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2068),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2068),
.Y(n_2366)
);

BUFx6f_ASAP7_75t_L g2367 ( 
.A(n_2180),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_2105),
.B(n_1977),
.Y(n_2368)
);

INVx4_ASAP7_75t_L g2369 ( 
.A(n_2136),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2138),
.B(n_2000),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_L g2371 ( 
.A(n_2032),
.B(n_1962),
.Y(n_2371)
);

NAND2x1p5_ASAP7_75t_L g2372 ( 
.A(n_2108),
.B(n_2126),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2138),
.B(n_1959),
.Y(n_2373)
);

AND2x4_ASAP7_75t_L g2374 ( 
.A(n_2038),
.B(n_1737),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_SL g2375 ( 
.A(n_2047),
.B(n_1799),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_2141),
.Y(n_2376)
);

INVx5_ASAP7_75t_L g2377 ( 
.A(n_2104),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2018),
.B(n_1985),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2069),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2145),
.B(n_1820),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2069),
.Y(n_2381)
);

CKINVDCx20_ASAP7_75t_R g2382 ( 
.A(n_2190),
.Y(n_2382)
);

OR2x6_ASAP7_75t_L g2383 ( 
.A(n_2171),
.B(n_1954),
.Y(n_2383)
);

BUFx3_ASAP7_75t_L g2384 ( 
.A(n_2190),
.Y(n_2384)
);

INVx4_ASAP7_75t_L g2385 ( 
.A(n_2136),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_SL g2386 ( 
.A(n_2143),
.B(n_1979),
.Y(n_2386)
);

BUFx10_ASAP7_75t_L g2387 ( 
.A(n_2241),
.Y(n_2387)
);

NAND2x1p5_ASAP7_75t_L g2388 ( 
.A(n_2126),
.B(n_1739),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2083),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2083),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2156),
.B(n_1765),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2084),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_SL g2393 ( 
.A(n_2237),
.B(n_1981),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2140),
.B(n_1779),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_2089),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2140),
.B(n_1782),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2163),
.B(n_1706),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2084),
.Y(n_2398)
);

INVx3_ASAP7_75t_L g2399 ( 
.A(n_2141),
.Y(n_2399)
);

AND2x4_ASAP7_75t_L g2400 ( 
.A(n_2201),
.B(n_2239),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_2171),
.B(n_1741),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2146),
.B(n_1785),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2086),
.Y(n_2403)
);

HB1xp67_ASAP7_75t_L g2404 ( 
.A(n_2249),
.Y(n_2404)
);

NAND2xp33_ASAP7_75t_L g2405 ( 
.A(n_2029),
.B(n_1825),
.Y(n_2405)
);

AND2x2_ASAP7_75t_SL g2406 ( 
.A(n_2063),
.B(n_1893),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2146),
.B(n_1896),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2182),
.B(n_2186),
.Y(n_2408)
);

INVx4_ASAP7_75t_L g2409 ( 
.A(n_2153),
.Y(n_2409)
);

INVx4_ASAP7_75t_L g2410 ( 
.A(n_2153),
.Y(n_2410)
);

BUFx3_ASAP7_75t_L g2411 ( 
.A(n_2246),
.Y(n_2411)
);

BUFx12f_ASAP7_75t_L g2412 ( 
.A(n_2290),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2287),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2259),
.B(n_2071),
.Y(n_2414)
);

BUFx3_ASAP7_75t_L g2415 ( 
.A(n_2266),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2289),
.Y(n_2416)
);

BUFx12f_ASAP7_75t_L g2417 ( 
.A(n_2263),
.Y(n_2417)
);

CKINVDCx20_ASAP7_75t_R g2418 ( 
.A(n_2264),
.Y(n_2418)
);

BUFx6f_ASAP7_75t_L g2419 ( 
.A(n_2348),
.Y(n_2419)
);

BUFx12f_ASAP7_75t_L g2420 ( 
.A(n_2273),
.Y(n_2420)
);

BUFx6f_ASAP7_75t_L g2421 ( 
.A(n_2348),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2305),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2312),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2314),
.Y(n_2424)
);

HB1xp67_ASAP7_75t_L g2425 ( 
.A(n_2265),
.Y(n_2425)
);

INVx4_ASAP7_75t_L g2426 ( 
.A(n_2367),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_2367),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2323),
.Y(n_2428)
);

OR2x6_ASAP7_75t_L g2429 ( 
.A(n_2265),
.B(n_2210),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_2254),
.Y(n_2430)
);

BUFx2_ASAP7_75t_SL g2431 ( 
.A(n_2256),
.Y(n_2431)
);

INVx3_ASAP7_75t_SL g2432 ( 
.A(n_2352),
.Y(n_2432)
);

BUFx3_ASAP7_75t_L g2433 ( 
.A(n_2357),
.Y(n_2433)
);

INVxp67_ASAP7_75t_SL g2434 ( 
.A(n_2316),
.Y(n_2434)
);

BUFx12f_ASAP7_75t_L g2435 ( 
.A(n_2357),
.Y(n_2435)
);

INVxp67_ASAP7_75t_SL g2436 ( 
.A(n_2317),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2278),
.B(n_2225),
.Y(n_2437)
);

BUFx3_ASAP7_75t_L g2438 ( 
.A(n_2302),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2282),
.Y(n_2439)
);

NAND2x1p5_ASAP7_75t_L g2440 ( 
.A(n_2269),
.B(n_2172),
.Y(n_2440)
);

INVx5_ASAP7_75t_L g2441 ( 
.A(n_2257),
.Y(n_2441)
);

BUFx2_ASAP7_75t_L g2442 ( 
.A(n_2279),
.Y(n_2442)
);

INVx5_ASAP7_75t_L g2443 ( 
.A(n_2257),
.Y(n_2443)
);

AND2x4_ASAP7_75t_L g2444 ( 
.A(n_2311),
.B(n_2180),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_2326),
.Y(n_2445)
);

AOI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2386),
.A2(n_2393),
.B1(n_2371),
.B2(n_2360),
.Y(n_2446)
);

AOI22xp5_ASAP7_75t_L g2447 ( 
.A1(n_2360),
.A2(n_2236),
.B1(n_2233),
.B2(n_2023),
.Y(n_2447)
);

BUFx2_ASAP7_75t_SL g2448 ( 
.A(n_2317),
.Y(n_2448)
);

CKINVDCx11_ASAP7_75t_R g2449 ( 
.A(n_2382),
.Y(n_2449)
);

BUFx2_ASAP7_75t_L g2450 ( 
.A(n_2279),
.Y(n_2450)
);

INVx2_ASAP7_75t_SL g2451 ( 
.A(n_2335),
.Y(n_2451)
);

BUFx2_ASAP7_75t_SL g2452 ( 
.A(n_2317),
.Y(n_2452)
);

AND2x4_ASAP7_75t_L g2453 ( 
.A(n_2318),
.B(n_2180),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_2281),
.Y(n_2454)
);

BUFx12f_ASAP7_75t_L g2455 ( 
.A(n_2384),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2277),
.B(n_2040),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2408),
.B(n_2175),
.Y(n_2457)
);

BUFx4_ASAP7_75t_SL g2458 ( 
.A(n_2340),
.Y(n_2458)
);

INVx2_ASAP7_75t_SL g2459 ( 
.A(n_2268),
.Y(n_2459)
);

INVx2_ASAP7_75t_SL g2460 ( 
.A(n_2333),
.Y(n_2460)
);

BUFx3_ASAP7_75t_L g2461 ( 
.A(n_2411),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2351),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2331),
.Y(n_2463)
);

INVx1_ASAP7_75t_SL g2464 ( 
.A(n_2297),
.Y(n_2464)
);

INVx6_ASAP7_75t_L g2465 ( 
.A(n_2252),
.Y(n_2465)
);

BUFx5_ASAP7_75t_L g2466 ( 
.A(n_2355),
.Y(n_2466)
);

BUFx12f_ASAP7_75t_L g2467 ( 
.A(n_2313),
.Y(n_2467)
);

INVx3_ASAP7_75t_L g2468 ( 
.A(n_2400),
.Y(n_2468)
);

BUFx2_ASAP7_75t_SL g2469 ( 
.A(n_2284),
.Y(n_2469)
);

INVx1_ASAP7_75t_SL g2470 ( 
.A(n_2286),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2332),
.Y(n_2471)
);

CKINVDCx16_ASAP7_75t_R g2472 ( 
.A(n_2280),
.Y(n_2472)
);

INVxp67_ASAP7_75t_SL g2473 ( 
.A(n_2317),
.Y(n_2473)
);

AOI22xp33_ASAP7_75t_L g2474 ( 
.A1(n_2309),
.A2(n_2104),
.B1(n_2231),
.B2(n_2206),
.Y(n_2474)
);

BUFx4f_ASAP7_75t_SL g2475 ( 
.A(n_2294),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2337),
.B(n_2034),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_L g2477 ( 
.A(n_2308),
.B(n_2031),
.Y(n_2477)
);

BUFx2_ASAP7_75t_L g2478 ( 
.A(n_2318),
.Y(n_2478)
);

NAND2x1p5_ASAP7_75t_L g2479 ( 
.A(n_2328),
.B(n_2172),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2361),
.Y(n_2480)
);

OAI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2359),
.A2(n_2363),
.B1(n_2385),
.B2(n_2369),
.Y(n_2481)
);

INVx4_ASAP7_75t_L g2482 ( 
.A(n_2288),
.Y(n_2482)
);

BUFx6f_ASAP7_75t_L g2483 ( 
.A(n_2267),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2364),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2341),
.Y(n_2485)
);

INVxp67_ASAP7_75t_SL g2486 ( 
.A(n_2310),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2345),
.Y(n_2487)
);

INVx1_ASAP7_75t_SL g2488 ( 
.A(n_2262),
.Y(n_2488)
);

BUFx2_ASAP7_75t_L g2489 ( 
.A(n_2301),
.Y(n_2489)
);

BUFx12f_ASAP7_75t_L g2490 ( 
.A(n_2313),
.Y(n_2490)
);

BUFx2_ASAP7_75t_L g2491 ( 
.A(n_2293),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2349),
.Y(n_2492)
);

BUFx6f_ASAP7_75t_L g2493 ( 
.A(n_2401),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2366),
.Y(n_2494)
);

BUFx10_ASAP7_75t_L g2495 ( 
.A(n_2274),
.Y(n_2495)
);

CKINVDCx20_ASAP7_75t_R g2496 ( 
.A(n_2322),
.Y(n_2496)
);

BUFx12f_ASAP7_75t_L g2497 ( 
.A(n_2336),
.Y(n_2497)
);

BUFx2_ASAP7_75t_SL g2498 ( 
.A(n_2404),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2381),
.Y(n_2499)
);

BUFx3_ASAP7_75t_L g2500 ( 
.A(n_2270),
.Y(n_2500)
);

OAI22xp33_ASAP7_75t_SL g2501 ( 
.A1(n_2375),
.A2(n_2168),
.B1(n_2223),
.B2(n_2085),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2260),
.B(n_2226),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2365),
.Y(n_2503)
);

HB1xp67_ASAP7_75t_L g2504 ( 
.A(n_2353),
.Y(n_2504)
);

INVx3_ASAP7_75t_L g2505 ( 
.A(n_2300),
.Y(n_2505)
);

INVx5_ASAP7_75t_L g2506 ( 
.A(n_2296),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2376),
.Y(n_2507)
);

INVx2_ASAP7_75t_SL g2508 ( 
.A(n_2342),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_L g2509 ( 
.A(n_2401),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2293),
.Y(n_2510)
);

BUFx6f_ASAP7_75t_L g2511 ( 
.A(n_2272),
.Y(n_2511)
);

BUFx6f_ASAP7_75t_L g2512 ( 
.A(n_2324),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2463),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2471),
.Y(n_2514)
);

OAI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2474),
.A2(n_2409),
.B1(n_2410),
.B2(n_2320),
.Y(n_2515)
);

CKINVDCx11_ASAP7_75t_R g2516 ( 
.A(n_2412),
.Y(n_2516)
);

OAI22xp5_ASAP7_75t_L g2517 ( 
.A1(n_2502),
.A2(n_2383),
.B1(n_2338),
.B2(n_2368),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2485),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2487),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2492),
.Y(n_2520)
);

INVx1_ASAP7_75t_SL g2521 ( 
.A(n_2432),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_2435),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2494),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2499),
.Y(n_2524)
);

OAI22xp33_ASAP7_75t_L g2525 ( 
.A1(n_2472),
.A2(n_2395),
.B1(n_2283),
.B2(n_2368),
.Y(n_2525)
);

OAI22xp5_ASAP7_75t_SL g2526 ( 
.A1(n_2475),
.A2(n_2406),
.B1(n_1865),
.B2(n_1919),
.Y(n_2526)
);

INVx6_ASAP7_75t_L g2527 ( 
.A(n_2454),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2439),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2413),
.Y(n_2529)
);

INVx5_ASAP7_75t_L g2530 ( 
.A(n_2454),
.Y(n_2530)
);

AOI22xp33_ASAP7_75t_SL g2531 ( 
.A1(n_2501),
.A2(n_2380),
.B1(n_2391),
.B2(n_2397),
.Y(n_2531)
);

INVx2_ASAP7_75t_SL g2532 ( 
.A(n_2419),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2416),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2423),
.Y(n_2534)
);

BUFx12f_ASAP7_75t_L g2535 ( 
.A(n_2449),
.Y(n_2535)
);

INVx4_ASAP7_75t_L g2536 ( 
.A(n_2441),
.Y(n_2536)
);

BUFx2_ASAP7_75t_SL g2537 ( 
.A(n_2418),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2428),
.Y(n_2538)
);

OAI22xp5_ASAP7_75t_L g2539 ( 
.A1(n_2437),
.A2(n_2383),
.B1(n_2354),
.B2(n_2334),
.Y(n_2539)
);

AOI22xp33_ASAP7_75t_L g2540 ( 
.A1(n_2476),
.A2(n_2319),
.B1(n_2378),
.B2(n_1713),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_SL g2541 ( 
.A1(n_2489),
.A2(n_2387),
.B1(n_2221),
.B2(n_2243),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2456),
.B(n_2253),
.Y(n_2542)
);

BUFx6f_ASAP7_75t_L g2543 ( 
.A(n_2441),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_2438),
.Y(n_2544)
);

INVx4_ASAP7_75t_L g2545 ( 
.A(n_2441),
.Y(n_2545)
);

AOI22xp33_ASAP7_75t_L g2546 ( 
.A1(n_2489),
.A2(n_2321),
.B1(n_2104),
.B2(n_1943),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_2478),
.A2(n_1948),
.B1(n_1990),
.B2(n_1965),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2422),
.Y(n_2548)
);

INVx8_ASAP7_75t_L g2549 ( 
.A(n_2443),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2424),
.Y(n_2550)
);

OAI22x1_ASAP7_75t_SL g2551 ( 
.A1(n_2430),
.A2(n_1693),
.B1(n_1967),
.B2(n_1952),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2462),
.Y(n_2552)
);

AOI22xp33_ASAP7_75t_L g2553 ( 
.A1(n_2478),
.A2(n_2006),
.B1(n_2291),
.B2(n_2292),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2480),
.Y(n_2554)
);

AOI22xp33_ASAP7_75t_SL g2555 ( 
.A1(n_2488),
.A2(n_2244),
.B1(n_2251),
.B2(n_2242),
.Y(n_2555)
);

CKINVDCx11_ASAP7_75t_R g2556 ( 
.A(n_2417),
.Y(n_2556)
);

BUFx8_ASAP7_75t_L g2557 ( 
.A(n_2420),
.Y(n_2557)
);

BUFx3_ASAP7_75t_L g2558 ( 
.A(n_2419),
.Y(n_2558)
);

INVx4_ASAP7_75t_L g2559 ( 
.A(n_2443),
.Y(n_2559)
);

AOI22xp33_ASAP7_75t_L g2560 ( 
.A1(n_2508),
.A2(n_2329),
.B1(n_2324),
.B2(n_2220),
.Y(n_2560)
);

AOI22xp33_ASAP7_75t_L g2561 ( 
.A1(n_2491),
.A2(n_2510),
.B1(n_2470),
.B2(n_2459),
.Y(n_2561)
);

CKINVDCx20_ASAP7_75t_R g2562 ( 
.A(n_2496),
.Y(n_2562)
);

CKINVDCx20_ASAP7_75t_R g2563 ( 
.A(n_2415),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_2495),
.Y(n_2564)
);

BUFx12f_ASAP7_75t_L g2565 ( 
.A(n_2455),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2484),
.Y(n_2566)
);

AOI22xp33_ASAP7_75t_L g2567 ( 
.A1(n_2491),
.A2(n_2227),
.B1(n_2224),
.B2(n_2377),
.Y(n_2567)
);

CKINVDCx20_ASAP7_75t_R g2568 ( 
.A(n_2445),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2503),
.Y(n_2569)
);

CKINVDCx14_ASAP7_75t_R g2570 ( 
.A(n_2461),
.Y(n_2570)
);

AOI22xp33_ASAP7_75t_L g2571 ( 
.A1(n_2510),
.A2(n_2377),
.B1(n_2115),
.B2(n_2339),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2460),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2442),
.Y(n_2573)
);

CKINVDCx16_ASAP7_75t_R g2574 ( 
.A(n_2433),
.Y(n_2574)
);

CKINVDCx11_ASAP7_75t_R g2575 ( 
.A(n_2467),
.Y(n_2575)
);

AOI22xp33_ASAP7_75t_L g2576 ( 
.A1(n_2464),
.A2(n_2414),
.B1(n_2450),
.B2(n_2442),
.Y(n_2576)
);

CKINVDCx6p67_ASAP7_75t_R g2577 ( 
.A(n_2443),
.Y(n_2577)
);

BUFx6f_ASAP7_75t_L g2578 ( 
.A(n_2421),
.Y(n_2578)
);

BUFx2_ASAP7_75t_SL g2579 ( 
.A(n_2421),
.Y(n_2579)
);

BUFx2_ASAP7_75t_L g2580 ( 
.A(n_2425),
.Y(n_2580)
);

OAI21xp33_ASAP7_75t_L g2581 ( 
.A1(n_2457),
.A2(n_2255),
.B(n_2258),
.Y(n_2581)
);

BUFx12f_ASAP7_75t_L g2582 ( 
.A(n_2490),
.Y(n_2582)
);

INVx6_ASAP7_75t_L g2583 ( 
.A(n_2483),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2450),
.B(n_2358),
.Y(n_2584)
);

AOI22xp33_ASAP7_75t_L g2585 ( 
.A1(n_2446),
.A2(n_2377),
.B1(n_2131),
.B2(n_2210),
.Y(n_2585)
);

INVx3_ASAP7_75t_SL g2586 ( 
.A(n_2465),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2434),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_2458),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2505),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2453),
.B(n_2358),
.Y(n_2590)
);

OAI22xp33_ASAP7_75t_L g2591 ( 
.A1(n_2429),
.A2(n_2356),
.B1(n_2340),
.B2(n_2362),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2444),
.Y(n_2592)
);

CKINVDCx20_ASAP7_75t_R g2593 ( 
.A(n_2500),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2584),
.B(n_2429),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2529),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2566),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2580),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2542),
.B(n_2477),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2513),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2514),
.Y(n_2600)
);

INVx4_ASAP7_75t_L g2601 ( 
.A(n_2549),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2530),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2525),
.B(n_2504),
.Y(n_2603)
);

AOI22xp33_ASAP7_75t_L g2604 ( 
.A1(n_2531),
.A2(n_2160),
.B1(n_2135),
.B2(n_2154),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2590),
.B(n_2216),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2540),
.B(n_2299),
.Y(n_2606)
);

AOI22xp33_ASAP7_75t_SL g2607 ( 
.A1(n_2526),
.A2(n_2120),
.B1(n_2207),
.B2(n_2195),
.Y(n_2607)
);

OAI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2541),
.A2(n_2447),
.B1(n_2486),
.B2(n_2343),
.Y(n_2608)
);

AOI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2555),
.A2(n_2213),
.B1(n_2053),
.B2(n_2070),
.Y(n_2609)
);

INVx3_ASAP7_75t_L g2610 ( 
.A(n_2536),
.Y(n_2610)
);

AOI22xp33_ASAP7_75t_L g2611 ( 
.A1(n_2546),
.A2(n_2049),
.B1(n_2183),
.B2(n_2149),
.Y(n_2611)
);

OAI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_2553),
.A2(n_2294),
.B1(n_2452),
.B2(n_2448),
.Y(n_2612)
);

AOI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_2517),
.A2(n_2581),
.B1(n_2585),
.B2(n_2539),
.Y(n_2613)
);

INVx3_ASAP7_75t_SL g2614 ( 
.A(n_2588),
.Y(n_2614)
);

INVxp67_ASAP7_75t_SL g2615 ( 
.A(n_2587),
.Y(n_2615)
);

AOI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2547),
.A2(n_2481),
.B1(n_2374),
.B2(n_2468),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2518),
.Y(n_2617)
);

AOI22xp5_ASAP7_75t_L g2618 ( 
.A1(n_2515),
.A2(n_2374),
.B1(n_1855),
.B2(n_1836),
.Y(n_2618)
);

AOI22xp33_ASAP7_75t_L g2619 ( 
.A1(n_2571),
.A2(n_2185),
.B1(n_2139),
.B2(n_2124),
.Y(n_2619)
);

OR2x2_ASAP7_75t_L g2620 ( 
.A(n_2576),
.B(n_2498),
.Y(n_2620)
);

AOI22xp33_ASAP7_75t_L g2621 ( 
.A1(n_2560),
.A2(n_2202),
.B1(n_2078),
.B2(n_2127),
.Y(n_2621)
);

CKINVDCx5p33_ASAP7_75t_R g2622 ( 
.A(n_2562),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_L g2623 ( 
.A1(n_2567),
.A2(n_2130),
.B1(n_2137),
.B2(n_2123),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2561),
.B(n_2370),
.Y(n_2624)
);

BUFx3_ASAP7_75t_L g2625 ( 
.A(n_2530),
.Y(n_2625)
);

OAI22xp5_ASAP7_75t_SL g2626 ( 
.A1(n_2593),
.A2(n_1767),
.B1(n_2336),
.B2(n_2497),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2551),
.B(n_2482),
.Y(n_2627)
);

AOI22xp33_ASAP7_75t_L g2628 ( 
.A1(n_2591),
.A2(n_2077),
.B1(n_2091),
.B2(n_2080),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2519),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2573),
.A2(n_2096),
.B1(n_2128),
.B2(n_2211),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2520),
.Y(n_2631)
);

OAI22xp5_ASAP7_75t_SL g2632 ( 
.A1(n_2564),
.A2(n_2493),
.B1(n_2509),
.B2(n_2350),
.Y(n_2632)
);

AOI22xp33_ASAP7_75t_L g2633 ( 
.A1(n_2537),
.A2(n_2075),
.B1(n_1842),
.B2(n_1884),
.Y(n_2633)
);

AOI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2572),
.A2(n_1861),
.B1(n_1856),
.B2(n_2373),
.Y(n_2634)
);

AOI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2521),
.A2(n_2509),
.B1(n_2493),
.B2(n_2315),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2523),
.Y(n_2636)
);

OAI21xp5_ASAP7_75t_L g2637 ( 
.A1(n_2548),
.A2(n_2076),
.B(n_2232),
.Y(n_2637)
);

AOI22xp33_ASAP7_75t_SL g2638 ( 
.A1(n_2549),
.A2(n_2452),
.B1(n_2448),
.B2(n_2315),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2592),
.B(n_2379),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_SL g2640 ( 
.A1(n_2535),
.A2(n_2344),
.B1(n_2347),
.B2(n_2346),
.Y(n_2640)
);

OAI21xp5_ASAP7_75t_SL g2641 ( 
.A1(n_2570),
.A2(n_1742),
.B(n_2179),
.Y(n_2641)
);

OAI22xp5_ASAP7_75t_L g2642 ( 
.A1(n_2533),
.A2(n_2346),
.B1(n_2347),
.B2(n_2344),
.Y(n_2642)
);

AOI22xp33_ASAP7_75t_L g2643 ( 
.A1(n_2550),
.A2(n_2389),
.B1(n_2390),
.B2(n_2133),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2552),
.B(n_2407),
.Y(n_2644)
);

AOI22xp33_ASAP7_75t_L g2645 ( 
.A1(n_2554),
.A2(n_2261),
.B1(n_2219),
.B2(n_2177),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2524),
.Y(n_2646)
);

OAI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2528),
.A2(n_2398),
.B1(n_2403),
.B2(n_2392),
.Y(n_2647)
);

OAI21xp33_ASAP7_75t_L g2648 ( 
.A1(n_2534),
.A2(n_2396),
.B(n_2394),
.Y(n_2648)
);

AOI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2569),
.A2(n_2219),
.B1(n_2178),
.B2(n_2167),
.Y(n_2649)
);

BUFx12f_ASAP7_75t_L g2650 ( 
.A(n_2516),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2538),
.B(n_2451),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2589),
.Y(n_2652)
);

OAI222xp33_ASAP7_75t_L g2653 ( 
.A1(n_2563),
.A2(n_2214),
.B1(n_2247),
.B2(n_2402),
.C1(n_2276),
.C2(n_2330),
.Y(n_2653)
);

INVx3_ASAP7_75t_L g2654 ( 
.A(n_2536),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_L g2655 ( 
.A(n_2574),
.B(n_2511),
.Y(n_2655)
);

INVx4_ASAP7_75t_L g2656 ( 
.A(n_2530),
.Y(n_2656)
);

NOR2x1_ASAP7_75t_SL g2657 ( 
.A(n_2545),
.B(n_2431),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2543),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2543),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2543),
.Y(n_2660)
);

OAI21xp33_ASAP7_75t_L g2661 ( 
.A1(n_2544),
.A2(n_2098),
.B(n_2086),
.Y(n_2661)
);

BUFx4f_ASAP7_75t_SL g2662 ( 
.A(n_2568),
.Y(n_2662)
);

BUFx2_ASAP7_75t_L g2663 ( 
.A(n_2558),
.Y(n_2663)
);

OAI21xp5_ASAP7_75t_SL g2664 ( 
.A1(n_2532),
.A2(n_2111),
.B(n_2208),
.Y(n_2664)
);

AOI22xp33_ASAP7_75t_SL g2665 ( 
.A1(n_2582),
.A2(n_2029),
.B1(n_2469),
.B2(n_2405),
.Y(n_2665)
);

AOI22xp33_ASAP7_75t_L g2666 ( 
.A1(n_2575),
.A2(n_2099),
.B1(n_2101),
.B2(n_2098),
.Y(n_2666)
);

AOI22xp33_ASAP7_75t_L g2667 ( 
.A1(n_2522),
.A2(n_2101),
.B1(n_2103),
.B2(n_2099),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2583),
.A2(n_2110),
.B1(n_2114),
.B2(n_2103),
.Y(n_2668)
);

OAI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2577),
.A2(n_2306),
.B1(n_2307),
.B2(n_2303),
.Y(n_2669)
);

AOI22xp33_ASAP7_75t_L g2670 ( 
.A1(n_2607),
.A2(n_2114),
.B1(n_2110),
.B2(n_2229),
.Y(n_2670)
);

AOI22xp33_ASAP7_75t_SL g2671 ( 
.A1(n_2606),
.A2(n_2557),
.B1(n_2029),
.B2(n_2565),
.Y(n_2671)
);

AOI22xp33_ASAP7_75t_L g2672 ( 
.A1(n_2613),
.A2(n_2165),
.B1(n_2181),
.B2(n_2164),
.Y(n_2672)
);

OAI22xp5_ASAP7_75t_L g2673 ( 
.A1(n_2598),
.A2(n_2325),
.B1(n_2327),
.B2(n_2436),
.Y(n_2673)
);

NAND3xp33_ASAP7_75t_L g2674 ( 
.A(n_2611),
.B(n_2155),
.C(n_2147),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_SL g2675 ( 
.A1(n_2608),
.A2(n_2557),
.B1(n_2029),
.B2(n_2545),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2599),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2629),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2600),
.Y(n_2678)
);

OAI222xp33_ASAP7_75t_L g2679 ( 
.A1(n_2618),
.A2(n_2285),
.B1(n_2295),
.B2(n_2147),
.C1(n_2157),
.C2(n_2155),
.Y(n_2679)
);

BUFx2_ASAP7_75t_SL g2680 ( 
.A(n_2625),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2615),
.B(n_2473),
.Y(n_2681)
);

OAI221xp5_ASAP7_75t_SL g2682 ( 
.A1(n_2641),
.A2(n_2209),
.B1(n_2193),
.B2(n_2162),
.C(n_2188),
.Y(n_2682)
);

AOI22xp33_ASAP7_75t_L g2683 ( 
.A1(n_2604),
.A2(n_2603),
.B1(n_2609),
.B2(n_2619),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_L g2684 ( 
.A1(n_2648),
.A2(n_2196),
.B1(n_2197),
.B2(n_2189),
.Y(n_2684)
);

INVx3_ASAP7_75t_L g2685 ( 
.A(n_2610),
.Y(n_2685)
);

AOI22xp33_ASAP7_75t_L g2686 ( 
.A1(n_2605),
.A2(n_2212),
.B1(n_2217),
.B2(n_2203),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2594),
.B(n_2158),
.Y(n_2687)
);

AOI22xp33_ASAP7_75t_L g2688 ( 
.A1(n_2621),
.A2(n_2235),
.B1(n_2240),
.B2(n_2230),
.Y(n_2688)
);

OAI222xp33_ASAP7_75t_L g2689 ( 
.A1(n_2628),
.A2(n_2157),
.B1(n_2159),
.B2(n_2440),
.C1(n_2205),
.C2(n_2162),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_2620),
.A2(n_2669),
.B1(n_2624),
.B2(n_2630),
.Y(n_2690)
);

AND2x4_ASAP7_75t_SL g2691 ( 
.A(n_2656),
.B(n_2559),
.Y(n_2691)
);

AOI22xp33_ASAP7_75t_L g2692 ( 
.A1(n_2669),
.A2(n_2159),
.B1(n_2144),
.B2(n_2125),
.Y(n_2692)
);

OAI222xp33_ASAP7_75t_L g2693 ( 
.A1(n_2640),
.A2(n_2193),
.B1(n_2479),
.B2(n_2399),
.C1(n_2506),
.C2(n_2271),
.Y(n_2693)
);

AOI22xp33_ASAP7_75t_L g2694 ( 
.A1(n_2632),
.A2(n_2355),
.B1(n_2059),
.B2(n_2066),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2595),
.B(n_2427),
.Y(n_2695)
);

OA21x2_ASAP7_75t_L g2696 ( 
.A1(n_2637),
.A2(n_2109),
.B(n_2245),
.Y(n_2696)
);

OAI22xp5_ASAP7_75t_SL g2697 ( 
.A1(n_2626),
.A2(n_2527),
.B1(n_2586),
.B2(n_2583),
.Y(n_2697)
);

AOI22xp33_ASAP7_75t_SL g2698 ( 
.A1(n_2612),
.A2(n_2029),
.B1(n_2506),
.B2(n_2431),
.Y(n_2698)
);

OAI221xp5_ASAP7_75t_L g2699 ( 
.A1(n_2641),
.A2(n_2117),
.B1(n_2065),
.B2(n_2072),
.C(n_2079),
.Y(n_2699)
);

AOI22xp33_ASAP7_75t_L g2700 ( 
.A1(n_2633),
.A2(n_2355),
.B1(n_2090),
.B2(n_2093),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2612),
.B(n_2275),
.Y(n_2701)
);

OA21x2_ASAP7_75t_L g2702 ( 
.A1(n_2637),
.A2(n_1745),
.B(n_1743),
.Y(n_2702)
);

AOI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2616),
.A2(n_2556),
.B1(n_2511),
.B2(n_2483),
.Y(n_2703)
);

AOI22xp33_ASAP7_75t_L g2704 ( 
.A1(n_2623),
.A2(n_2094),
.B1(n_2113),
.B2(n_2088),
.Y(n_2704)
);

AOI22xp33_ASAP7_75t_L g2705 ( 
.A1(n_2661),
.A2(n_2118),
.B1(n_1753),
.B2(n_1747),
.Y(n_2705)
);

OAI221xp5_ASAP7_75t_SL g2706 ( 
.A1(n_2664),
.A2(n_2116),
.B1(n_2507),
.B2(n_2122),
.C(n_2039),
.Y(n_2706)
);

BUFx2_ASAP7_75t_L g2707 ( 
.A(n_2597),
.Y(n_2707)
);

AOI22xp33_ASAP7_75t_L g2708 ( 
.A1(n_2627),
.A2(n_2037),
.B1(n_2095),
.B2(n_2020),
.Y(n_2708)
);

AOI22xp33_ASAP7_75t_L g2709 ( 
.A1(n_2666),
.A2(n_2095),
.B1(n_2020),
.B2(n_2028),
.Y(n_2709)
);

OAI21x1_ASAP7_75t_L g2710 ( 
.A1(n_2649),
.A2(n_2372),
.B(n_2304),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_SL g2711 ( 
.A1(n_2642),
.A2(n_2506),
.B1(n_2466),
.B2(n_2579),
.Y(n_2711)
);

OR2x2_ASAP7_75t_L g2712 ( 
.A(n_2617),
.B(n_2578),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2631),
.B(n_2298),
.Y(n_2713)
);

AOI22xp33_ASAP7_75t_L g2714 ( 
.A1(n_2634),
.A2(n_2028),
.B1(n_2014),
.B2(n_2512),
.Y(n_2714)
);

AOI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2664),
.A2(n_2512),
.B1(n_2465),
.B2(n_2527),
.Y(n_2715)
);

AOI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2655),
.A2(n_2635),
.B1(n_2667),
.B2(n_2622),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2596),
.B(n_2652),
.Y(n_2717)
);

AOI221xp5_ASAP7_75t_L g2718 ( 
.A1(n_2653),
.A2(n_2014),
.B1(n_2578),
.B2(n_2426),
.C(n_2388),
.Y(n_2718)
);

AOI22xp33_ASAP7_75t_L g2719 ( 
.A1(n_2643),
.A2(n_2296),
.B1(n_2466),
.B2(n_2578),
.Y(n_2719)
);

AOI22xp33_ASAP7_75t_SL g2720 ( 
.A1(n_2662),
.A2(n_2466),
.B1(n_2296),
.B2(n_193),
.Y(n_2720)
);

AOI22xp33_ASAP7_75t_SL g2721 ( 
.A1(n_2650),
.A2(n_2466),
.B1(n_195),
.B2(n_191),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2707),
.B(n_2636),
.Y(n_2722)
);

NAND3xp33_ASAP7_75t_L g2723 ( 
.A(n_2683),
.B(n_2668),
.C(n_2665),
.Y(n_2723)
);

OAI21xp5_ASAP7_75t_SL g2724 ( 
.A1(n_2721),
.A2(n_2638),
.B(n_2644),
.Y(n_2724)
);

NAND4xp25_ASAP7_75t_L g2725 ( 
.A(n_2690),
.B(n_2682),
.C(n_2715),
.D(n_2686),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2676),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2678),
.B(n_2646),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2717),
.B(n_2651),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2687),
.B(n_2658),
.Y(n_2729)
);

OAI221xp5_ASAP7_75t_L g2730 ( 
.A1(n_2703),
.A2(n_2639),
.B1(n_2663),
.B2(n_2602),
.C(n_2645),
.Y(n_2730)
);

AOI22xp33_ASAP7_75t_L g2731 ( 
.A1(n_2674),
.A2(n_2670),
.B1(n_2720),
.B2(n_2675),
.Y(n_2731)
);

OAI21xp5_ASAP7_75t_L g2732 ( 
.A1(n_2679),
.A2(n_2647),
.B(n_2659),
.Y(n_2732)
);

NAND3xp33_ASAP7_75t_L g2733 ( 
.A(n_2706),
.B(n_2656),
.C(n_2647),
.Y(n_2733)
);

NAND3xp33_ASAP7_75t_L g2734 ( 
.A(n_2718),
.B(n_2660),
.C(n_2654),
.Y(n_2734)
);

OAI21xp5_ASAP7_75t_L g2735 ( 
.A1(n_2673),
.A2(n_2654),
.B(n_2610),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2677),
.B(n_2601),
.Y(n_2736)
);

OAI21xp5_ASAP7_75t_SL g2737 ( 
.A1(n_2671),
.A2(n_2601),
.B(n_2657),
.Y(n_2737)
);

OAI221xp5_ASAP7_75t_SL g2738 ( 
.A1(n_2716),
.A2(n_2694),
.B1(n_2700),
.B2(n_2719),
.C(n_2684),
.Y(n_2738)
);

OAI221xp5_ASAP7_75t_L g2739 ( 
.A1(n_2672),
.A2(n_2699),
.B1(n_2708),
.B2(n_2692),
.C(n_2688),
.Y(n_2739)
);

NAND3xp33_ASAP7_75t_L g2740 ( 
.A(n_2673),
.B(n_191),
.C(n_192),
.Y(n_2740)
);

OR2x2_ASAP7_75t_L g2741 ( 
.A(n_2701),
.B(n_2614),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2712),
.B(n_192),
.Y(n_2742)
);

NAND3xp33_ASAP7_75t_L g2743 ( 
.A(n_2714),
.B(n_196),
.C(n_197),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2681),
.B(n_197),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_SL g2745 ( 
.A1(n_2701),
.A2(n_201),
.B1(n_198),
.B2(n_199),
.Y(n_2745)
);

OA21x2_ASAP7_75t_L g2746 ( 
.A1(n_2681),
.A2(n_198),
.B(n_202),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2698),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2711),
.B(n_1772),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2695),
.B(n_203),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2713),
.B(n_204),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2713),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2685),
.B(n_206),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_SL g2753 ( 
.A(n_2685),
.B(n_1829),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2680),
.B(n_206),
.Y(n_2754)
);

NAND3xp33_ASAP7_75t_L g2755 ( 
.A(n_2704),
.B(n_207),
.C(n_208),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2702),
.B(n_208),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2702),
.B(n_209),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2691),
.B(n_210),
.Y(n_2758)
);

OR2x2_ASAP7_75t_L g2759 ( 
.A(n_2722),
.B(n_2696),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2741),
.B(n_2710),
.Y(n_2760)
);

NAND4xp75_ASAP7_75t_L g2761 ( 
.A(n_2746),
.B(n_2696),
.C(n_2693),
.D(n_2697),
.Y(n_2761)
);

NAND3xp33_ASAP7_75t_L g2762 ( 
.A(n_2740),
.B(n_2745),
.C(n_2755),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2751),
.B(n_211),
.Y(n_2763)
);

NAND4xp75_ASAP7_75t_L g2764 ( 
.A(n_2746),
.B(n_2756),
.C(n_2757),
.D(n_2732),
.Y(n_2764)
);

OAI211xp5_ASAP7_75t_SL g2765 ( 
.A1(n_2745),
.A2(n_2705),
.B(n_2709),
.C(n_2689),
.Y(n_2765)
);

OR2x2_ASAP7_75t_L g2766 ( 
.A(n_2728),
.B(n_211),
.Y(n_2766)
);

BUFx2_ASAP7_75t_L g2767 ( 
.A(n_2736),
.Y(n_2767)
);

AOI22xp33_ASAP7_75t_SL g2768 ( 
.A1(n_2723),
.A2(n_213),
.B1(n_215),
.B2(n_217),
.Y(n_2768)
);

AOI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2725),
.A2(n_2731),
.B1(n_2739),
.B2(n_2747),
.Y(n_2769)
);

BUFx2_ASAP7_75t_L g2770 ( 
.A(n_2726),
.Y(n_2770)
);

OR2x2_ASAP7_75t_L g2771 ( 
.A(n_2727),
.B(n_213),
.Y(n_2771)
);

AOI22xp33_ASAP7_75t_L g2772 ( 
.A1(n_2731),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_2772)
);

OAI211xp5_ASAP7_75t_SL g2773 ( 
.A1(n_2724),
.A2(n_218),
.B(n_219),
.C(n_220),
.Y(n_2773)
);

NOR2x1_ASAP7_75t_SL g2774 ( 
.A(n_2737),
.B(n_221),
.Y(n_2774)
);

NAND3xp33_ASAP7_75t_L g2775 ( 
.A(n_2734),
.B(n_222),
.C(n_223),
.Y(n_2775)
);

AOI221xp5_ASAP7_75t_L g2776 ( 
.A1(n_2747),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.C(n_227),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2744),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2729),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2742),
.B(n_225),
.Y(n_2779)
);

NAND4xp75_ASAP7_75t_L g2780 ( 
.A(n_2735),
.B(n_229),
.C(n_230),
.D(n_231),
.Y(n_2780)
);

NAND3xp33_ASAP7_75t_L g2781 ( 
.A(n_2750),
.B(n_229),
.C(n_230),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2749),
.B(n_232),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2770),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2767),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2760),
.B(n_2758),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2759),
.B(n_2752),
.Y(n_2786)
);

INVx3_ASAP7_75t_L g2787 ( 
.A(n_2778),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2777),
.Y(n_2788)
);

INVxp67_ASAP7_75t_L g2789 ( 
.A(n_2764),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2779),
.B(n_2754),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2773),
.A2(n_2743),
.B1(n_2733),
.B2(n_2730),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2763),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2763),
.Y(n_2793)
);

XNOR2x1_ASAP7_75t_L g2794 ( 
.A(n_2782),
.B(n_232),
.Y(n_2794)
);

XOR2x2_ASAP7_75t_L g2795 ( 
.A(n_2774),
.B(n_2738),
.Y(n_2795)
);

XNOR2xp5_ASAP7_75t_L g2796 ( 
.A(n_2794),
.B(n_2769),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2788),
.Y(n_2797)
);

INVxp67_ASAP7_75t_L g2798 ( 
.A(n_2792),
.Y(n_2798)
);

INVxp67_ASAP7_75t_L g2799 ( 
.A(n_2793),
.Y(n_2799)
);

AOI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2789),
.A2(n_2773),
.B1(n_2762),
.B2(n_2780),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2786),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2797),
.Y(n_2802)
);

XNOR2xp5_ASAP7_75t_L g2803 ( 
.A(n_2796),
.B(n_2795),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2798),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2800),
.A2(n_2789),
.B1(n_2791),
.B2(n_2761),
.Y(n_2805)
);

INVx1_ASAP7_75t_SL g2806 ( 
.A(n_2801),
.Y(n_2806)
);

XNOR2xp5_ASAP7_75t_L g2807 ( 
.A(n_2799),
.B(n_2790),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2797),
.Y(n_2808)
);

INVx1_ASAP7_75t_SL g2809 ( 
.A(n_2807),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2802),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2802),
.Y(n_2811)
);

INVx1_ASAP7_75t_SL g2812 ( 
.A(n_2803),
.Y(n_2812)
);

OAI322xp33_ASAP7_75t_L g2813 ( 
.A1(n_2805),
.A2(n_2791),
.A3(n_2781),
.B1(n_2786),
.B2(n_2766),
.C1(n_2775),
.C2(n_2771),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2808),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2810),
.Y(n_2815)
);

OAI322xp33_ASAP7_75t_L g2816 ( 
.A1(n_2809),
.A2(n_2806),
.A3(n_2804),
.B1(n_2784),
.B2(n_2783),
.C1(n_2768),
.C2(n_2776),
.Y(n_2816)
);

AOI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2812),
.A2(n_2776),
.B1(n_2772),
.B2(n_2785),
.Y(n_2817)
);

INVx2_ASAP7_75t_SL g2818 ( 
.A(n_2814),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2818),
.Y(n_2819)
);

HB1xp67_ASAP7_75t_L g2820 ( 
.A(n_2815),
.Y(n_2820)
);

OAI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2817),
.A2(n_2811),
.B1(n_2738),
.B2(n_2813),
.Y(n_2821)
);

A2O1A1Ixp33_ASAP7_75t_SL g2822 ( 
.A1(n_2816),
.A2(n_2765),
.B(n_2787),
.C(n_235),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2815),
.Y(n_2823)
);

NOR2x1_ASAP7_75t_L g2824 ( 
.A(n_2819),
.B(n_2748),
.Y(n_2824)
);

AOI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2821),
.A2(n_2765),
.B1(n_2748),
.B2(n_2787),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2820),
.Y(n_2826)
);

AOI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2823),
.A2(n_2753),
.B1(n_234),
.B2(n_235),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2822),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2822),
.B(n_233),
.Y(n_2829)
);

NOR2x1_ASAP7_75t_L g2830 ( 
.A(n_2819),
.B(n_236),
.Y(n_2830)
);

AOI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2821),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2828),
.B(n_242),
.Y(n_2832)
);

NOR2x1_ASAP7_75t_L g2833 ( 
.A(n_2830),
.B(n_244),
.Y(n_2833)
);

AO22x2_ASAP7_75t_L g2834 ( 
.A1(n_2826),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_2834)
);

INVx3_ASAP7_75t_L g2835 ( 
.A(n_2829),
.Y(n_2835)
);

INVxp67_ASAP7_75t_SL g2836 ( 
.A(n_2824),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2827),
.Y(n_2837)
);

AOI22xp33_ASAP7_75t_SL g2838 ( 
.A1(n_2831),
.A2(n_246),
.B1(n_249),
.B2(n_250),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2825),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2833),
.B(n_2835),
.Y(n_2840)
);

AO22x2_ASAP7_75t_L g2841 ( 
.A1(n_2836),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2834),
.Y(n_2842)
);

OR3x2_ASAP7_75t_L g2843 ( 
.A(n_2839),
.B(n_251),
.C(n_252),
.Y(n_2843)
);

AOI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2837),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2832),
.Y(n_2845)
);

AOI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2838),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_2846)
);

OAI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2838),
.A2(n_257),
.B1(n_259),
.B2(n_261),
.Y(n_2847)
);

INVx2_ASAP7_75t_SL g2848 ( 
.A(n_2841),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2841),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2840),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2842),
.Y(n_2851)
);

BUFx8_ASAP7_75t_L g2852 ( 
.A(n_2845),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2843),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2844),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2847),
.Y(n_2855)
);

AO22x2_ASAP7_75t_L g2856 ( 
.A1(n_2848),
.A2(n_2846),
.B1(n_263),
.B2(n_264),
.Y(n_2856)
);

AO22x2_ASAP7_75t_L g2857 ( 
.A1(n_2849),
.A2(n_262),
.B1(n_263),
.B2(n_266),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2853),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_2858)
);

AOI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_2851),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2852),
.Y(n_2860)
);

AO22x2_ASAP7_75t_L g2861 ( 
.A1(n_2855),
.A2(n_270),
.B1(n_271),
.B2(n_274),
.Y(n_2861)
);

OAI22xp5_ASAP7_75t_L g2862 ( 
.A1(n_2854),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2850),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2857),
.Y(n_2864)
);

INVxp67_ASAP7_75t_SL g2865 ( 
.A(n_2860),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2861),
.Y(n_2866)
);

XNOR2xp5_ASAP7_75t_L g2867 ( 
.A(n_2856),
.B(n_277),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2858),
.Y(n_2868)
);

INVxp67_ASAP7_75t_SL g2869 ( 
.A(n_2862),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2859),
.Y(n_2870)
);

AOI221xp5_ASAP7_75t_L g2871 ( 
.A1(n_2865),
.A2(n_2863),
.B1(n_282),
.B2(n_283),
.C(n_285),
.Y(n_2871)
);

AOI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2869),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_2872)
);

AOI22xp5_ASAP7_75t_L g2873 ( 
.A1(n_2868),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2872),
.Y(n_2874)
);

AOI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2874),
.A2(n_2864),
.B1(n_2866),
.B2(n_2870),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2875),
.Y(n_2876)
);

AOI221xp5_ASAP7_75t_L g2877 ( 
.A1(n_2876),
.A2(n_2867),
.B1(n_2871),
.B2(n_2873),
.C(n_292),
.Y(n_2877)
);

AOI211xp5_ASAP7_75t_L g2878 ( 
.A1(n_2877),
.A2(n_287),
.B(n_289),
.C(n_291),
.Y(n_2878)
);


endmodule