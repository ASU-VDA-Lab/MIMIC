module real_jpeg_21905_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_346, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_346;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_0),
.A2(n_22),
.B1(n_24),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_0),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_0),
.A2(n_68),
.B1(n_69),
.B2(n_92),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_0),
.A2(n_50),
.B1(n_52),
.B2(n_92),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_1),
.A2(n_22),
.B1(n_24),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_61),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_1),
.A2(n_61),
.B1(n_68),
.B2(n_69),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_1),
.A2(n_50),
.B1(n_52),
.B2(n_61),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_21),
.B1(n_31),
.B2(n_32),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_2),
.A2(n_21),
.B1(n_68),
.B2(n_69),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_2),
.A2(n_21),
.B1(n_50),
.B2(n_52),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_22),
.B1(n_24),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_3),
.A2(n_34),
.B1(n_50),
.B2(n_52),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_3),
.A2(n_34),
.B1(n_68),
.B2(n_69),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_4),
.A2(n_68),
.B1(n_69),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_4),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_4),
.A2(n_50),
.B1(n_52),
.B2(n_128),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_128),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_4),
.A2(n_22),
.B1(n_24),
.B2(n_128),
.Y(n_264)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_6),
.A2(n_52),
.B(n_64),
.C(n_108),
.D(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_6),
.B(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_6),
.B(n_49),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_6),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_6),
.A2(n_129),
.B(n_131),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_6),
.A2(n_31),
.B(n_46),
.C(n_167),
.D(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_6),
.B(n_31),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_35),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_6),
.A2(n_22),
.B1(n_24),
.B2(n_147),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_6),
.A2(n_30),
.B(n_32),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_7),
.A2(n_22),
.B1(n_24),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_7),
.A2(n_59),
.B1(n_68),
.B2(n_69),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_7),
.A2(n_50),
.B1(n_52),
.B2(n_59),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_59),
.Y(n_280)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_8),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_8),
.A2(n_140),
.B1(n_177),
.B2(n_192),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_50),
.B1(n_52),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_10),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_10),
.A2(n_68),
.B1(n_69),
.B2(n_111),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_111),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_10),
.A2(n_22),
.B1(n_24),
.B2(n_111),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_12),
.A2(n_50),
.B1(n_52),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_12),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_12),
.A2(n_68),
.B1(n_69),
.B2(n_123),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_123),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_12),
.A2(n_22),
.B1(n_24),
.B2(n_123),
.Y(n_235)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_38),
.B(n_341),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_36),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_19),
.B(n_40),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_19),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_25),
.B1(n_33),
.B2(n_35),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_20),
.A2(n_25),
.B1(n_35),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_27),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_22),
.A2(n_27),
.B(n_147),
.C(n_219),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_33),
.B(n_35),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_25),
.B(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_26),
.A2(n_29),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_26),
.A2(n_29),
.B1(n_58),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_26),
.A2(n_29),
.B1(n_235),
.B2(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_26),
.A2(n_213),
.B(n_264),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_29),
.A2(n_235),
.B(n_236),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_29),
.A2(n_91),
.B(n_236),
.Y(n_306)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_35),
.B(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_37),
.B(n_343),
.Y(n_342)
);

OAI21x1_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_78),
.B(n_340),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_73),
.C(n_75),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_42),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_56),
.C(n_62),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_44),
.B1(n_62),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_45),
.A2(n_53),
.B1(n_54),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_45),
.A2(n_54),
.B1(n_186),
.B2(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_45),
.A2(n_208),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_49),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_46),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_46),
.A2(n_49),
.B1(n_261),
.B2(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_46),
.A2(n_49),
.B1(n_97),
.B2(n_280),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_48),
.Y(n_175)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_50),
.B(n_51),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_52),
.A2(n_167),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_54),
.B(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_54),
.A2(n_186),
.B(n_187),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_54),
.A2(n_187),
.B(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_57),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_62),
.A2(n_89),
.B1(n_94),
.B2(n_95),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_71),
.B(n_72),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_63),
.A2(n_71),
.B1(n_122),
.B2(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_63),
.A2(n_165),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_63),
.A2(n_71),
.B1(n_205),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_63),
.A2(n_71),
.B1(n_246),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_63),
.A2(n_71),
.B1(n_255),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_64),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_64),
.A2(n_67),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx9p33_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_65),
.B(n_69),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_68),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_68),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_69),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_71),
.B(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_71),
.A2(n_124),
.B(n_205),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_72),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_98),
.B(n_339),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_80),
.B(n_84),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.C(n_93),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_325),
.Y(n_331)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_90),
.C(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_90),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_90),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_93),
.B(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI321xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_322),
.A3(n_332),
.B1(n_337),
.B2(n_338),
.C(n_345),
.Y(n_98)
);

AOI321xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_272),
.A3(n_310),
.B1(n_316),
.B2(n_321),
.C(n_346),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_229),
.C(n_268),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_199),
.B(n_228),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_180),
.B(n_198),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_159),
.B(n_179),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_135),
.B(n_158),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_106),
.B(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_112),
.B1(n_113),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_109),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_121),
.C(n_126),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_129),
.B(n_131),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_133),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_129),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_129),
.A2(n_223),
.B1(n_224),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_129),
.A2(n_149),
.B1(n_244),
.B2(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_129),
.A2(n_149),
.B(n_253),
.Y(n_285)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_151),
.B(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_134),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_144),
.B(n_157),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_142),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_152),
.B(n_156),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_148),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_149),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_172),
.B2(n_178),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_166),
.B1(n_170),
.B2(n_171),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_171),
.C(n_178),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_168),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_172),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_181),
.B(n_182),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_194),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_195),
.C(n_196),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_189),
.B2(n_193),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_190),
.C(n_191),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_189),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_201),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_215),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_202),
.B(n_216),
.C(n_227),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_204),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_209),
.C(n_210),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_216),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_221),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_230),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_248),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_231),
.B(n_248),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_242),
.C(n_247),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_241),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_234),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_247),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_245),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_266),
.B2(n_267),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_251),
.B(n_256),
.C(n_267),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_254),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_262),
.C(n_265),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_259),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_269),
.B(n_270),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_290),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_273),
.B(n_290),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.C(n_289),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_274),
.A2(n_275),
.B1(n_283),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_288),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_285),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_284),
.A2(n_302),
.B(n_306),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_286),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_287),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_308),
.B2(n_309),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_300),
.B2(n_301),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_301),
.C(n_309),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_298),
.B(n_299),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_298),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_299),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_299),
.A2(n_324),
.B1(n_328),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_307),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_304),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_308),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_311),
.A2(n_317),
.B(n_320),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_313),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_330),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_330),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.C(n_329),
.Y(n_323)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_324),
.Y(n_336)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);


endmodule