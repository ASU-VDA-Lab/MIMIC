module fake_jpeg_29190_n_138 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_138);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_19),
.B(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_30),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_79),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_57),
.B1(n_45),
.B2(n_48),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_46),
.B1(n_22),
.B2(n_23),
.Y(n_86)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_80),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_42),
.B1(n_57),
.B2(n_45),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_85)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_51),
.B(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_58),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_55),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_87),
.C(n_25),
.Y(n_114)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_18),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_20),
.B1(n_39),
.B2(n_35),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_96),
.Y(n_103)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_74),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_101),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_89),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_29),
.C(n_31),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_6),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_7),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_110),
.B1(n_113),
.B2(n_9),
.Y(n_119)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_7),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_8),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_114),
.B(n_115),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_8),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_27),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_117)
);

NOR2xp67_ASAP7_75t_R g126 ( 
.A(n_117),
.B(n_119),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_9),
.B1(n_17),
.B2(n_24),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_125),
.C(n_114),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_33),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_125),
.B1(n_120),
.B2(n_117),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_103),
.C(n_109),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_131),
.B(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_124),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_118),
.B(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_130),
.B(n_121),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_137),
.Y(n_138)
);


endmodule