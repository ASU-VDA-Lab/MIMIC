module real_jpeg_7431_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_3;

output n_7;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_11;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_8;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_1),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_16),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_4),
.B(n_66),
.C(n_69),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_4),
.A2(n_26),
.B1(n_79),
.B2(n_82),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_24),
.B1(n_32),
.B2(n_36),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_6),
.A2(n_36),
.B1(n_73),
.B2(n_76),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_56),
.Y(n_7)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_37),
.B(n_55),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_17),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_15),
.Y(n_10)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_12),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_20),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_28),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_19),
.B(n_43),
.Y(n_99)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_24),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_51),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_50),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_72),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_100),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_96),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_70),
.B1(n_94),
.B2(n_95),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_60),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_86),
.B1(n_89),
.B2(n_91),
.Y(n_85)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_84),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);


endmodule