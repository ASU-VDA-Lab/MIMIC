module fake_jpeg_23547_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_4),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx6_ASAP7_75t_SL g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_1),
.B(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_16),
.B(n_18),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_12),
.B1(n_9),
.B2(n_8),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_17),
.B1(n_21),
.B2(n_19),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_0),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx10_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_6),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_13),
.C(n_8),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_13),
.C(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_27),
.B(n_28),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_SL g27 ( 
.A1(n_17),
.A2(n_1),
.B(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_25),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_31),
.A3(n_29),
.B1(n_27),
.B2(n_24),
.C1(n_17),
.C2(n_16),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_34),
.C(n_33),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_35),
.Y(n_38)
);


endmodule