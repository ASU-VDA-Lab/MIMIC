module fake_netlist_1_6243_n_694 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_694);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_694;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g81 ( .A(n_1), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_30), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_67), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_66), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_23), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_65), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_36), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_69), .Y(n_89) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_32), .Y(n_90) );
CKINVDCx14_ASAP7_75t_R g91 ( .A(n_61), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_5), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_78), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_18), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_57), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_55), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_48), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_35), .Y(n_98) );
INVx3_ASAP7_75t_L g99 ( .A(n_72), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_38), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_75), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_74), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_53), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_76), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_52), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_54), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_68), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_44), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_7), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_56), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_47), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_6), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_39), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_43), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_3), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_45), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_1), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_29), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_24), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_7), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_70), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_25), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_46), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_16), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_37), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_99), .B(n_0), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_91), .Y(n_131) );
NOR2xp33_ASAP7_75t_SL g132 ( .A(n_93), .B(n_28), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_128), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_91), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_99), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_88), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_99), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_88), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_83), .A2(n_27), .B(n_79), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_128), .Y(n_142) );
NOR2xp67_ASAP7_75t_L g143 ( .A(n_94), .B(n_0), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_104), .B(n_2), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_96), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_104), .B(n_2), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_96), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_89), .B(n_4), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_94), .B(n_4), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_92), .B(n_5), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_85), .Y(n_152) );
NOR2xp67_ASAP7_75t_L g153 ( .A(n_105), .B(n_6), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_97), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_86), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_106), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_89), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_97), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_111), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_98), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_114), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_108), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g163 ( .A(n_93), .B(n_34), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_100), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_118), .B(n_8), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_119), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_108), .Y(n_167) );
AND2x6_ASAP7_75t_L g168 ( .A(n_101), .B(n_40), .Y(n_168) );
INVx5_ASAP7_75t_L g169 ( .A(n_89), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_121), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_84), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_124), .B(n_9), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_121), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_144), .B(n_81), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_131), .B(n_113), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
OR2x2_ASAP7_75t_L g177 ( .A(n_144), .B(n_116), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_146), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_151), .B(n_121), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_131), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_169), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
OAI21xp33_ASAP7_75t_L g185 ( .A1(n_160), .A2(n_113), .B(n_109), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_137), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_169), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
AO22x2_ASAP7_75t_L g190 ( .A1(n_151), .A2(n_129), .B1(n_127), .B2(n_126), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_169), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_171), .B(n_84), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_172), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_169), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_172), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_169), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_140), .B(n_109), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_146), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_172), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_140), .B(n_112), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_171), .A2(n_121), .B1(n_95), .B2(n_115), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_169), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_133), .Y(n_205) );
OAI21xp33_ASAP7_75t_L g206 ( .A1(n_160), .A2(n_110), .B(n_123), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_134), .B(n_107), .Y(n_207) );
AO22x2_ASAP7_75t_L g208 ( .A1(n_149), .A2(n_122), .B1(n_120), .B2(n_117), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_133), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_142), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_152), .B(n_121), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_142), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_130), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_150), .B(n_125), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_138), .Y(n_215) );
OR2x6_ASAP7_75t_L g216 ( .A(n_149), .B(n_103), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_134), .B(n_102), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_156), .B(n_89), .Y(n_218) );
INVxp67_ASAP7_75t_L g219 ( .A(n_136), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_152), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_159), .B(n_90), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_138), .Y(n_222) );
OR2x2_ASAP7_75t_L g223 ( .A(n_161), .B(n_9), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_166), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_155), .B(n_90), .Y(n_225) );
INVx5_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_155), .B(n_90), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_164), .B(n_90), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_164), .B(n_90), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_168), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_143), .B(n_10), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_165), .Y(n_233) );
AND2x6_ASAP7_75t_L g234 ( .A(n_168), .B(n_41), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_138), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_213), .B(n_168), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_205), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_233), .B(n_136), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_180), .B(n_153), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_228), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_216), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_205), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_221), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_228), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_205), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_231), .Y(n_247) );
BUFx8_ASAP7_75t_L g248 ( .A(n_182), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_213), .B(n_168), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_210), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_186), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_199), .B(n_168), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_180), .B(n_167), .Y(n_254) );
INVxp67_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_186), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_219), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_212), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_191), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_191), .Y(n_260) );
BUFx2_ASAP7_75t_SL g261 ( .A(n_226), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_216), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_226), .B(n_132), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_181), .Y(n_265) );
NOR3xp33_ASAP7_75t_SL g266 ( .A(n_185), .B(n_158), .C(n_139), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_176), .A2(n_141), .B(n_148), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_181), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_216), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_189), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_181), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_200), .B(n_173), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_225), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_200), .B(n_170), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_214), .B(n_163), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_214), .B(n_167), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_216), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_226), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_226), .Y(n_279) );
INVx3_ASAP7_75t_L g280 ( .A(n_211), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_174), .B(n_10), .Y(n_281) );
NOR2xp33_ASAP7_75t_SL g282 ( .A(n_234), .B(n_139), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_174), .B(n_158), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_177), .B(n_162), .Y(n_284) );
NOR2xp33_ASAP7_75t_R g285 ( .A(n_189), .B(n_145), .Y(n_285) );
NOR3xp33_ASAP7_75t_SL g286 ( .A(n_193), .B(n_147), .C(n_154), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_224), .B(n_141), .Y(n_287) );
BUFx8_ASAP7_75t_L g288 ( .A(n_234), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_190), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_177), .Y(n_290) );
NAND2x1p5_ASAP7_75t_L g291 ( .A(n_189), .B(n_141), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_208), .B(n_141), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_176), .B(n_157), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_223), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_225), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_220), .Y(n_296) );
AND3x1_ASAP7_75t_SL g297 ( .A(n_208), .B(n_11), .C(n_13), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_211), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_194), .A2(n_157), .B(n_14), .C(n_15), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_190), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_211), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_248), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_294), .B(n_208), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_289), .B(n_226), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_248), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_289), .A2(n_194), .B1(n_196), .B2(n_197), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_300), .A2(n_208), .B1(n_190), .B2(n_232), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_236), .A2(n_196), .B(n_179), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_250), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_300), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_281), .A2(n_190), .B1(n_232), .B2(n_201), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_240), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_281), .B(n_232), .Y(n_313) );
CKINVDCx6p67_ASAP7_75t_R g314 ( .A(n_262), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_252), .Y(n_315) );
OAI21xp33_ASAP7_75t_L g316 ( .A1(n_292), .A2(n_202), .B(n_209), .Y(n_316) );
CKINVDCx16_ASAP7_75t_R g317 ( .A(n_262), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_265), .Y(n_318) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_241), .B(n_223), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_241), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_248), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_237), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_237), .Y(n_323) );
BUFx10_ASAP7_75t_L g324 ( .A(n_269), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_265), .Y(n_325) );
BUFx4f_ASAP7_75t_SL g326 ( .A(n_257), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_290), .B(n_203), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_282), .B(n_207), .Y(n_328) );
BUFx12f_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_281), .B(n_217), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_242), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_242), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_277), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_239), .B(n_178), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_265), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_277), .A2(n_220), .B1(n_178), .B2(n_206), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_268), .B(n_218), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_240), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_254), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_268), .B(n_240), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_255), .B(n_175), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_268), .B(n_234), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_239), .B(n_234), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_288), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_270), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_239), .B(n_234), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_249), .A2(n_229), .B(n_230), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_292), .A2(n_234), .B1(n_227), .B2(n_195), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_254), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_276), .A2(n_195), .B1(n_183), .B2(n_187), .C(n_204), .Y(n_350) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_283), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_288), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_251), .B(n_183), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_275), .B(n_187), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_288), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_319), .A2(n_257), .B1(n_283), .B2(n_238), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_319), .B(n_251), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_339), .B(n_284), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_339), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_308), .A2(n_253), .B(n_287), .Y(n_360) );
OAI33xp33_ASAP7_75t_L g361 ( .A1(n_330), .A2(n_274), .A3(n_272), .B1(n_243), .B2(n_245), .B3(n_273), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_313), .B(n_261), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_343), .A2(n_263), .B(n_258), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_346), .A2(n_267), .B(n_270), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_326), .A2(n_284), .B1(n_295), .B2(n_296), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_319), .B(n_256), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_349), .Y(n_367) );
NAND2xp33_ASAP7_75t_R g368 ( .A(n_313), .B(n_285), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_347), .A2(n_246), .B(n_291), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_349), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_303), .B(n_295), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_309), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_309), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_315), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_328), .A2(n_291), .B(n_293), .Y(n_375) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_316), .A2(n_299), .B(n_264), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_315), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_334), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_351), .A2(n_271), .B1(n_280), .B2(n_301), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_322), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_351), .A2(n_280), .B1(n_301), .B2(n_298), .Y(n_381) );
A2O1A1Ixp33_ASAP7_75t_L g382 ( .A1(n_316), .A2(n_256), .B(n_259), .C(n_260), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_333), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_322), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_311), .A2(n_260), .B1(n_259), .B2(n_298), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_302), .A2(n_297), .B1(n_266), .B2(n_286), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_305), .A2(n_280), .B1(n_291), .B2(n_247), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_305), .Y(n_388) );
AND2x6_ASAP7_75t_L g389 ( .A(n_342), .B(n_244), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_356), .A2(n_307), .B1(n_313), .B2(n_310), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_372), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_383), .B(n_303), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_357), .A2(n_317), .B1(n_324), .B2(n_355), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_373), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_374), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_365), .A2(n_313), .B1(n_355), .B2(n_344), .Y(n_396) );
NAND3xp33_ASAP7_75t_L g397 ( .A(n_386), .B(n_348), .C(n_336), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
AOI222xp33_ASAP7_75t_L g399 ( .A1(n_358), .A2(n_321), .B1(n_341), .B2(n_327), .C1(n_378), .C2(n_361), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_357), .B(n_333), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_380), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_362), .A2(n_310), .B1(n_320), .B2(n_314), .Y(n_402) );
BUFx4f_ASAP7_75t_L g403 ( .A(n_362), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_377), .B(n_341), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_359), .A2(n_336), .B1(n_350), .B2(n_306), .C(n_317), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_366), .A2(n_344), .B1(n_314), .B2(n_352), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_362), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_366), .A2(n_352), .B1(n_329), .B2(n_320), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_369), .A2(n_354), .B(n_323), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_384), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_367), .A2(n_352), .B1(n_329), .B2(n_342), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_370), .B(n_353), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_371), .A2(n_342), .B1(n_324), .B2(n_325), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_385), .A2(n_318), .B1(n_335), .B2(n_325), .C(n_353), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_384), .Y(n_416) );
OR2x6_ASAP7_75t_L g417 ( .A(n_363), .B(n_342), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_324), .B1(n_318), .B2(n_335), .C1(n_325), .C2(n_345), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_403), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_416), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_397), .B(n_399), .C(n_405), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_403), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_401), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_403), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_398), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_401), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_402), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_409), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_409), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_416), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_391), .Y(n_431) );
NAND5xp2_ASAP7_75t_L g432 ( .A(n_393), .B(n_379), .C(n_381), .D(n_368), .E(n_324), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_411), .B(n_382), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_398), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
AO21x2_ASAP7_75t_L g436 ( .A1(n_410), .A2(n_382), .B(n_376), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
OAI31xp33_ASAP7_75t_SL g438 ( .A1(n_390), .A2(n_387), .A3(n_368), .B(n_375), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_411), .Y(n_439) );
INVx4_ASAP7_75t_L g440 ( .A(n_407), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_395), .B(n_376), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_394), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_400), .B(n_345), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_413), .Y(n_444) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_404), .A2(n_360), .B(n_364), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_392), .B(n_388), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_400), .A2(n_389), .B1(n_318), .B2(n_335), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_417), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_407), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_413), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g451 ( .A1(n_396), .A2(n_323), .B1(n_332), .B2(n_331), .C(n_340), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_417), .Y(n_452) );
OR2x6_ASAP7_75t_L g453 ( .A(n_417), .B(n_375), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_429), .B(n_392), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_431), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_429), .B(n_417), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_450), .B(n_406), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_431), .B(n_11), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_435), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_450), .B(n_408), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g461 ( .A1(n_421), .A2(n_412), .B1(n_414), .B2(n_418), .C(n_415), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_435), .B(n_14), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_437), .B(n_389), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_421), .A2(n_337), .B1(n_340), .B2(n_304), .C(n_332), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_423), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_437), .B(n_389), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_444), .B(n_389), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_443), .B(n_15), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_420), .B(n_16), .Y(n_469) );
BUFx3_ASAP7_75t_L g470 ( .A(n_434), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_428), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_428), .Y(n_472) );
AND2x2_ASAP7_75t_SL g473 ( .A(n_427), .B(n_389), .Y(n_473) );
OAI31xp33_ASAP7_75t_L g474 ( .A1(n_432), .A2(n_340), .A3(n_331), .B(n_19), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_444), .B(n_389), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_443), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_423), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_438), .B(n_157), .C(n_184), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_443), .B(n_17), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_427), .A2(n_338), .B1(n_312), .B2(n_337), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_420), .B(n_17), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_444), .B(n_18), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_430), .B(n_19), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_434), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_423), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_449), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_432), .A2(n_312), .B1(n_338), .B2(n_157), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_430), .B(n_157), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_426), .Y(n_489) );
OAI33xp33_ASAP7_75t_L g490 ( .A1(n_442), .A2(n_235), .A3(n_222), .B1(n_215), .B2(n_204), .B3(n_198), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_422), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_446), .B(n_235), .C(n_222), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_441), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_426), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_426), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_448), .B(n_338), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_439), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g499 ( .A1(n_442), .A2(n_215), .B1(n_188), .B2(n_184), .C(n_337), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_439), .B(n_20), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_439), .B(n_338), .Y(n_501) );
AOI33xp33_ASAP7_75t_L g502 ( .A1(n_447), .A2(n_198), .A3(n_192), .B1(n_26), .B2(n_31), .B3(n_33), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_446), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_476), .B(n_449), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_465), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_484), .B(n_446), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_454), .B(n_503), .Y(n_507) );
INVx4_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_455), .B(n_452), .Y(n_509) );
BUFx3_ASAP7_75t_L g510 ( .A(n_470), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_455), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_470), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_465), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_459), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_468), .B(n_440), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_459), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_469), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_474), .A2(n_448), .B1(n_452), .B2(n_451), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_495), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_456), .B(n_448), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_495), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_498), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_456), .B(n_452), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_461), .B(n_451), .C(n_422), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_479), .B(n_440), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_479), .B(n_440), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_465), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_491), .B(n_448), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_474), .A2(n_448), .B1(n_440), .B2(n_419), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_469), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_498), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_491), .B(n_494), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_471), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_487), .A2(n_419), .B1(n_422), .B2(n_424), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_494), .B(n_453), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_484), .B(n_422), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_471), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_477), .B(n_453), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_477), .Y(n_539) );
INVx1_ASAP7_75t_SL g540 ( .A(n_470), .Y(n_540) );
OAI21xp33_ASAP7_75t_L g541 ( .A1(n_478), .A2(n_438), .B(n_425), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_481), .B(n_424), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_458), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_458), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_477), .B(n_453), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_485), .B(n_453), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
NAND2xp33_ASAP7_75t_R g548 ( .A(n_481), .B(n_424), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_485), .B(n_453), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_489), .B(n_453), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_489), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_472), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_473), .B(n_422), .Y(n_553) );
AND2x6_ASAP7_75t_SL g554 ( .A(n_462), .B(n_424), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_489), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_496), .B(n_433), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_496), .B(n_433), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_486), .B(n_472), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_483), .B(n_440), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_488), .B(n_433), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_511), .Y(n_562) );
OAI322xp33_ASAP7_75t_SL g563 ( .A1(n_507), .A2(n_460), .A3(n_457), .B1(n_482), .B2(n_463), .C1(n_466), .C2(n_475), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_511), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_541), .A2(n_478), .B(n_480), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_524), .A2(n_473), .B1(n_493), .B2(n_462), .Y(n_566) );
AOI211x1_ASAP7_75t_SL g567 ( .A1(n_534), .A2(n_480), .B(n_463), .C(n_466), .Y(n_567) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_517), .A2(n_483), .B1(n_490), .B2(n_488), .C(n_464), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_514), .Y(n_569) );
AOI222xp33_ASAP7_75t_L g570 ( .A1(n_543), .A2(n_424), .B1(n_467), .B2(n_425), .C1(n_492), .C2(n_500), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_532), .B(n_492), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_506), .B(n_502), .C(n_499), .Y(n_572) );
OAI211xp5_ASAP7_75t_SL g573 ( .A1(n_529), .A2(n_447), .B(n_425), .C(n_501), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_540), .B(n_497), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_537), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_532), .B(n_445), .Y(n_576) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_558), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_516), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_530), .B(n_445), .Y(n_579) );
AO22x1_ASAP7_75t_L g580 ( .A1(n_508), .A2(n_497), .B1(n_500), .B2(n_501), .Y(n_580) );
NAND2xp33_ASAP7_75t_L g581 ( .A(n_542), .B(n_497), .Y(n_581) );
NOR2xp67_ASAP7_75t_SL g582 ( .A(n_508), .B(n_338), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_519), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_544), .B(n_445), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_515), .B(n_497), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_512), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_523), .B(n_445), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_525), .B(n_436), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_521), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_521), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_553), .A2(n_436), .B(n_312), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_509), .B(n_436), .Y(n_592) );
XNOR2x1_ASAP7_75t_L g593 ( .A(n_510), .B(n_21), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_552), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_509), .B(n_436), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_558), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g597 ( .A1(n_508), .A2(n_312), .B(n_42), .C(n_49), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_505), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_522), .Y(n_599) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_518), .A2(n_188), .B1(n_184), .B2(n_312), .C(n_192), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_561), .B(n_22), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_561), .B(n_50), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_522), .Y(n_603) );
NOR2xp67_ASAP7_75t_L g604 ( .A(n_533), .B(n_51), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_531), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_556), .B(n_58), .Y(n_606) );
AOI21xp33_ASAP7_75t_SL g607 ( .A1(n_548), .A2(n_59), .B(n_60), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_531), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_536), .B(n_62), .Y(n_609) );
NOR3xp33_ASAP7_75t_SL g610 ( .A(n_573), .B(n_504), .C(n_526), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_586), .B(n_552), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_596), .B(n_523), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_562), .Y(n_613) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_604), .B(n_559), .Y(n_614) );
NOR4xp25_ASAP7_75t_SL g615 ( .A(n_607), .B(n_554), .C(n_539), .D(n_547), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_577), .B(n_557), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_594), .B(n_575), .Y(n_617) );
AND4x1_ASAP7_75t_L g618 ( .A(n_566), .B(n_535), .C(n_550), .D(n_549), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_573), .A2(n_520), .B1(n_535), .B2(n_528), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_587), .B(n_557), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_564), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_574), .B(n_520), .Y(n_622) );
NOR2xp33_ASAP7_75t_R g623 ( .A(n_581), .B(n_550), .Y(n_623) );
NOR2x1_ASAP7_75t_L g624 ( .A(n_597), .B(n_555), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_565), .B(n_528), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_576), .B(n_556), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_597), .B(n_539), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g628 ( .A1(n_594), .A2(n_545), .B(n_538), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_569), .Y(n_629) );
AND3x2_ASAP7_75t_L g630 ( .A(n_568), .B(n_609), .C(n_593), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_571), .B(n_520), .Y(n_631) );
O2A1O1Ixp5_ASAP7_75t_SL g632 ( .A1(n_601), .A2(n_555), .B(n_547), .C(n_551), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_568), .B(n_551), .C(n_538), .Y(n_633) );
NOR2xp33_ASAP7_75t_R g634 ( .A(n_602), .B(n_545), .Y(n_634) );
INVxp33_ASAP7_75t_L g635 ( .A(n_582), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_579), .B(n_549), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_598), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_585), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_584), .B(n_546), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_578), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_583), .B(n_546), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_608), .B(n_527), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_610), .A2(n_567), .B1(n_565), .B2(n_572), .C(n_570), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_624), .B(n_591), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_633), .A2(n_563), .B1(n_605), .B2(n_603), .C(n_589), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_630), .A2(n_588), .B1(n_600), .B2(n_606), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_613), .Y(n_647) );
XOR2xp5_ASAP7_75t_L g648 ( .A(n_619), .B(n_580), .Y(n_648) );
XOR2xp5_ASAP7_75t_L g649 ( .A(n_616), .B(n_590), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_617), .B(n_599), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_621), .Y(n_651) );
NAND3xp33_ASAP7_75t_SL g652 ( .A(n_615), .B(n_600), .C(n_591), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_622), .B(n_595), .Y(n_653) );
INVxp33_ASAP7_75t_SL g654 ( .A(n_611), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_629), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_638), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_627), .A2(n_592), .B1(n_560), .B2(n_527), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_637), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_611), .Y(n_659) );
NOR2xp33_ASAP7_75t_R g660 ( .A(n_630), .B(n_63), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_625), .A2(n_513), .B(n_71), .C(n_73), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_628), .A2(n_184), .B1(n_188), .B2(n_80), .Y(n_662) );
AOI22xp33_ASAP7_75t_R g663 ( .A1(n_660), .A2(n_623), .B1(n_634), .B2(n_640), .Y(n_663) );
AND2x2_ASAP7_75t_SL g664 ( .A(n_646), .B(n_618), .Y(n_664) );
OAI311xp33_ASAP7_75t_L g665 ( .A1(n_643), .A2(n_636), .A3(n_639), .B1(n_631), .C1(n_641), .Y(n_665) );
CKINVDCx16_ASAP7_75t_R g666 ( .A(n_659), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_645), .B(n_617), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_656), .B(n_614), .Y(n_668) );
AOI322xp5_ASAP7_75t_L g669 ( .A1(n_646), .A2(n_620), .A3(n_612), .B1(n_626), .B2(n_642), .C1(n_632), .C2(n_635), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_654), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_649), .B(n_64), .Y(n_671) );
AOI221xp5_ASAP7_75t_SL g672 ( .A1(n_648), .A2(n_184), .B1(n_188), .B2(n_77), .C(n_261), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_647), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_644), .A2(n_240), .B(n_244), .C(n_247), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_660), .A2(n_650), .B1(n_651), .B2(n_655), .C(n_652), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_661), .A2(n_278), .B1(n_279), .B2(n_662), .C(n_658), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g677 ( .A1(n_653), .A2(n_278), .B(n_279), .C(n_660), .Y(n_677) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_657), .B(n_278), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_645), .B(n_278), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_643), .A2(n_279), .B1(n_645), .B2(n_657), .C(n_563), .Y(n_680) );
NOR2x1_ASAP7_75t_L g681 ( .A(n_677), .B(n_678), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_673), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_666), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_670), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_679), .Y(n_685) );
INVx5_ASAP7_75t_SL g686 ( .A(n_684), .Y(n_686) );
NAND3xp33_ASAP7_75t_SL g687 ( .A(n_683), .B(n_675), .C(n_669), .Y(n_687) );
NOR4xp25_ASAP7_75t_SL g688 ( .A(n_685), .B(n_680), .C(n_676), .D(n_665), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_686), .Y(n_689) );
OAI22x1_ASAP7_75t_L g690 ( .A1(n_687), .A2(n_681), .B1(n_684), .B2(n_667), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_689), .Y(n_691) );
OAI222xp33_ASAP7_75t_L g692 ( .A1(n_690), .A2(n_663), .B1(n_688), .B2(n_682), .C1(n_668), .C2(n_671), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_691), .A2(n_664), .B1(n_668), .B2(n_672), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_693), .A2(n_692), .B(n_674), .Y(n_694) );
endmodule