module fake_ibex_1172_n_2257 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2257);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2257;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_641;
wire n_557;
wire n_1937;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2163;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2189;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_1326;
wire n_971;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_2256;
wire n_406;
wire n_737;
wire n_606;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_399;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2162;
wire n_2236;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_864;
wire n_608;
wire n_412;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_878;
wire n_474;
wire n_594;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_585;
wire n_1982;
wire n_2252;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_650;
wire n_409;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_2243;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_1830;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1642;
wire n_1455;
wire n_1871;
wire n_480;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2078;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_415;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2222;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_753;
wire n_2126;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_417;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1397;
wire n_1211;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2092;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_405;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_408;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_349),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_232),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_142),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_86),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_63),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_224),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_248),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_236),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_292),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_201),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_5),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_133),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_341),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_388),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_348),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_215),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_7),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_251),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_383),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_363),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_129),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_318),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_329),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_59),
.Y(n_422)
);

BUFx10_ASAP7_75t_L g423 ( 
.A(n_56),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_130),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_362),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_357),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_376),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_352),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_182),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_386),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_206),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_340),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_398),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_375),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_351),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_30),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_47),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_28),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_280),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_214),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_285),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_41),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_267),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_233),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_257),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_219),
.Y(n_448)
);

BUFx10_ASAP7_75t_L g449 ( 
.A(n_189),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_247),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_70),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_11),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_237),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_315),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_59),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_6),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_303),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_2),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_177),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_109),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_305),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_274),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_67),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_306),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_326),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_93),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_207),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_217),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_90),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_269),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_205),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_14),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_277),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_185),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_290),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_138),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_283),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_275),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_239),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_133),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_221),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_307),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_225),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_332),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_175),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_365),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_60),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_263),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_314),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_255),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_322),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_331),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_197),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_286),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_366),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_170),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_359),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_11),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_92),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_354),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_6),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_276),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_241),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_231),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_188),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_268),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_199),
.Y(n_509)
);

BUFx10_ASAP7_75t_L g510 ( 
.A(n_27),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_220),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_32),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_186),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_191),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_44),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_73),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_202),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_353),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_369),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_160),
.B(n_2),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_86),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_310),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_156),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_238),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_112),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_380),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_194),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_227),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_208),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_320),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_379),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_67),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_112),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_70),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_252),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_139),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_195),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_126),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_261),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_300),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_119),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_262),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_284),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_377),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_0),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_37),
.Y(n_546)
);

BUFx5_ASAP7_75t_L g547 ( 
.A(n_390),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_142),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_106),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_9),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_3),
.Y(n_551)
);

BUFx8_ASAP7_75t_SL g552 ( 
.A(n_166),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_155),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_167),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_68),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_226),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_395),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_216),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_222),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_254),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_66),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_218),
.Y(n_562)
);

BUFx8_ASAP7_75t_SL g563 ( 
.A(n_336),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_323),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_288),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_382),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_179),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_311),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_393),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_316),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_397),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_360),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_92),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_125),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_330),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_94),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_171),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_161),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_384),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_287),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_187),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_296),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_125),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_9),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_213),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_209),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_137),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_99),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_108),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_279),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_12),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_127),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_356),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_371),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_40),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_228),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_174),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_151),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_313),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_278),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_245),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_211),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_1),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_256),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_342),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_324),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_102),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_328),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_103),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_22),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_14),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_192),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_347),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_344),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_249),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_337),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_169),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_312),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_41),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_325),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_350),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_114),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_144),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_17),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_135),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_99),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_301),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_295),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_162),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_372),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_32),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_389),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_141),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_355),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_60),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_4),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_293),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_327),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_136),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_137),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_161),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_149),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_240),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_230),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_253),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_264),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_156),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_243),
.Y(n_648)
);

BUFx5_ASAP7_75t_L g649 ( 
.A(n_116),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_47),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_148),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_49),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_138),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_136),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_338),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_94),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_281),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_346),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_84),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_364),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_335),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_129),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_294),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_25),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_339),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_418),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_420),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_440),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_649),
.Y(n_669)
);

INVx5_ASAP7_75t_L g670 ( 
.A(n_449),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_514),
.B(n_5),
.Y(n_671)
);

BUFx8_ASAP7_75t_SL g672 ( 
.A(n_410),
.Y(n_672)
);

BUFx8_ASAP7_75t_L g673 ( 
.A(n_582),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_489),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_512),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_462),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_462),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_489),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_649),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_462),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_449),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_SL g682 ( 
.A(n_552),
.B(n_165),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_449),
.Y(n_683)
);

CKINVDCx16_ASAP7_75t_R g684 ( 
.A(n_549),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_440),
.B(n_8),
.Y(n_685)
);

BUFx8_ASAP7_75t_SL g686 ( 
.A(n_410),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_562),
.Y(n_687)
);

BUFx8_ASAP7_75t_SL g688 ( 
.A(n_470),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_525),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_445),
.B(n_8),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_450),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_423),
.B(n_10),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_423),
.B(n_12),
.Y(n_693)
);

AND2x6_ASAP7_75t_L g694 ( 
.A(n_494),
.B(n_168),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_462),
.Y(n_695)
);

BUFx8_ASAP7_75t_L g696 ( 
.A(n_445),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_476),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_470),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_525),
.B(n_13),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_546),
.Y(n_700)
);

OA21x2_ASAP7_75t_L g701 ( 
.A1(n_414),
.A2(n_173),
.B(n_172),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_649),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_649),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_450),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_546),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_649),
.Y(n_706)
);

OA21x2_ASAP7_75t_L g707 ( 
.A1(n_414),
.A2(n_178),
.B(n_176),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_450),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_622),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_510),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_622),
.B(n_15),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_468),
.B(n_15),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_510),
.Y(n_713)
);

OAI22x1_ASAP7_75t_SL g714 ( 
.A1(n_545),
.A2(n_573),
.B1(n_550),
.B2(n_619),
.Y(n_714)
);

INVx5_ASAP7_75t_L g715 ( 
.A(n_476),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_510),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_399),
.B(n_655),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_468),
.B(n_16),
.Y(n_718)
);

BUFx8_ASAP7_75t_L g719 ( 
.A(n_649),
.Y(n_719)
);

INVx5_ASAP7_75t_L g720 ( 
.A(n_476),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_451),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_451),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_409),
.B(n_16),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_456),
.B(n_494),
.Y(n_724)
);

OAI21x1_ASAP7_75t_L g725 ( 
.A1(n_509),
.A2(n_181),
.B(n_180),
.Y(n_725)
);

AOI22x1_ASAP7_75t_SL g726 ( 
.A1(n_545),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_451),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_451),
.Y(n_728)
);

INVxp33_ASAP7_75t_SL g729 ( 
.A(n_664),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_517),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_649),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_547),
.Y(n_732)
);

BUFx12f_ASAP7_75t_L g733 ( 
.A(n_616),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_533),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_422),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_547),
.Y(n_736)
);

AOI22x1_ASAP7_75t_SL g737 ( 
.A1(n_550),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_737)
);

INVx5_ASAP7_75t_L g738 ( 
.A(n_517),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_509),
.B(n_20),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_524),
.B(n_21),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_405),
.B(n_22),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_533),
.Y(n_742)
);

BUFx2_ASAP7_75t_L g743 ( 
.A(n_664),
.Y(n_743)
);

OA21x2_ASAP7_75t_L g744 ( 
.A1(n_518),
.A2(n_184),
.B(n_183),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_533),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_401),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_533),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_405),
.B(n_23),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_439),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_402),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_452),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_600),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_574),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_600),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_455),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_574),
.Y(n_756)
);

OA21x2_ASAP7_75t_L g757 ( 
.A1(n_518),
.A2(n_193),
.B(n_190),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_522),
.A2(n_198),
.B(n_196),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_574),
.Y(n_759)
);

AND2x6_ASAP7_75t_L g760 ( 
.A(n_617),
.B(n_200),
.Y(n_760)
);

BUFx12f_ASAP7_75t_L g761 ( 
.A(n_616),
.Y(n_761)
);

BUFx8_ASAP7_75t_SL g762 ( 
.A(n_573),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_574),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_733),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_685),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_733),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_698),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_761),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_743),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_676),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_717),
.B(n_416),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_685),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_729),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_685),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_761),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_729),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_669),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_672),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_750),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_672),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_699),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_686),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_686),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_698),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_688),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_688),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_750),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_762),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_762),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_675),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_684),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_675),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_699),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_669),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_746),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_673),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_673),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_679),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_673),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_SL g800 ( 
.A(n_740),
.B(n_428),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_667),
.B(n_416),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_714),
.Y(n_802)
);

NOR2xp67_ASAP7_75t_L g803 ( 
.A(n_670),
.B(n_404),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_719),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_711),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_719),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_719),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_670),
.B(n_406),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_689),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_716),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_670),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_683),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_741),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_711),
.Y(n_814)
);

INVx6_ASAP7_75t_L g815 ( 
.A(n_683),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_R g816 ( 
.A(n_713),
.B(n_428),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_694),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_711),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_674),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_683),
.Y(n_820)
);

BUFx10_ASAP7_75t_L g821 ( 
.A(n_710),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_691),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_679),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_691),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_691),
.B(n_411),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_691),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_678),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_704),
.B(n_522),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_702),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_704),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_704),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_R g832 ( 
.A(n_713),
.B(n_432),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_748),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_R g834 ( 
.A(n_710),
.B(n_432),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_692),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_678),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_694),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_708),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_R g839 ( 
.A(n_708),
.B(n_478),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_708),
.B(n_403),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_700),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_696),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_703),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_696),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_705),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_693),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_676),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_696),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_709),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_724),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_681),
.Y(n_851)
);

XOR2xp5_ASAP7_75t_L g852 ( 
.A(n_726),
.B(n_478),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_681),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_724),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_737),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_666),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_R g857 ( 
.A(n_682),
.B(n_490),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_687),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_690),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_712),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_703),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_735),
.B(n_417),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_671),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_730),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_749),
.B(n_426),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_730),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_751),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_668),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_706),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_755),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_718),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_752),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_752),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_723),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_739),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_739),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_732),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_738),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_706),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_732),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_694),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_694),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_760),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_731),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_738),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_738),
.B(n_431),
.Y(n_886)
);

INVx8_ASAP7_75t_L g887 ( 
.A(n_760),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_760),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_760),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_738),
.Y(n_890)
);

BUFx10_ASAP7_75t_L g891 ( 
.A(n_760),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_736),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_R g893 ( 
.A(n_754),
.B(n_490),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_754),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_754),
.B(n_415),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_R g896 ( 
.A(n_754),
.B(n_491),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_727),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_727),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_R g899 ( 
.A(n_763),
.B(n_491),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_763),
.B(n_419),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_701),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_753),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_676),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_753),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_701),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_SL g906 ( 
.A1(n_707),
.A2(n_528),
.B1(n_531),
.B2(n_502),
.Y(n_906)
);

CKINVDCx16_ASAP7_75t_R g907 ( 
.A(n_721),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_759),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_715),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_759),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_759),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_725),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_725),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_758),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_707),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_715),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_715),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_676),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_715),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_758),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_721),
.B(n_502),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_R g922 ( 
.A(n_721),
.B(n_528),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_721),
.Y(n_923)
);

INVx11_ASAP7_75t_L g924 ( 
.A(n_720),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_744),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_SL g926 ( 
.A(n_720),
.B(n_552),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_720),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_722),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_722),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_677),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_744),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_722),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_859),
.B(n_744),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_860),
.B(n_434),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_771),
.B(n_531),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_910),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_858),
.B(n_757),
.Y(n_937)
);

AOI221xp5_ASAP7_75t_L g938 ( 
.A1(n_819),
.A2(n_500),
.B1(n_501),
.B2(n_467),
.C(n_460),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_817),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_795),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_769),
.B(n_520),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_871),
.B(n_400),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_827),
.B(n_540),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_850),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_765),
.B(n_757),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_841),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_SL g947 ( 
.A(n_773),
.B(n_601),
.C(n_540),
.Y(n_947)
);

OA21x2_ASAP7_75t_L g948 ( 
.A1(n_912),
.A2(n_566),
.B(n_527),
.Y(n_948)
);

XOR2xp5_ASAP7_75t_L g949 ( 
.A(n_767),
.B(n_601),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_854),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_772),
.B(n_774),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_867),
.B(n_407),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_801),
.B(n_620),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_845),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_870),
.B(n_408),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_875),
.B(n_412),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_864),
.B(n_866),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_817),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_900),
.B(n_413),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_913),
.A2(n_757),
.B(n_441),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_851),
.B(n_421),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_842),
.B(n_425),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_779),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_853),
.B(n_427),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_781),
.B(n_436),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_844),
.B(n_429),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_836),
.B(n_430),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_821),
.B(n_433),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_848),
.B(n_435),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_849),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_779),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_877),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_787),
.Y(n_973)
);

INVxp33_ASAP7_75t_L g974 ( 
.A(n_834),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_821),
.B(n_863),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_L g976 ( 
.A(n_800),
.B(n_503),
.C(n_481),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_846),
.B(n_437),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_892),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_807),
.Y(n_979)
);

AND2x6_ASAP7_75t_L g980 ( 
.A(n_837),
.B(n_617),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_887),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_887),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_813),
.B(n_443),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_793),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_805),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_874),
.B(n_447),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_809),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_815),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_797),
.B(n_23),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_L g990 ( 
.A(n_887),
.B(n_547),
.Y(n_990)
);

NOR2x1p5_ASAP7_75t_L g991 ( 
.A(n_799),
.B(n_424),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_814),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_876),
.B(n_448),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_810),
.B(n_454),
.Y(n_994)
);

NOR2xp67_ASAP7_75t_L g995 ( 
.A(n_764),
.B(n_24),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_L g996 ( 
.A(n_881),
.B(n_547),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_818),
.B(n_442),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_909),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_880),
.B(n_446),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_856),
.B(n_457),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_862),
.Y(n_1001)
);

NAND3xp33_ASAP7_75t_L g1002 ( 
.A(n_882),
.B(n_444),
.C(n_438),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_SL g1003 ( 
.A(n_891),
.B(n_645),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_840),
.B(n_461),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_891),
.Y(n_1005)
);

INVxp33_ASAP7_75t_L g1006 ( 
.A(n_834),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_865),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_776),
.B(n_465),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_909),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_815),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_878),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_902),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_872),
.B(n_466),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_873),
.B(n_469),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_879),
.B(n_453),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_815),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_777),
.B(n_459),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_811),
.B(n_812),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_777),
.B(n_463),
.Y(n_1019)
);

XOR2xp5_ASAP7_75t_L g1020 ( 
.A(n_784),
.B(n_645),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_904),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_820),
.B(n_471),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_920),
.A2(n_532),
.B(n_555),
.C(n_523),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_790),
.B(n_515),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_822),
.B(n_472),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_883),
.B(n_474),
.Y(n_1026)
);

BUFx2_ASAP7_75t_R g1027 ( 
.A(n_778),
.Y(n_1027)
);

NOR3xp33_ASAP7_75t_L g1028 ( 
.A(n_906),
.B(n_625),
.C(n_607),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_792),
.B(n_458),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_895),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_L g1031 ( 
.A(n_855),
.B(n_473),
.C(n_464),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_888),
.B(n_889),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_804),
.B(n_806),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_L g1034 ( 
.A(n_802),
.B(n_516),
.C(n_477),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_824),
.B(n_475),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_908),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_911),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_794),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_826),
.B(n_480),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_830),
.B(n_483),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_831),
.B(n_486),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_905),
.A2(n_583),
.B1(n_584),
.B2(n_576),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_828),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_838),
.B(n_487),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_828),
.Y(n_1045)
);

NOR2x1p5_ASAP7_75t_L g1046 ( 
.A(n_780),
.B(n_521),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_897),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_898),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_L g1049 ( 
.A(n_782),
.B(n_536),
.C(n_534),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_907),
.B(n_496),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_798),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_803),
.B(n_498),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_808),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_798),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_825),
.B(n_505),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_886),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_766),
.B(n_538),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_893),
.B(n_511),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_893),
.B(n_519),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_896),
.B(n_526),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_926),
.B(n_548),
.C(n_541),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_783),
.B(n_553),
.C(n_551),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_835),
.B(n_529),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_914),
.B(n_530),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_823),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_833),
.B(n_535),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_839),
.B(n_539),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_823),
.B(n_829),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_816),
.B(n_561),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_931),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_925),
.B(n_588),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_925),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_839),
.B(n_543),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_L g1074 ( 
.A(n_768),
.B(n_24),
.Y(n_1074)
);

BUFx5_ASAP7_75t_L g1075 ( 
.A(n_923),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_770),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_775),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_785),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_832),
.B(n_578),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_885),
.B(n_560),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_843),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_861),
.B(n_565),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_861),
.B(n_567),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_786),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_L g1085 ( 
.A(n_788),
.B(n_589),
.C(n_587),
.Y(n_1085)
);

NOR2x1p5_ASAP7_75t_L g1086 ( 
.A(n_789),
.B(n_796),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_899),
.B(n_595),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_852),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_869),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_884),
.B(n_479),
.Y(n_1090)
);

NOR2xp67_ASAP7_75t_L g1091 ( 
.A(n_916),
.B(n_25),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_890),
.B(n_568),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_L g1093 ( 
.A(n_857),
.B(n_610),
.C(n_609),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_L g1094 ( 
.A(n_857),
.B(n_623),
.C(n_611),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_917),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_901),
.B(n_569),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_894),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_915),
.B(n_572),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_903),
.A2(n_484),
.B(n_482),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_921),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_922),
.B(n_485),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_922),
.B(n_488),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_919),
.B(n_492),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_770),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_924),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_927),
.B(n_575),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_928),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_929),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_932),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_918),
.B(n_493),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_791),
.B(n_579),
.Y(n_1111)
);

OR2x6_ASAP7_75t_L g1112 ( 
.A(n_930),
.B(n_591),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_930),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_770),
.B(n_580),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_770),
.B(n_581),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_847),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_859),
.B(n_495),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_871),
.B(n_586),
.Y(n_1118)
);

AO221x1_ASAP7_75t_L g1119 ( 
.A1(n_906),
.A2(n_563),
.B1(n_598),
.B2(n_603),
.C(n_592),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_859),
.B(n_497),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_910),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_850),
.Y(n_1122)
);

NOR2x1p5_ASAP7_75t_L g1123 ( 
.A(n_797),
.B(n_624),
.Y(n_1123)
);

INVxp67_ASAP7_75t_L g1124 ( 
.A(n_795),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_859),
.B(n_499),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_910),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_859),
.B(n_504),
.Y(n_1127)
);

NOR3xp33_ASAP7_75t_L g1128 ( 
.A(n_800),
.B(n_633),
.C(n_626),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_817),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_871),
.B(n_594),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_871),
.B(n_596),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_910),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_910),
.Y(n_1133)
);

AND2x6_ASAP7_75t_SL g1134 ( 
.A(n_767),
.B(n_629),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_859),
.B(n_506),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_859),
.B(n_507),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_859),
.B(n_508),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_SL g1138 ( 
.A(n_779),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_795),
.B(n_635),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_910),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_910),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_850),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_859),
.B(n_513),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_859),
.B(n_597),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_871),
.B(n_605),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_859),
.A2(n_636),
.B1(n_641),
.B2(n_631),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_871),
.B(n_606),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_795),
.B(n_639),
.Y(n_1148)
);

NOR3xp33_ASAP7_75t_L g1149 ( 
.A(n_800),
.B(n_642),
.C(n_640),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_871),
.B(n_612),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_859),
.B(n_613),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_859),
.B(n_614),
.Y(n_1152)
);

NOR2xp67_ASAP7_75t_L g1153 ( 
.A(n_797),
.B(n_26),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_779),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_779),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_859),
.B(n_537),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_871),
.B(n_621),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_871),
.B(n_628),
.Y(n_1158)
);

OR2x4_ASAP7_75t_L g1159 ( 
.A(n_947),
.B(n_650),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_963),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_972),
.B(n_647),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_981),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_981),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_981),
.B(n_632),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1139),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_971),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_982),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_933),
.A2(n_656),
.B(n_662),
.C(n_651),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_978),
.B(n_652),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1117),
.B(n_653),
.Y(n_1170)
);

OR2x6_ASAP7_75t_L g1171 ( 
.A(n_1124),
.B(n_563),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1117),
.B(n_654),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1154),
.B(n_663),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1028),
.A2(n_659),
.B1(n_544),
.B2(n_554),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_982),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1148),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1030),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_933),
.A2(n_556),
.B(n_542),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1071),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_984),
.B(n_557),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1155),
.B(n_634),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1047),
.B(n_558),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_973),
.B(n_637),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_975),
.B(n_646),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_935),
.B(n_648),
.Y(n_1185)
);

AND2x6_ASAP7_75t_L g1186 ( 
.A(n_1005),
.B(n_663),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1071),
.Y(n_1187)
);

AO22x1_ASAP7_75t_L g1188 ( 
.A1(n_974),
.A2(n_1006),
.B1(n_943),
.B2(n_935),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_SL g1189 ( 
.A(n_979),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_944),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1048),
.B(n_559),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_950),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_939),
.B(n_657),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_980),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1023),
.A2(n_1120),
.B(n_1127),
.C(n_1125),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1011),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1125),
.B(n_658),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1024),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1127),
.B(n_661),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_939),
.B(n_665),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1135),
.B(n_564),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1012),
.B(n_570),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1135),
.B(n_571),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_946),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1136),
.A2(n_585),
.B(n_590),
.C(n_577),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1122),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1142),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1119),
.A2(n_604),
.B1(n_608),
.B2(n_593),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1136),
.B(n_618),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1095),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_993),
.B(n_627),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_980),
.Y(n_1212)
);

INVx8_ASAP7_75t_L g1213 ( 
.A(n_1138),
.Y(n_1213)
);

INVx6_ASAP7_75t_L g1214 ( 
.A(n_1086),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_954),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1021),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_943),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1042),
.A2(n_638),
.B1(n_643),
.B2(n_630),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1029),
.B(n_660),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_949),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1063),
.B(n_26),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1036),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_970),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1020),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_L g1225 ( 
.A(n_958),
.B(n_547),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1138),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1037),
.Y(n_1227)
);

OA22x2_ASAP7_75t_L g1228 ( 
.A1(n_987),
.A2(n_566),
.B1(n_602),
.B2(n_599),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_985),
.A2(n_602),
.B1(n_615),
.B2(n_599),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1129),
.B(n_644),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1128),
.A2(n_547),
.B1(n_728),
.B2(n_722),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_992),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1134),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1129),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1137),
.B(n_28),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_951),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_R g1237 ( 
.A(n_1003),
.B(n_29),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1027),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_951),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1087),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_988),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_960),
.A2(n_680),
.B(n_677),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1137),
.B(n_29),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_988),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1143),
.B(n_30),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1069),
.B(n_1079),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1057),
.B(n_31),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1015),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_986),
.B(n_31),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1143),
.B(n_33),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1015),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1077),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1078),
.Y(n_1253)
);

NAND2xp33_ASAP7_75t_L g1254 ( 
.A(n_980),
.B(n_680),
.Y(n_1254)
);

NAND2xp33_ASAP7_75t_L g1255 ( 
.A(n_980),
.B(n_680),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1156),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1149),
.A2(n_734),
.B1(n_742),
.B2(n_728),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1038),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1098),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1100),
.B(n_756),
.Y(n_1260)
);

NAND2x1p5_ASAP7_75t_L g1261 ( 
.A(n_1105),
.B(n_728),
.Y(n_1261)
);

OAI21xp33_ASAP7_75t_L g1262 ( 
.A1(n_1156),
.A2(n_734),
.B(n_728),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1017),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1017),
.Y(n_1264)
);

NAND3xp33_ASAP7_75t_L g1265 ( 
.A(n_938),
.B(n_742),
.C(n_734),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1019),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_934),
.B(n_34),
.Y(n_1267)
);

INVx5_ASAP7_75t_L g1268 ( 
.A(n_1112),
.Y(n_1268)
);

BUFx2_ASAP7_75t_SL g1269 ( 
.A(n_989),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1144),
.B(n_35),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1112),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_1050),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_991),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_976),
.A2(n_742),
.B1(n_745),
.B2(n_734),
.Y(n_1274)
);

AOI22x1_ASAP7_75t_R g1275 ( 
.A1(n_1088),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1070),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1090),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1151),
.B(n_36),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1000),
.B(n_1066),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1090),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_965),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1084),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1093),
.A2(n_747),
.B1(n_756),
.B2(n_745),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_965),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_L g1285 ( 
.A(n_941),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1152),
.B(n_38),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1097),
.B(n_39),
.Y(n_1287)
);

OR2x6_ASAP7_75t_L g1288 ( 
.A(n_1123),
.B(n_745),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_997),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1094),
.A2(n_756),
.B1(n_747),
.B2(n_695),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1072),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1072),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1046),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_997),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1051),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1092),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_999),
.B(n_39),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1001),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_942),
.B(n_40),
.Y(n_1299)
);

AO22x1_ASAP7_75t_L g1300 ( 
.A1(n_1049),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_962),
.B(n_42),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1008),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1007),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_937),
.B(n_43),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1072),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1043),
.Y(n_1306)
);

OR2x2_ASAP7_75t_SL g1307 ( 
.A(n_1061),
.B(n_45),
.Y(n_1307)
);

NOR3xp33_ASAP7_75t_SL g1308 ( 
.A(n_1111),
.B(n_45),
.C(n_46),
.Y(n_1308)
);

INVx4_ASAP7_75t_L g1309 ( 
.A(n_1112),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1045),
.A2(n_756),
.B(n_747),
.C(n_695),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_999),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1118),
.B(n_46),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1146),
.B(n_48),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_966),
.B(n_48),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1005),
.B(n_747),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1054),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1065),
.Y(n_1317)
);

NOR3xp33_ASAP7_75t_SL g1318 ( 
.A(n_1033),
.B(n_49),
.C(n_50),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1081),
.Y(n_1319)
);

OR2x4_ASAP7_75t_L g1320 ( 
.A(n_994),
.B(n_50),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_941),
.Y(n_1321)
);

NOR2x1p5_ASAP7_75t_L g1322 ( 
.A(n_983),
.B(n_51),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1053),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1089),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_968),
.B(n_953),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_977),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_956),
.B(n_51),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1130),
.B(n_52),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1110),
.Y(n_1329)
);

NOR2xp67_ASAP7_75t_L g1330 ( 
.A(n_1064),
.B(n_203),
.Y(n_1330)
);

AND2x2_ASAP7_75t_SL g1331 ( 
.A(n_1062),
.B(n_52),
.Y(n_1331)
);

AND3x1_ASAP7_75t_L g1332 ( 
.A(n_1034),
.B(n_1031),
.C(n_1085),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_961),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_964),
.B(n_53),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1080),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_941),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1056),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_959),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_967),
.B(n_54),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_936),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_969),
.B(n_55),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1131),
.B(n_56),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1002),
.B(n_697),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_945),
.B(n_57),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1103),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_945),
.B(n_57),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1145),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_998),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1147),
.B(n_58),
.Y(n_1349)
);

NAND2xp33_ASAP7_75t_L g1350 ( 
.A(n_1096),
.B(n_1068),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_948),
.B(n_58),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1121),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1126),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_948),
.B(n_61),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1091),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_960),
.A2(n_210),
.B(n_204),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1132),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1009),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1099),
.A2(n_65),
.B(n_62),
.C(n_64),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1133),
.Y(n_1360)
);

BUFx4f_ASAP7_75t_L g1361 ( 
.A(n_1105),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1140),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1101),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1153),
.B(n_69),
.Y(n_1364)
);

BUFx2_ASAP7_75t_SL g1365 ( 
.A(n_995),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1141),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1103),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1150),
.B(n_71),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1102),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1010),
.Y(n_1370)
);

CKINVDCx16_ASAP7_75t_R g1371 ( 
.A(n_1018),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1074),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1016),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1052),
.Y(n_1374)
);

INVx5_ASAP7_75t_L g1375 ( 
.A(n_1076),
.Y(n_1375)
);

NAND3xp33_ASAP7_75t_SL g1376 ( 
.A(n_1013),
.B(n_1014),
.C(n_957),
.Y(n_1376)
);

AND2x6_ASAP7_75t_L g1377 ( 
.A(n_990),
.B(n_212),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1075),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_952),
.B(n_955),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1157),
.B(n_72),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1158),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1082),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1075),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1106),
.B(n_74),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1083),
.Y(n_1385)
);

INVx5_ASAP7_75t_L g1386 ( 
.A(n_1076),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1040),
.Y(n_1387)
);

CKINVDCx14_ASAP7_75t_R g1388 ( 
.A(n_1022),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1004),
.B(n_75),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1067),
.B(n_75),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_1055),
.B(n_223),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1025),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1114),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1058),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1073),
.B(n_76),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1026),
.B(n_76),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1035),
.B(n_77),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1039),
.B(n_1041),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1115),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1059),
.B(n_77),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1060),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1044),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1032),
.B(n_78),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1104),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_996),
.B(n_78),
.Y(n_1405)
);

NAND2xp33_ASAP7_75t_L g1406 ( 
.A(n_1108),
.B(n_229),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1109),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1113),
.B(n_79),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1107),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1116),
.A2(n_80),
.B(n_81),
.C(n_82),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1104),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1198),
.B(n_83),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1306),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1256),
.B(n_84),
.Y(n_1414)
);

AND2x2_ASAP7_75t_SL g1415 ( 
.A(n_1285),
.B(n_85),
.Y(n_1415)
);

NOR3xp33_ASAP7_75t_L g1416 ( 
.A(n_1188),
.B(n_87),
.C(n_88),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1226),
.B(n_88),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1345),
.B(n_1311),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1268),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1268),
.B(n_89),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1171),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1236),
.B(n_91),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1248),
.A2(n_93),
.B(n_95),
.C(n_96),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1242),
.A2(n_235),
.B(n_234),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1268),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_SL g1426 ( 
.A1(n_1304),
.A2(n_1346),
.B(n_1344),
.C(n_1389),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1178),
.A2(n_95),
.B(n_96),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1271),
.B(n_97),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1239),
.B(n_98),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1198),
.B(n_98),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1271),
.B(n_100),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1215),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1309),
.B(n_100),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1367),
.B(n_101),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1238),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1281),
.B(n_101),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1165),
.B(n_1176),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_L g1438 ( 
.A(n_1171),
.B(n_103),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1309),
.B(n_104),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1246),
.A2(n_105),
.B(n_106),
.C(n_107),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1251),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1304),
.A2(n_110),
.B(n_111),
.Y(n_1442)
);

BUFx4f_ASAP7_75t_L g1443 ( 
.A(n_1213),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1237),
.B(n_110),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1284),
.B(n_111),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1242),
.A2(n_1294),
.B(n_1289),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1205),
.A2(n_113),
.B(n_114),
.C(n_115),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1165),
.B(n_113),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1176),
.B(n_115),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1259),
.B(n_116),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1263),
.A2(n_1266),
.B(n_1264),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1277),
.B(n_117),
.Y(n_1452)
);

INVx4_ASAP7_75t_L g1453 ( 
.A(n_1213),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1223),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1265),
.B(n_117),
.C(n_118),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1280),
.B(n_118),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1338),
.B(n_119),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1190),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1192),
.B(n_120),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1213),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1217),
.B(n_121),
.Y(n_1461)
);

INVx4_ASAP7_75t_L g1462 ( 
.A(n_1171),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1206),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1166),
.B(n_121),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1207),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1245),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1232),
.B(n_1369),
.Y(n_1467)
);

NOR3xp33_ASAP7_75t_SL g1468 ( 
.A(n_1293),
.B(n_122),
.C(n_123),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1240),
.B(n_124),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1326),
.B(n_126),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1177),
.B(n_127),
.Y(n_1471)
);

BUFx4f_ASAP7_75t_L g1472 ( 
.A(n_1214),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1313),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_SL g1474 ( 
.A(n_1208),
.B(n_128),
.C(n_130),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_SL g1475 ( 
.A1(n_1344),
.A2(n_304),
.B(n_396),
.C(n_394),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1252),
.B(n_128),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_SL g1477 ( 
.A(n_1194),
.B(n_242),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1258),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1379),
.B(n_131),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1160),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1313),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1170),
.B(n_131),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1329),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1296),
.B(n_132),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1245),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1253),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1172),
.B(n_134),
.Y(n_1487)
);

AOI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1351),
.A2(n_309),
.B(n_391),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1235),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1243),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1250),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1210),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1272),
.B(n_146),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1287),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1218),
.B(n_147),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1325),
.B(n_147),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1201),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1385),
.A2(n_150),
.B(n_151),
.C(n_152),
.Y(n_1498)
);

A2O1A1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1219),
.A2(n_152),
.B(n_153),
.C(n_154),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1382),
.B(n_153),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1295),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1189),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_SL g1503 ( 
.A(n_1194),
.B(n_244),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1387),
.B(n_154),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1297),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1203),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_1506)
);

O2A1O1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1359),
.A2(n_157),
.B(n_158),
.C(n_159),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1316),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1202),
.B(n_159),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1202),
.B(n_160),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1279),
.B(n_163),
.Y(n_1511)
);

NOR3xp33_ASAP7_75t_L g1512 ( 
.A(n_1376),
.B(n_164),
.C(n_246),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1197),
.A2(n_333),
.B(n_250),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1276),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1361),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1199),
.A2(n_1209),
.B(n_1180),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1162),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1282),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1317),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1302),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1319),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1180),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1336),
.B(n_265),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1287),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1389),
.A2(n_266),
.B(n_270),
.C(n_271),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1229),
.A2(n_272),
.B1(n_273),
.B2(n_282),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1276),
.Y(n_1527)
);

A2O1A1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1221),
.A2(n_289),
.B(n_291),
.C(n_297),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1407),
.A2(n_298),
.B1(n_299),
.B2(n_302),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1288),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1392),
.B(n_1185),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_R g1532 ( 
.A(n_1321),
.B(n_308),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1233),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1183),
.A2(n_317),
.B1(n_319),
.B2(n_321),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1196),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1163),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1379),
.B(n_334),
.Y(n_1537)
);

CKINVDCx10_ASAP7_75t_R g1538 ( 
.A(n_1371),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1324),
.Y(n_1539)
);

NOR3xp33_ASAP7_75t_L g1540 ( 
.A(n_1300),
.B(n_343),
.C(n_345),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1182),
.B(n_361),
.Y(n_1541)
);

O2A1O1Ixp33_ASAP7_75t_SL g1542 ( 
.A1(n_1351),
.A2(n_367),
.B(n_368),
.C(n_370),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_SL g1543 ( 
.A(n_1194),
.B(n_373),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1229),
.A2(n_374),
.B1(n_381),
.B2(n_385),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1409),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_SL g1546 ( 
.A1(n_1354),
.A2(n_1270),
.B(n_1278),
.C(n_1286),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1402),
.B(n_1216),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1355),
.A2(n_1407),
.B1(n_1267),
.B2(n_1339),
.Y(n_1548)
);

NOR3xp33_ASAP7_75t_L g1549 ( 
.A(n_1247),
.B(n_1398),
.C(n_1312),
.Y(n_1549)
);

INVx4_ASAP7_75t_L g1550 ( 
.A(n_1167),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1222),
.B(n_1227),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1298),
.Y(n_1552)
);

NOR3xp33_ASAP7_75t_SL g1553 ( 
.A(n_1347),
.B(n_1328),
.C(n_1299),
.Y(n_1553)
);

CKINVDCx10_ASAP7_75t_R g1554 ( 
.A(n_1364),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1182),
.B(n_1191),
.Y(n_1555)
);

OAI21xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1355),
.A2(n_1228),
.B(n_1322),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1331),
.B(n_1191),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1406),
.A2(n_1327),
.B(n_1230),
.Y(n_1558)
);

INVx4_ASAP7_75t_L g1559 ( 
.A(n_1175),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1249),
.B(n_1301),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1410),
.A2(n_1397),
.B(n_1169),
.C(n_1161),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1301),
.B(n_1314),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1291),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1390),
.A2(n_1395),
.B(n_1265),
.C(n_1354),
.Y(n_1564)
);

A2O1A1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1334),
.A2(n_1330),
.B(n_1380),
.C(n_1342),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1357),
.A2(n_1360),
.B(n_1340),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1352),
.A2(n_1353),
.B(n_1362),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1341),
.B(n_1403),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_R g1569 ( 
.A(n_1285),
.B(n_1388),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1374),
.B(n_1401),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1303),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1356),
.A2(n_1305),
.B(n_1292),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1358),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1214),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1384),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1173),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1292),
.A2(n_1305),
.B(n_1405),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1384),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1403),
.B(n_1349),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1292),
.A2(n_1305),
.B(n_1330),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1335),
.A2(n_1400),
.B1(n_1396),
.B2(n_1332),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1378),
.A2(n_1383),
.B(n_1225),
.Y(n_1582)
);

BUFx8_ASAP7_75t_L g1583 ( 
.A(n_1273),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1364),
.A2(n_1307),
.B1(n_1363),
.B2(n_1320),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1396),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1368),
.A2(n_1408),
.B(n_1400),
.C(n_1231),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_SL g1587 ( 
.A(n_1181),
.B(n_1184),
.C(n_1399),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1364),
.A2(n_1212),
.B1(n_1159),
.B2(n_1333),
.Y(n_1588)
);

OAI22x1_ASAP7_75t_L g1589 ( 
.A1(n_1220),
.A2(n_1224),
.B1(n_1275),
.B2(n_1372),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1348),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1174),
.B(n_1394),
.Y(n_1591)
);

O2A1O1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1308),
.A2(n_1318),
.B(n_1288),
.C(n_1381),
.Y(n_1592)
);

NOR2xp67_ASAP7_75t_L g1593 ( 
.A(n_1393),
.B(n_1373),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1332),
.B(n_1288),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1375),
.Y(n_1595)
);

O2A1O1Ixp5_ASAP7_75t_L g1596 ( 
.A1(n_1260),
.A2(n_1343),
.B(n_1315),
.C(n_1193),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1323),
.B(n_1370),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1269),
.B(n_1365),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_R g1599 ( 
.A(n_1337),
.B(n_1186),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1254),
.A2(n_1255),
.B(n_1366),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1186),
.B(n_1244),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1186),
.B(n_1244),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1373),
.B(n_1212),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1375),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1366),
.Y(n_1605)
);

BUFx12f_ASAP7_75t_L g1606 ( 
.A(n_1186),
.Y(n_1606)
);

CKINVDCx11_ASAP7_75t_R g1607 ( 
.A(n_1241),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1164),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1404),
.A2(n_1411),
.B(n_1262),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_R g1610 ( 
.A(n_1375),
.B(n_1386),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1200),
.Y(n_1611)
);

BUFx12f_ASAP7_75t_L g1612 ( 
.A(n_1261),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1274),
.B(n_1257),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1283),
.B(n_1290),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1310),
.A2(n_1391),
.B(n_1234),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1377),
.Y(n_1616)
);

INVx4_ASAP7_75t_L g1617 ( 
.A(n_1213),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1195),
.A2(n_1256),
.B(n_1248),
.C(n_1251),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1168),
.A2(n_1195),
.B(n_1246),
.C(n_1205),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1198),
.B(n_940),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1252),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1265),
.B(n_1028),
.C(n_1211),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1204),
.Y(n_1625)
);

AND2x6_ASAP7_75t_L g1626 ( 
.A(n_1179),
.B(n_1187),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1268),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1204),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1268),
.B(n_1271),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1268),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1178),
.A2(n_933),
.B(n_945),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1345),
.B(n_940),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1198),
.B(n_940),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_R g1636 ( 
.A(n_1213),
.B(n_1226),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1268),
.B(n_1271),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1213),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1350),
.A2(n_901),
.B(n_933),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1168),
.A2(n_1195),
.B(n_1246),
.C(n_1205),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1198),
.B(n_940),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1350),
.A2(n_901),
.B(n_933),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1268),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1345),
.B(n_940),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1195),
.A2(n_1256),
.B(n_1248),
.C(n_1251),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1268),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1213),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1256),
.A2(n_1251),
.B1(n_1248),
.B2(n_1239),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1268),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1268),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1198),
.B(n_940),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1268),
.B(n_1271),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1178),
.A2(n_933),
.B(n_945),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_SL g1657 ( 
.A(n_1238),
.B(n_780),
.C(n_778),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1252),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_SL g1659 ( 
.A(n_1238),
.B(n_780),
.C(n_778),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1198),
.B(n_940),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1661)
);

BUFx3_ASAP7_75t_L g1662 ( 
.A(n_1213),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1198),
.A2(n_1028),
.B1(n_906),
.B2(n_868),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1198),
.B(n_940),
.Y(n_1664)
);

AND2x2_ASAP7_75t_SL g1665 ( 
.A(n_1285),
.B(n_1003),
.Y(n_1665)
);

CKINVDCx16_ASAP7_75t_R g1666 ( 
.A(n_1171),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1443),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1443),
.Y(n_1668)
);

INVx4_ASAP7_75t_L g1669 ( 
.A(n_1453),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1634),
.B(n_1644),
.Y(n_1670)
);

NAND2x1p5_ASAP7_75t_L g1671 ( 
.A(n_1453),
.B(n_1617),
.Y(n_1671)
);

AO21x2_ASAP7_75t_L g1672 ( 
.A1(n_1426),
.A2(n_1564),
.B(n_1546),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1610),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1604),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1612),
.Y(n_1675)
);

INVx6_ASAP7_75t_L g1676 ( 
.A(n_1617),
.Y(n_1676)
);

BUFx2_ASAP7_75t_SL g1677 ( 
.A(n_1502),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1418),
.B(n_1618),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1572),
.A2(n_1577),
.B(n_1580),
.Y(n_1679)
);

OAI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1609),
.A2(n_1615),
.B(n_1488),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1568),
.B(n_1562),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1624),
.Y(n_1682)
);

BUFx2_ASAP7_75t_SL g1683 ( 
.A(n_1662),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1631),
.B(n_1632),
.Y(n_1684)
);

AO21x1_ASAP7_75t_L g1685 ( 
.A1(n_1584),
.A2(n_1529),
.B(n_1526),
.Y(n_1685)
);

INVx6_ASAP7_75t_L g1686 ( 
.A(n_1583),
.Y(n_1686)
);

AO21x2_ASAP7_75t_L g1687 ( 
.A1(n_1633),
.A2(n_1656),
.B(n_1639),
.Y(n_1687)
);

AO21x2_ASAP7_75t_L g1688 ( 
.A1(n_1633),
.A2(n_1656),
.B(n_1642),
.Y(n_1688)
);

INVx4_ASAP7_75t_L g1689 ( 
.A(n_1460),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1607),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1619),
.A2(n_1645),
.B(n_1516),
.Y(n_1691)
);

INVx6_ASAP7_75t_SL g1692 ( 
.A(n_1570),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1606),
.Y(n_1693)
);

OAI21x1_ASAP7_75t_SL g1694 ( 
.A1(n_1650),
.A2(n_1442),
.B(n_1588),
.Y(n_1694)
);

NAND2x1p5_ASAP7_75t_L g1695 ( 
.A(n_1629),
.B(n_1637),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1584),
.A2(n_1415),
.B1(n_1650),
.B2(n_1665),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1636),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1646),
.B(n_1649),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1595),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1652),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1554),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_SL g1702 ( 
.A1(n_1442),
.A2(n_1588),
.B(n_1427),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1437),
.Y(n_1703)
);

OR2x6_ASAP7_75t_L g1704 ( 
.A(n_1462),
.B(n_1638),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1661),
.Y(n_1705)
);

OAI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1446),
.A2(n_1451),
.B(n_1485),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1522),
.B(n_1473),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1413),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1582),
.A2(n_1600),
.B(n_1424),
.Y(n_1709)
);

INVx4_ASAP7_75t_L g1710 ( 
.A(n_1486),
.Y(n_1710)
);

INVx3_ASAP7_75t_SL g1711 ( 
.A(n_1666),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1481),
.B(n_1467),
.Y(n_1712)
);

BUFx12f_ASAP7_75t_L g1713 ( 
.A(n_1583),
.Y(n_1713)
);

INVx5_ASAP7_75t_SL g1714 ( 
.A(n_1616),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1489),
.B(n_1458),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1538),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1530),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1575),
.B(n_1578),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1463),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1472),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1585),
.B(n_1419),
.Y(n_1721)
);

BUFx2_ASAP7_75t_SL g1722 ( 
.A(n_1648),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1432),
.Y(n_1723)
);

INVx8_ASAP7_75t_L g1724 ( 
.A(n_1626),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1512),
.B(n_1623),
.C(n_1416),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1454),
.Y(n_1726)
);

INVx6_ASAP7_75t_L g1727 ( 
.A(n_1517),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1472),
.Y(n_1728)
);

NAND2x1p5_ASAP7_75t_L g1729 ( 
.A(n_1655),
.B(n_1419),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1505),
.B(n_1548),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1552),
.Y(n_1731)
);

BUFx4f_ASAP7_75t_L g1732 ( 
.A(n_1435),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1571),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1595),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1620),
.A2(n_1640),
.B(n_1548),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1478),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1425),
.B(n_1643),
.Y(n_1737)
);

AO21x2_ASAP7_75t_L g1738 ( 
.A1(n_1455),
.A2(n_1565),
.B(n_1542),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1664),
.B(n_1621),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1425),
.B(n_1643),
.Y(n_1740)
);

INVx8_ASAP7_75t_L g1741 ( 
.A(n_1626),
.Y(n_1741)
);

NAND2x1p5_ASAP7_75t_L g1742 ( 
.A(n_1647),
.B(n_1517),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1635),
.B(n_1641),
.Y(n_1743)
);

BUFx2_ASAP7_75t_SL g1744 ( 
.A(n_1535),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1479),
.Y(n_1745)
);

BUFx12f_ASAP7_75t_L g1746 ( 
.A(n_1518),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1579),
.B(n_1555),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1560),
.B(n_1496),
.Y(n_1748)
);

AO21x2_ASAP7_75t_L g1749 ( 
.A1(n_1586),
.A2(n_1623),
.B(n_1475),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_1599),
.Y(n_1750)
);

OAI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1561),
.A2(n_1556),
.B(n_1456),
.Y(n_1751)
);

INVx4_ASAP7_75t_L g1752 ( 
.A(n_1514),
.Y(n_1752)
);

BUFx12f_ASAP7_75t_L g1753 ( 
.A(n_1574),
.Y(n_1753)
);

OAI21x1_ASAP7_75t_L g1754 ( 
.A1(n_1601),
.A2(n_1602),
.B(n_1596),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1479),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1471),
.Y(n_1756)
);

AO21x2_ASAP7_75t_L g1757 ( 
.A1(n_1540),
.A2(n_1525),
.B(n_1614),
.Y(n_1757)
);

INVx6_ASAP7_75t_L g1758 ( 
.A(n_1536),
.Y(n_1758)
);

NAND2x1p5_ASAP7_75t_L g1759 ( 
.A(n_1536),
.B(n_1550),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1550),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1559),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1452),
.A2(n_1429),
.B(n_1422),
.Y(n_1762)
);

INVx5_ASAP7_75t_L g1763 ( 
.A(n_1527),
.Y(n_1763)
);

BUFx4f_ASAP7_75t_L g1764 ( 
.A(n_1616),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1654),
.B(n_1660),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1414),
.A2(n_1445),
.B(n_1436),
.Y(n_1766)
);

AO21x2_ASAP7_75t_L g1767 ( 
.A1(n_1528),
.A2(n_1459),
.B(n_1482),
.Y(n_1767)
);

BUFx4f_ASAP7_75t_L g1768 ( 
.A(n_1524),
.Y(n_1768)
);

INVx4_ASAP7_75t_L g1769 ( 
.A(n_1559),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1504),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1434),
.A2(n_1507),
.B(n_1566),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1511),
.B(n_1549),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1622),
.B(n_1658),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1545),
.Y(n_1774)
);

CKINVDCx16_ASAP7_75t_R g1775 ( 
.A(n_1569),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1487),
.A2(n_1567),
.B(n_1495),
.Y(n_1776)
);

BUFx12f_ASAP7_75t_L g1777 ( 
.A(n_1608),
.Y(n_1777)
);

OR2x6_ASAP7_75t_L g1778 ( 
.A(n_1515),
.B(n_1494),
.Y(n_1778)
);

BUFx8_ASAP7_75t_L g1779 ( 
.A(n_1570),
.Y(n_1779)
);

AO21x2_ASAP7_75t_L g1780 ( 
.A1(n_1474),
.A2(n_1544),
.B(n_1423),
.Y(n_1780)
);

NOR2xp67_ASAP7_75t_SL g1781 ( 
.A(n_1576),
.B(n_1627),
.Y(n_1781)
);

OAI21x1_ASAP7_75t_SL g1782 ( 
.A1(n_1466),
.A2(n_1592),
.B(n_1497),
.Y(n_1782)
);

AO21x2_ASAP7_75t_L g1783 ( 
.A1(n_1509),
.A2(n_1510),
.B(n_1498),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1663),
.A2(n_1557),
.B1(n_1594),
.B2(n_1421),
.Y(n_1784)
);

NOR2x1_ASAP7_75t_L g1785 ( 
.A(n_1438),
.B(n_1417),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1447),
.A2(n_1613),
.B(n_1537),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1625),
.B(n_1628),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1591),
.B(n_1531),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1630),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1581),
.B(n_1547),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1626),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1480),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1493),
.B(n_1470),
.Y(n_1793)
);

INVxp67_ASAP7_75t_SL g1794 ( 
.A(n_1563),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1603),
.B(n_1492),
.Y(n_1795)
);

OAI21x1_ASAP7_75t_L g1796 ( 
.A1(n_1590),
.A2(n_1521),
.B(n_1539),
.Y(n_1796)
);

OAI22x1_ASAP7_75t_L g1797 ( 
.A1(n_1444),
.A2(n_1412),
.B1(n_1430),
.B2(n_1476),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1497),
.Y(n_1798)
);

AO21x2_ASAP7_75t_L g1799 ( 
.A1(n_1541),
.A2(n_1534),
.B(n_1499),
.Y(n_1799)
);

OR2x6_ASAP7_75t_L g1800 ( 
.A(n_1533),
.B(n_1598),
.Y(n_1800)
);

AO21x2_ASAP7_75t_L g1801 ( 
.A1(n_1420),
.A2(n_1428),
.B(n_1431),
.Y(n_1801)
);

OA21x2_ASAP7_75t_L g1802 ( 
.A1(n_1433),
.A2(n_1439),
.B(n_1520),
.Y(n_1802)
);

INVx6_ASAP7_75t_L g1803 ( 
.A(n_1603),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1651),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1448),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1657),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1466),
.Y(n_1807)
);

AO21x2_ASAP7_75t_L g1808 ( 
.A1(n_1490),
.A2(n_1491),
.B(n_1440),
.Y(n_1808)
);

AO21x2_ASAP7_75t_L g1809 ( 
.A1(n_1490),
.A2(n_1491),
.B(n_1500),
.Y(n_1809)
);

BUFx2_ASAP7_75t_SL g1810 ( 
.A(n_1653),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1457),
.B(n_1450),
.Y(n_1811)
);

OAI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1501),
.A2(n_1508),
.B(n_1519),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1484),
.B(n_1469),
.Y(n_1813)
);

OR2x6_ASAP7_75t_L g1814 ( 
.A(n_1573),
.B(n_1593),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1553),
.B(n_1605),
.Y(n_1815)
);

OAI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1611),
.A2(n_1573),
.B(n_1483),
.Y(n_1816)
);

OAI21x1_ASAP7_75t_L g1817 ( 
.A1(n_1441),
.A2(n_1506),
.B(n_1464),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1449),
.A2(n_1461),
.B(n_1523),
.Y(n_1818)
);

INVx5_ASAP7_75t_L g1819 ( 
.A(n_1477),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1477),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1503),
.Y(n_1821)
);

NAND2x1p5_ASAP7_75t_L g1822 ( 
.A(n_1551),
.B(n_1597),
.Y(n_1822)
);

AOI22x1_ASAP7_75t_L g1823 ( 
.A1(n_1543),
.A2(n_1587),
.B1(n_1468),
.B2(n_1532),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1659),
.Y(n_1824)
);

AOI22x1_ASAP7_75t_L g1825 ( 
.A1(n_1516),
.A2(n_1558),
.B1(n_1589),
.B2(n_1513),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1618),
.Y(n_1826)
);

OAI21x1_ASAP7_75t_L g1827 ( 
.A1(n_1572),
.A2(n_1577),
.B(n_1580),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1568),
.B(n_1562),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1572),
.A2(n_1577),
.B(n_1580),
.Y(n_1829)
);

NOR2xp67_ASAP7_75t_R g1830 ( 
.A(n_1606),
.B(n_1616),
.Y(n_1830)
);

BUFx3_ASAP7_75t_L g1831 ( 
.A(n_1443),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1522),
.B(n_1256),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1618),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1443),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1616),
.B(n_1650),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1618),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1443),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1465),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1618),
.Y(n_1839)
);

INVxp67_ASAP7_75t_SL g1840 ( 
.A(n_1650),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1618),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1708),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1730),
.Y(n_1843)
);

INVx5_ASAP7_75t_L g1844 ( 
.A(n_1713),
.Y(n_1844)
);

INVx6_ASAP7_75t_L g1845 ( 
.A(n_1675),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1675),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1705),
.Y(n_1847)
);

NOR2xp67_ASAP7_75t_L g1848 ( 
.A(n_1669),
.B(n_1701),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1705),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1730),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1707),
.Y(n_1851)
);

INVx6_ASAP7_75t_L g1852 ( 
.A(n_1686),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1684),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1707),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1686),
.Y(n_1855)
);

BUFx2_ASAP7_75t_R g1856 ( 
.A(n_1716),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1696),
.A2(n_1685),
.B1(n_1790),
.B2(n_1784),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1736),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1838),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1686),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1696),
.A2(n_1790),
.B1(n_1784),
.B2(n_1694),
.Y(n_1861)
);

OAI21x1_ASAP7_75t_L g1862 ( 
.A1(n_1679),
.A2(n_1829),
.B(n_1827),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1669),
.Y(n_1863)
);

AO21x1_ASAP7_75t_SL g1864 ( 
.A1(n_1745),
.A2(n_1755),
.B(n_1819),
.Y(n_1864)
);

BUFx3_ASAP7_75t_L g1865 ( 
.A(n_1673),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1788),
.A2(n_1782),
.B1(n_1702),
.B2(n_1811),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1840),
.A2(n_1682),
.B1(n_1826),
.B2(n_1755),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_SL g1868 ( 
.A1(n_1745),
.A2(n_1823),
.B1(n_1840),
.B2(n_1819),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1739),
.A2(n_1743),
.B1(n_1765),
.B2(n_1772),
.Y(n_1869)
);

CKINVDCx11_ASAP7_75t_R g1870 ( 
.A(n_1697),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1787),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1819),
.A2(n_1770),
.B1(n_1698),
.B2(n_1678),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_SL g1873 ( 
.A1(n_1820),
.A2(n_1821),
.B1(n_1770),
.B2(n_1768),
.Y(n_1873)
);

BUFx8_ASAP7_75t_L g1874 ( 
.A(n_1690),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1810),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_SL g1876 ( 
.A1(n_1820),
.A2(n_1768),
.B1(n_1703),
.B2(n_1741),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1671),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1676),
.Y(n_1878)
);

BUFx12f_ASAP7_75t_L g1879 ( 
.A(n_1716),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1832),
.A2(n_1712),
.B1(n_1772),
.B2(n_1805),
.Y(n_1880)
);

AO21x2_ASAP7_75t_L g1881 ( 
.A1(n_1735),
.A2(n_1691),
.B(n_1749),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1813),
.A2(n_1798),
.B1(n_1807),
.B2(n_1793),
.Y(n_1882)
);

OR2x6_ASAP7_75t_L g1883 ( 
.A(n_1677),
.B(n_1683),
.Y(n_1883)
);

INVx4_ASAP7_75t_SL g1884 ( 
.A(n_1711),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1670),
.B(n_1700),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1719),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1731),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1779),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1676),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1813),
.A2(n_1747),
.B1(n_1681),
.B2(n_1828),
.Y(n_1890)
);

AOI21x1_ASAP7_75t_L g1891 ( 
.A1(n_1835),
.A2(n_1680),
.B(n_1709),
.Y(n_1891)
);

AOI21x1_ASAP7_75t_L g1892 ( 
.A1(n_1835),
.A2(n_1735),
.B(n_1691),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1748),
.A2(n_1805),
.B1(n_1747),
.B2(n_1809),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1748),
.A2(n_1809),
.B1(n_1681),
.B2(n_1828),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1787),
.Y(n_1895)
);

INVx2_ASAP7_75t_SL g1896 ( 
.A(n_1676),
.Y(n_1896)
);

NAND2x1p5_ASAP7_75t_L g1897 ( 
.A(n_1668),
.B(n_1831),
.Y(n_1897)
);

NAND2x1p5_ASAP7_75t_L g1898 ( 
.A(n_1668),
.B(n_1831),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1733),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1833),
.B(n_1836),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1723),
.Y(n_1901)
);

BUFx4f_ASAP7_75t_L g1902 ( 
.A(n_1711),
.Y(n_1902)
);

INVx6_ASAP7_75t_L g1903 ( 
.A(n_1779),
.Y(n_1903)
);

BUFx2_ASAP7_75t_L g1904 ( 
.A(n_1692),
.Y(n_1904)
);

INVx4_ASAP7_75t_L g1905 ( 
.A(n_1834),
.Y(n_1905)
);

CKINVDCx11_ASAP7_75t_R g1906 ( 
.A(n_1697),
.Y(n_1906)
);

INVx6_ASAP7_75t_L g1907 ( 
.A(n_1753),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1726),
.Y(n_1908)
);

AO21x1_ASAP7_75t_L g1909 ( 
.A1(n_1751),
.A2(n_1786),
.B(n_1706),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1832),
.A2(n_1703),
.B1(n_1839),
.B2(n_1841),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_1750),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1706),
.Y(n_1912)
);

BUFx10_ASAP7_75t_L g1913 ( 
.A(n_1667),
.Y(n_1913)
);

BUFx2_ASAP7_75t_L g1914 ( 
.A(n_1692),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1715),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1715),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1812),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1774),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1796),
.Y(n_1919)
);

OAI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1775),
.A2(n_1800),
.B1(n_1822),
.B2(n_1773),
.Y(n_1920)
);

OAI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1800),
.A2(n_1750),
.B1(n_1792),
.B2(n_1704),
.Y(n_1921)
);

CKINVDCx11_ASAP7_75t_R g1922 ( 
.A(n_1710),
.Y(n_1922)
);

INVx4_ASAP7_75t_L g1923 ( 
.A(n_1834),
.Y(n_1923)
);

BUFx2_ASAP7_75t_SL g1924 ( 
.A(n_1837),
.Y(n_1924)
);

INVx8_ASAP7_75t_L g1925 ( 
.A(n_1746),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1789),
.B(n_1804),
.Y(n_1926)
);

AOI21xp33_ASAP7_75t_L g1927 ( 
.A1(n_1725),
.A2(n_1751),
.B(n_1825),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1718),
.Y(n_1928)
);

BUFx12f_ASAP7_75t_L g1929 ( 
.A(n_1710),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1724),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1815),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1789),
.Y(n_1932)
);

INVx3_ASAP7_75t_L g1933 ( 
.A(n_1724),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1815),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1754),
.Y(n_1935)
);

BUFx2_ASAP7_75t_R g1936 ( 
.A(n_1806),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1785),
.B(n_1704),
.Y(n_1937)
);

INVx3_ASAP7_75t_L g1938 ( 
.A(n_1724),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1741),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1672),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1804),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1756),
.A2(n_1797),
.B1(n_1818),
.B2(n_1808),
.Y(n_1942)
);

BUFx2_ASAP7_75t_R g1943 ( 
.A(n_1806),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1744),
.Y(n_1944)
);

OAI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1818),
.A2(n_1800),
.B1(n_1704),
.B2(n_1717),
.Y(n_1945)
);

BUFx2_ASAP7_75t_L g1946 ( 
.A(n_1837),
.Y(n_1946)
);

OR2x6_ASAP7_75t_L g1947 ( 
.A(n_1741),
.B(n_1690),
.Y(n_1947)
);

INVx8_ASAP7_75t_L g1948 ( 
.A(n_1777),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1687),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1808),
.A2(n_1780),
.B1(n_1783),
.B2(n_1766),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1687),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1732),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1844),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1920),
.B(n_1769),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1883),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1843),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1900),
.B(n_1795),
.Y(n_1957)
);

OAI21xp5_ASAP7_75t_SL g1958 ( 
.A1(n_1888),
.A2(n_1824),
.B(n_1791),
.Y(n_1958)
);

NAND2xp33_ASAP7_75t_R g1959 ( 
.A(n_1883),
.B(n_1863),
.Y(n_1959)
);

INVx6_ASAP7_75t_L g1960 ( 
.A(n_1844),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1885),
.B(n_1795),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_R g1962 ( 
.A(n_1844),
.B(n_1732),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1857),
.A2(n_1814),
.B1(n_1778),
.B2(n_1742),
.Y(n_1963)
);

INVxp33_ASAP7_75t_L g1964 ( 
.A(n_1848),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1926),
.B(n_1737),
.Y(n_1965)
);

OR2x6_ASAP7_75t_L g1966 ( 
.A(n_1925),
.B(n_1722),
.Y(n_1966)
);

OR2x6_ASAP7_75t_L g1967 ( 
.A(n_1925),
.B(n_1693),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1869),
.B(n_1721),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1922),
.Y(n_1969)
);

NAND2xp33_ASAP7_75t_R g1970 ( 
.A(n_1863),
.B(n_1814),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1847),
.Y(n_1971)
);

O2A1O1Ixp33_ASAP7_75t_L g1972 ( 
.A1(n_1880),
.A2(n_1762),
.B(n_1766),
.C(n_1778),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1915),
.B(n_1916),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1843),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1850),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1932),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1877),
.B(n_1769),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1929),
.Y(n_1978)
);

NAND2xp33_ASAP7_75t_R g1979 ( 
.A(n_1877),
.B(n_1814),
.Y(n_1979)
);

BUFx4f_ASAP7_75t_SL g1980 ( 
.A(n_1879),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_SL g1981 ( 
.A(n_1875),
.B(n_1689),
.C(n_1742),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1859),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1870),
.Y(n_1983)
);

HB1xp67_ASAP7_75t_L g1984 ( 
.A(n_1849),
.Y(n_1984)
);

OAI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1942),
.A2(n_1817),
.B(n_1816),
.Y(n_1985)
);

BUFx3_ASAP7_75t_L g1986 ( 
.A(n_1845),
.Y(n_1986)
);

BUFx8_ASAP7_75t_L g1987 ( 
.A(n_1952),
.Y(n_1987)
);

CKINVDCx16_ASAP7_75t_R g1988 ( 
.A(n_1911),
.Y(n_1988)
);

NAND3xp33_ASAP7_75t_SL g1989 ( 
.A(n_1846),
.B(n_1689),
.C(n_1729),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_R g1990 ( 
.A(n_1903),
.B(n_1720),
.Y(n_1990)
);

NOR3xp33_ASAP7_75t_SL g1991 ( 
.A(n_1921),
.B(n_1762),
.C(n_1776),
.Y(n_1991)
);

CKINVDCx11_ASAP7_75t_R g1992 ( 
.A(n_1906),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1851),
.B(n_1760),
.Y(n_1993)
);

AO31x2_ASAP7_75t_L g1994 ( 
.A1(n_1909),
.A2(n_1752),
.A3(n_1749),
.B(n_1738),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1915),
.B(n_1737),
.Y(n_1995)
);

OR2x2_ASAP7_75t_SL g1996 ( 
.A(n_1903),
.B(n_1802),
.Y(n_1996)
);

NAND2xp33_ASAP7_75t_R g1997 ( 
.A(n_1947),
.B(n_1761),
.Y(n_1997)
);

CKINVDCx16_ASAP7_75t_R g1998 ( 
.A(n_1947),
.Y(n_1998)
);

AOI221xp5_ASAP7_75t_L g1999 ( 
.A1(n_1910),
.A2(n_1776),
.B1(n_1781),
.B2(n_1771),
.C(n_1740),
.Y(n_1999)
);

CKINVDCx20_ASAP7_75t_R g2000 ( 
.A(n_1874),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1853),
.Y(n_2001)
);

CKINVDCx8_ASAP7_75t_R g2002 ( 
.A(n_1884),
.Y(n_2002)
);

AOI21xp33_ASAP7_75t_L g2003 ( 
.A1(n_1893),
.A2(n_1801),
.B(n_1802),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1927),
.A2(n_1794),
.B(n_1771),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1845),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_R g2006 ( 
.A(n_1902),
.B(n_1728),
.Y(n_2006)
);

NAND3xp33_ASAP7_75t_SL g2007 ( 
.A(n_1890),
.B(n_1729),
.C(n_1695),
.Y(n_2007)
);

NOR2xp67_ASAP7_75t_R g2008 ( 
.A(n_1852),
.B(n_1693),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1854),
.B(n_1761),
.Y(n_2009)
);

NAND2xp33_ASAP7_75t_R g2010 ( 
.A(n_1946),
.B(n_1740),
.Y(n_2010)
);

OAI21xp33_ASAP7_75t_L g2011 ( 
.A1(n_1861),
.A2(n_1950),
.B(n_1866),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1931),
.A2(n_1780),
.B1(n_1799),
.B2(n_1801),
.Y(n_2012)
);

OR2x6_ASAP7_75t_L g2013 ( 
.A(n_1948),
.B(n_1803),
.Y(n_2013)
);

NOR3xp33_ASAP7_75t_SL g2014 ( 
.A(n_1945),
.B(n_1830),
.C(n_1794),
.Y(n_2014)
);

AO21x1_ASAP7_75t_L g2015 ( 
.A1(n_1872),
.A2(n_1695),
.B(n_1759),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1934),
.A2(n_1799),
.B1(n_1767),
.B2(n_1757),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_R g2017 ( 
.A(n_1904),
.B(n_1674),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1941),
.B(n_1918),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1899),
.Y(n_2019)
);

NAND2x1p5_ASAP7_75t_L g2020 ( 
.A(n_1902),
.B(n_1763),
.Y(n_2020)
);

OAI21x1_ASAP7_75t_SL g2021 ( 
.A1(n_1937),
.A2(n_1752),
.B(n_1714),
.Y(n_2021)
);

CKINVDCx8_ASAP7_75t_R g2022 ( 
.A(n_1884),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1854),
.B(n_1882),
.Y(n_2023)
);

NAND2xp33_ASAP7_75t_R g2024 ( 
.A(n_1914),
.B(n_1734),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1899),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1856),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_R g2027 ( 
.A(n_1948),
.B(n_1764),
.Y(n_2027)
);

INVx3_ASAP7_75t_SL g2028 ( 
.A(n_1907),
.Y(n_2028)
);

NOR3xp33_ASAP7_75t_SL g2029 ( 
.A(n_1874),
.B(n_1803),
.C(n_1727),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1901),
.Y(n_2030)
);

NAND2xp33_ASAP7_75t_R g2031 ( 
.A(n_1930),
.B(n_1933),
.Y(n_2031)
);

BUFx2_ASAP7_75t_R g2032 ( 
.A(n_1924),
.Y(n_2032)
);

NOR3xp33_ASAP7_75t_SL g2033 ( 
.A(n_1867),
.B(n_1727),
.C(n_1758),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1907),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1858),
.Y(n_2035)
);

AND2x6_ASAP7_75t_L g2036 ( 
.A(n_1864),
.B(n_1714),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1949),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_2010),
.A2(n_1894),
.B1(n_1895),
.B2(n_1871),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2037),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2018),
.B(n_1901),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2023),
.B(n_1908),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1956),
.B(n_1881),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_2037),
.B(n_1949),
.Y(n_2043)
);

INVx2_ASAP7_75t_SL g2044 ( 
.A(n_1960),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1956),
.B(n_1881),
.Y(n_2045)
);

CKINVDCx14_ASAP7_75t_R g2046 ( 
.A(n_2000),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1974),
.B(n_1912),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1975),
.B(n_1912),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_2019),
.B(n_1951),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_2025),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2030),
.B(n_1951),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2035),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_L g2053 ( 
.A1(n_2011),
.A2(n_1868),
.B1(n_1873),
.B2(n_1928),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2012),
.B(n_1892),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1971),
.B(n_1908),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2016),
.B(n_1940),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1985),
.B(n_1982),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_1959),
.Y(n_2058)
);

BUFx2_ASAP7_75t_L g2059 ( 
.A(n_1996),
.Y(n_2059)
);

INVx2_ASAP7_75t_SL g2060 ( 
.A(n_1960),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1994),
.B(n_1862),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1984),
.B(n_2001),
.Y(n_2062)
);

OAI221xp5_ASAP7_75t_L g2063 ( 
.A1(n_1991),
.A2(n_1876),
.B1(n_1944),
.B2(n_1860),
.C(n_1855),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_1976),
.B(n_1842),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1973),
.Y(n_2065)
);

INVx8_ASAP7_75t_L g2066 ( 
.A(n_2036),
.Y(n_2066)
);

INVx5_ASAP7_75t_SL g2067 ( 
.A(n_1966),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_1970),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1965),
.B(n_1917),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_2032),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1995),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_2036),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1993),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1993),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_2009),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_1957),
.B(n_1886),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2003),
.B(n_1919),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2043),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2071),
.B(n_1972),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2069),
.B(n_1935),
.Y(n_2080)
);

BUFx2_ASAP7_75t_L g2081 ( 
.A(n_2059),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2043),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2071),
.B(n_1887),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_2059),
.B(n_2014),
.Y(n_2084)
);

NAND3xp33_ASAP7_75t_L g2085 ( 
.A(n_2053),
.B(n_2063),
.C(n_2038),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2039),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2069),
.B(n_2042),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2042),
.B(n_1935),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2043),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2045),
.B(n_1919),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_2061),
.B(n_1891),
.Y(n_2091)
);

NAND3xp33_ASAP7_75t_L g2092 ( 
.A(n_2038),
.B(n_1999),
.C(n_2033),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2045),
.B(n_2004),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2055),
.B(n_1968),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2057),
.B(n_1688),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2057),
.B(n_2049),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_2066),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2065),
.B(n_2009),
.Y(n_2098)
);

INVx2_ASAP7_75t_SL g2099 ( 
.A(n_2066),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_2055),
.B(n_1688),
.Y(n_2100)
);

NAND2x1p5_ASAP7_75t_L g2101 ( 
.A(n_2072),
.B(n_1954),
.Y(n_2101)
);

NAND2x1_ASAP7_75t_SL g2102 ( 
.A(n_2072),
.B(n_1977),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2050),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2065),
.B(n_1961),
.Y(n_2104)
);

NAND4xp25_ASAP7_75t_L g2105 ( 
.A(n_2058),
.B(n_2062),
.C(n_2041),
.D(n_1963),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2040),
.B(n_2076),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2096),
.B(n_2077),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2096),
.B(n_2087),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2103),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2093),
.B(n_2052),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2086),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2086),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_2091),
.Y(n_2113)
);

AOI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_2085),
.A2(n_2068),
.B(n_1962),
.C(n_1981),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2087),
.B(n_2077),
.Y(n_2115)
);

AOI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_2092),
.A2(n_2007),
.B1(n_2074),
.B2(n_2073),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2093),
.B(n_2054),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2090),
.B(n_2052),
.Y(n_2118)
);

INVxp67_ASAP7_75t_SL g2119 ( 
.A(n_2081),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2094),
.B(n_2064),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2081),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2095),
.B(n_2054),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2090),
.B(n_2051),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2095),
.B(n_2056),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2078),
.B(n_2056),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2094),
.B(n_2064),
.Y(n_2126)
);

INVxp67_ASAP7_75t_L g2127 ( 
.A(n_2105),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2078),
.B(n_2047),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2082),
.B(n_2047),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2082),
.B(n_2048),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2118),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_2110),
.B(n_2123),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2118),
.Y(n_2133)
);

INVxp67_ASAP7_75t_L g2134 ( 
.A(n_2121),
.Y(n_2134)
);

INVx3_ASAP7_75t_SL g2135 ( 
.A(n_2120),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2117),
.B(n_2088),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2107),
.B(n_2084),
.Y(n_2137)
);

NAND2x1_ASAP7_75t_SL g2138 ( 
.A(n_2113),
.B(n_2084),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2110),
.Y(n_2139)
);

O2A1O1Ixp33_ASAP7_75t_SL g2140 ( 
.A1(n_2114),
.A2(n_2070),
.B(n_2099),
.C(n_2097),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2117),
.B(n_2088),
.Y(n_2141)
);

INVxp67_ASAP7_75t_SL g2142 ( 
.A(n_2119),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2120),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2127),
.A2(n_2079),
.B1(n_2084),
.B2(n_2098),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_2114),
.A2(n_1998),
.B1(n_2106),
.B2(n_2080),
.Y(n_2145)
);

OAI211xp5_ASAP7_75t_SL g2146 ( 
.A1(n_2116),
.A2(n_1992),
.B(n_2046),
.C(n_2022),
.Y(n_2146)
);

A2O1A1Ixp33_ASAP7_75t_L g2147 ( 
.A1(n_2113),
.A2(n_2102),
.B(n_1955),
.C(n_1964),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2109),
.Y(n_2148)
);

AOI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_2122),
.A2(n_2080),
.B1(n_2097),
.B2(n_2099),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2126),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2109),
.Y(n_2151)
);

AOI211xp5_ASAP7_75t_L g2152 ( 
.A1(n_2113),
.A2(n_2028),
.B(n_1953),
.C(n_1958),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2126),
.Y(n_2153)
);

XNOR2x2_ASAP7_75t_L g2154 ( 
.A(n_2108),
.B(n_1989),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2122),
.B(n_2100),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2107),
.B(n_2089),
.Y(n_2156)
);

AOI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_2140),
.A2(n_2101),
.B(n_2066),
.Y(n_2157)
);

INVxp67_ASAP7_75t_SL g2158 ( 
.A(n_2142),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2143),
.Y(n_2159)
);

NOR3xp33_ASAP7_75t_L g2160 ( 
.A(n_2146),
.B(n_1988),
.C(n_2113),
.Y(n_2160)
);

NAND3xp33_ASAP7_75t_SL g2161 ( 
.A(n_2152),
.B(n_2002),
.C(n_2101),
.Y(n_2161)
);

INVxp67_ASAP7_75t_L g2162 ( 
.A(n_2154),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2150),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2135),
.Y(n_2164)
);

NOR2x1_ASAP7_75t_L g2165 ( 
.A(n_2146),
.B(n_1966),
.Y(n_2165)
);

OAI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2145),
.A2(n_2101),
.B1(n_2067),
.B2(n_2123),
.Y(n_2166)
);

INVx1_ASAP7_75t_SL g2167 ( 
.A(n_2138),
.Y(n_2167)
);

INVxp67_ASAP7_75t_L g2168 ( 
.A(n_2144),
.Y(n_2168)
);

OAI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_2134),
.A2(n_2102),
.B(n_2060),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2139),
.B(n_2124),
.Y(n_2170)
);

OAI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_2149),
.A2(n_2072),
.B1(n_2066),
.B2(n_2075),
.Y(n_2171)
);

NAND3xp33_ASAP7_75t_L g2172 ( 
.A(n_2134),
.B(n_2112),
.C(n_2111),
.Y(n_2172)
);

AOI22xp33_ASAP7_75t_L g2173 ( 
.A1(n_2162),
.A2(n_2153),
.B1(n_2067),
.B2(n_2074),
.Y(n_2173)
);

AO21x1_ASAP7_75t_L g2174 ( 
.A1(n_2158),
.A2(n_2024),
.B(n_1997),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_SL g2175 ( 
.A(n_2165),
.B(n_2026),
.Y(n_2175)
);

NAND3x2_ASAP7_75t_L g2176 ( 
.A(n_2160),
.B(n_2137),
.C(n_2159),
.Y(n_2176)
);

OAI21xp33_ASAP7_75t_L g2177 ( 
.A1(n_2168),
.A2(n_2133),
.B(n_2131),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2164),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2163),
.Y(n_2179)
);

OAI321xp33_ASAP7_75t_L g2180 ( 
.A1(n_2166),
.A2(n_2147),
.A3(n_2044),
.B1(n_2060),
.B2(n_2155),
.C(n_2100),
.Y(n_2180)
);

INVxp67_ASAP7_75t_L g2181 ( 
.A(n_2172),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2167),
.B(n_2108),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2170),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2169),
.B(n_2155),
.Y(n_2184)
);

AOI322xp5_ASAP7_75t_L g2185 ( 
.A1(n_2161),
.A2(n_2136),
.A3(n_2141),
.B1(n_2115),
.B2(n_2124),
.C1(n_2156),
.C2(n_2104),
.Y(n_2185)
);

NOR2xp67_ASAP7_75t_L g2186 ( 
.A(n_2157),
.B(n_2072),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2171),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2157),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2158),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2158),
.B(n_2132),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2158),
.Y(n_2191)
);

NOR2x1_ASAP7_75t_SL g2192 ( 
.A(n_2188),
.B(n_1967),
.Y(n_2192)
);

INVx2_ASAP7_75t_SL g2193 ( 
.A(n_2178),
.Y(n_2193)
);

OAI21xp33_ASAP7_75t_SL g2194 ( 
.A1(n_2185),
.A2(n_2141),
.B(n_2136),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2178),
.B(n_2115),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_2175),
.B(n_1969),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2189),
.B(n_2151),
.Y(n_2197)
);

OAI322xp33_ASAP7_75t_L g2198 ( 
.A1(n_2181),
.A2(n_2191),
.A3(n_2187),
.B1(n_2190),
.B2(n_2184),
.C1(n_2183),
.C2(n_2179),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_2181),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_2173),
.Y(n_2200)
);

NOR3x1_ASAP7_75t_L g2201 ( 
.A(n_2174),
.B(n_1980),
.C(n_2044),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2182),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2182),
.B(n_2148),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2177),
.Y(n_2204)
);

OR2x2_ASAP7_75t_L g2205 ( 
.A(n_2173),
.B(n_2128),
.Y(n_2205)
);

AOI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_2176),
.A2(n_2067),
.B1(n_2125),
.B2(n_2015),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2202),
.Y(n_2207)
);

NOR3x1_ASAP7_75t_L g2208 ( 
.A(n_2204),
.B(n_2180),
.C(n_2186),
.Y(n_2208)
);

AO21x1_ASAP7_75t_L g2209 ( 
.A1(n_2206),
.A2(n_2196),
.B(n_2199),
.Y(n_2209)
);

NOR2x1_ASAP7_75t_L g2210 ( 
.A(n_2198),
.B(n_1967),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_2200),
.B(n_2034),
.Y(n_2211)
);

OAI21xp5_ASAP7_75t_SL g2212 ( 
.A1(n_2193),
.A2(n_2020),
.B(n_1898),
.Y(n_2212)
);

INVx2_ASAP7_75t_SL g2213 ( 
.A(n_2197),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2194),
.B(n_2128),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_2192),
.A2(n_1983),
.B(n_1978),
.Y(n_2215)
);

AND3x4_ASAP7_75t_L g2216 ( 
.A(n_2201),
.B(n_2029),
.C(n_2005),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2197),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2195),
.B(n_2129),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2205),
.B(n_2203),
.Y(n_2219)
);

NAND5xp2_ASAP7_75t_L g2220 ( 
.A(n_2215),
.B(n_1897),
.C(n_2008),
.D(n_2067),
.E(n_2027),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_R g2221 ( 
.A(n_2207),
.B(n_1852),
.Y(n_2221)
);

OAI222xp33_ASAP7_75t_L g2222 ( 
.A1(n_2210),
.A2(n_2013),
.B1(n_2083),
.B2(n_1923),
.C1(n_1905),
.C2(n_1986),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_2210),
.B(n_2209),
.Y(n_2223)
);

AOI211xp5_ASAP7_75t_L g2224 ( 
.A1(n_2212),
.A2(n_1990),
.B(n_2006),
.C(n_1865),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2213),
.B(n_2129),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2211),
.A2(n_2013),
.B(n_2066),
.Y(n_2226)
);

INVxp67_ASAP7_75t_SL g2227 ( 
.A(n_2217),
.Y(n_2227)
);

INVx1_ASAP7_75t_SL g2228 ( 
.A(n_2219),
.Y(n_2228)
);

NAND4xp25_ASAP7_75t_SL g2229 ( 
.A(n_2214),
.B(n_1936),
.C(n_1943),
.D(n_2067),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2228),
.Y(n_2230)
);

NOR2x1_ASAP7_75t_L g2231 ( 
.A(n_2223),
.B(n_2220),
.Y(n_2231)
);

NOR2x1_ASAP7_75t_L g2232 ( 
.A(n_2222),
.B(n_2216),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2227),
.Y(n_2233)
);

HB1xp67_ASAP7_75t_L g2234 ( 
.A(n_2221),
.Y(n_2234)
);

INVxp67_ASAP7_75t_SL g2235 ( 
.A(n_2224),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2229),
.A2(n_2218),
.B1(n_2208),
.B2(n_1987),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_2226),
.B(n_2225),
.Y(n_2237)
);

NAND4xp75_ASAP7_75t_L g2238 ( 
.A(n_2231),
.B(n_1896),
.C(n_1987),
.D(n_1913),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2230),
.B(n_2111),
.Y(n_2239)
);

CKINVDCx16_ASAP7_75t_R g2240 ( 
.A(n_2234),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2232),
.B(n_2130),
.Y(n_2241)
);

AND3x4_ASAP7_75t_L g2242 ( 
.A(n_2237),
.B(n_2235),
.C(n_2236),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_2240),
.Y(n_2243)
);

NOR2xp67_ASAP7_75t_L g2244 ( 
.A(n_2239),
.B(n_2233),
.Y(n_2244)
);

NOR2x1_ASAP7_75t_L g2245 ( 
.A(n_2242),
.B(n_1905),
.Y(n_2245)
);

NAND4xp25_ASAP7_75t_L g2246 ( 
.A(n_2241),
.B(n_1923),
.C(n_1979),
.D(n_2017),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2243),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2245),
.A2(n_2238),
.B1(n_1878),
.B2(n_1889),
.Y(n_2248)
);

AO22x2_ASAP7_75t_L g2249 ( 
.A1(n_2247),
.A2(n_2248),
.B1(n_2244),
.B2(n_2246),
.Y(n_2249)
);

A2O1A1Ixp33_ASAP7_75t_SL g2250 ( 
.A1(n_2247),
.A2(n_1889),
.B(n_1878),
.C(n_1734),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2249),
.A2(n_1977),
.B1(n_1933),
.B2(n_1939),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2250),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2251),
.Y(n_2253)
);

AOI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2253),
.A2(n_2252),
.B(n_2021),
.Y(n_2254)
);

AOI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_2254),
.A2(n_1913),
.B1(n_1938),
.B2(n_1939),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2255),
.B(n_1699),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2256),
.A2(n_2031),
.B1(n_1758),
.B2(n_1727),
.Y(n_2257)
);


endmodule