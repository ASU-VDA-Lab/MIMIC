module real_aes_7210_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_617;
wire n_552;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g181 ( .A1(n_0), .A2(n_182), .B(n_183), .C(n_187), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_1), .B(n_176), .Y(n_189) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_3), .B(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_4), .A2(n_170), .B(n_476), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_5), .A2(n_150), .B(n_167), .C(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_6), .A2(n_170), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_7), .B(n_176), .Y(n_482) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_8), .A2(n_142), .B(n_264), .Y(n_263) );
AND2x6_ASAP7_75t_L g167 ( .A(n_9), .B(n_168), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_10), .A2(n_150), .B(n_167), .C(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g573 ( .A(n_11), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_12), .B(n_41), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_12), .B(n_41), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_13), .B(n_186), .Y(n_522) );
INVx1_ASAP7_75t_L g147 ( .A(n_14), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_15), .B(n_161), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_16), .A2(n_162), .B(n_531), .C(n_533), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_17), .B(n_176), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_18), .A2(n_105), .B1(n_113), .B2(n_739), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_19), .B(n_204), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_20), .A2(n_150), .B(n_196), .C(n_203), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_21), .A2(n_185), .B(n_238), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_22), .B(n_186), .Y(n_504) );
AOI222xp33_ASAP7_75t_L g451 ( .A1(n_23), .A2(n_452), .B1(n_722), .B2(n_723), .C1(n_732), .C2(n_736), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_24), .B(n_186), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_25), .Y(n_500) );
INVx1_ASAP7_75t_L g470 ( .A(n_26), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_27), .A2(n_150), .B(n_203), .C(n_267), .Y(n_266) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_28), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_29), .Y(n_518) );
INVx1_ASAP7_75t_L g494 ( .A(n_30), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_31), .A2(n_170), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_32), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g152 ( .A(n_33), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_34), .A2(n_165), .B(n_219), .C(n_220), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_35), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_36), .A2(n_185), .B(n_479), .C(n_481), .Y(n_478) );
INVxp67_ASAP7_75t_L g495 ( .A(n_37), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_38), .B(n_269), .Y(n_268) );
CKINVDCx14_ASAP7_75t_R g477 ( .A(n_39), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_40), .A2(n_150), .B(n_203), .C(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_42), .A2(n_187), .B(n_571), .C(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_43), .B(n_194), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_44), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_45), .B(n_161), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_46), .B(n_170), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_47), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_48), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_49), .A2(n_165), .B(n_219), .C(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g184 ( .A(n_50), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_51), .A2(n_67), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_51), .Y(n_130) );
INVx1_ASAP7_75t_L g248 ( .A(n_52), .Y(n_248) );
INVx1_ASAP7_75t_L g538 ( .A(n_53), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_54), .B(n_170), .Y(n_245) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_55), .A2(n_72), .B1(n_133), .B2(n_134), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_55), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_56), .Y(n_208) );
CKINVDCx14_ASAP7_75t_R g569 ( .A(n_57), .Y(n_569) );
INVx1_ASAP7_75t_L g168 ( .A(n_58), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_59), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_60), .B(n_176), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_61), .A2(n_157), .B(n_202), .C(n_259), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_62), .A2(n_71), .B1(n_729), .B2(n_730), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_62), .Y(n_729) );
INVx1_ASAP7_75t_L g146 ( .A(n_63), .Y(n_146) );
INVx1_ASAP7_75t_SL g480 ( .A(n_64), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_66), .B(n_161), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_67), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_67), .B(n_176), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_68), .B(n_162), .Y(n_235) );
INVx1_ASAP7_75t_L g503 ( .A(n_69), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_70), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_71), .Y(n_730) );
INVx1_ASAP7_75t_L g134 ( .A(n_72), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_73), .B(n_198), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_74), .A2(n_150), .B(n_155), .C(n_165), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_75), .Y(n_257) );
INVx1_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_77), .A2(n_170), .B(n_568), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_78), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_79), .A2(n_170), .B(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_80), .A2(n_194), .B(n_490), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_81), .Y(n_467) );
INVx1_ASAP7_75t_L g529 ( .A(n_82), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_83), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_83), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_84), .B(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_85), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_86), .A2(n_170), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g532 ( .A(n_87), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_88), .A2(n_724), .B1(n_725), .B2(n_731), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_88), .Y(n_724) );
INVx2_ASAP7_75t_L g144 ( .A(n_89), .Y(n_144) );
INVx1_ASAP7_75t_L g521 ( .A(n_90), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_91), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_92), .B(n_186), .Y(n_236) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_93), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g123 ( .A(n_93), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g456 ( .A(n_93), .B(n_125), .Y(n_456) );
INVx2_ASAP7_75t_L g721 ( .A(n_93), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_94), .A2(n_150), .B(n_165), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_95), .B(n_170), .Y(n_217) );
INVx1_ASAP7_75t_L g221 ( .A(n_96), .Y(n_221) );
INVxp67_ASAP7_75t_L g260 ( .A(n_97), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_98), .B(n_142), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g156 ( .A(n_100), .Y(n_156) );
INVx1_ASAP7_75t_L g231 ( .A(n_101), .Y(n_231) );
INVx2_ASAP7_75t_L g541 ( .A(n_102), .Y(n_541) );
AND2x2_ASAP7_75t_L g250 ( .A(n_103), .B(n_206), .Y(n_250) );
INVx1_ASAP7_75t_L g739 ( .A(n_105), .Y(n_739) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g125 ( .A(n_109), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_450), .Y(n_113) );
BUFx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_115), .B(n_447), .C(n_451), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_127), .B(n_447), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_123), .Y(n_449) );
NOR2x2_ASAP7_75t_L g738 ( .A(n_124), .B(n_721), .Y(n_738) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g720 ( .A(n_125), .B(n_721), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_131), .B1(n_445), .B2(n_446), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_128), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_131), .Y(n_446) );
XNOR2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_135), .Y(n_131) );
INVx1_ASAP7_75t_L g453 ( .A(n_135), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_135), .A2(n_458), .B1(n_733), .B2(n_734), .Y(n_732) );
OR3x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_353), .C(n_402), .Y(n_135) );
NAND5xp2_ASAP7_75t_L g136 ( .A(n_137), .B(n_287), .C(n_316), .D(n_324), .E(n_339), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_210), .B(n_226), .C(n_271), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_190), .Y(n_138) );
AND2x2_ASAP7_75t_L g282 ( .A(n_139), .B(n_279), .Y(n_282) );
AND2x2_ASAP7_75t_L g315 ( .A(n_139), .B(n_191), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_139), .B(n_214), .Y(n_408) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_175), .Y(n_139) );
INVx2_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
BUFx2_ASAP7_75t_L g382 ( .A(n_140), .Y(n_382) );
AO21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_148), .B(n_173), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_141), .B(n_174), .Y(n_173) );
INVx3_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_141), .B(n_225), .Y(n_224) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_141), .A2(n_230), .B(n_240), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_141), .B(n_473), .Y(n_472) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_141), .A2(n_499), .B(n_506), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_141), .B(n_524), .Y(n_523) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_142), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_142), .A2(n_265), .B(n_266), .Y(n_264) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g242 ( .A(n_143), .Y(n_242) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_144), .B(n_145), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_169), .Y(n_148) );
INVx5_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
BUFx3_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
INVx1_ASAP7_75t_L g239 ( .A(n_152), .Y(n_239) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_154), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
AND2x2_ASAP7_75t_L g171 ( .A(n_154), .B(n_172), .Y(n_171) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
INVx1_ASAP7_75t_L g269 ( .A(n_154), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_160), .C(n_163), .Y(n_155) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_158), .A2(n_161), .B1(n_494), .B2(n_495), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_158), .B(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_158), .B(n_541), .Y(n_540) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g198 ( .A(n_159), .Y(n_198) );
INVx2_ASAP7_75t_L g182 ( .A(n_161), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_161), .B(n_260), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_161), .A2(n_201), .B(n_470), .C(n_471), .Y(n_469) );
INVx5_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_162), .B(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g481 ( .A(n_164), .Y(n_481) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g178 ( .A1(n_166), .A2(n_179), .B(n_180), .C(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_166), .A2(n_180), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_166), .A2(n_180), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_166), .A2(n_180), .B(n_491), .C(n_492), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_166), .A2(n_180), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g537 ( .A1(n_166), .A2(n_180), .B(n_538), .C(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_SL g568 ( .A1(n_166), .A2(n_180), .B(n_569), .C(n_570), .Y(n_568) );
INVx4_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g170 ( .A(n_167), .B(n_171), .Y(n_170) );
BUFx3_ASAP7_75t_L g203 ( .A(n_167), .Y(n_203) );
NAND2x1p5_ASAP7_75t_L g232 ( .A(n_167), .B(n_171), .Y(n_232) );
BUFx2_ASAP7_75t_L g194 ( .A(n_170), .Y(n_194) );
INVx1_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
AND2x2_ASAP7_75t_L g190 ( .A(n_175), .B(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g280 ( .A(n_175), .Y(n_280) );
AND2x2_ASAP7_75t_L g366 ( .A(n_175), .B(n_279), .Y(n_366) );
AND2x2_ASAP7_75t_L g421 ( .A(n_175), .B(n_213), .Y(n_421) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_189), .Y(n_175) );
INVx2_ASAP7_75t_L g219 ( .A(n_180), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_185), .B(n_480), .Y(n_479) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g571 ( .A(n_186), .Y(n_571) );
INVx2_ASAP7_75t_L g505 ( .A(n_187), .Y(n_505) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_188), .Y(n_223) );
INVx1_ASAP7_75t_L g533 ( .A(n_188), .Y(n_533) );
INVx1_ASAP7_75t_L g338 ( .A(n_190), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_190), .B(n_214), .Y(n_385) );
INVx5_ASAP7_75t_L g279 ( .A(n_191), .Y(n_279) );
AND2x4_ASAP7_75t_L g300 ( .A(n_191), .B(n_280), .Y(n_300) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_191), .Y(n_322) );
AND2x2_ASAP7_75t_L g397 ( .A(n_191), .B(n_382), .Y(n_397) );
AND2x2_ASAP7_75t_L g400 ( .A(n_191), .B(n_215), .Y(n_400) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_207), .Y(n_191) );
AOI21xp5_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_195), .B(n_204), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_199), .B(n_201), .Y(n_196) );
INVx2_ASAP7_75t_L g200 ( .A(n_198), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_200), .A2(n_221), .B(n_222), .C(n_223), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_200), .A2(n_223), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_200), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
O2A1O1Ixp5_ASAP7_75t_L g520 ( .A1(n_200), .A2(n_505), .B(n_521), .C(n_522), .Y(n_520) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_202), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_205), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g209 ( .A(n_206), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_206), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_206), .A2(n_245), .B(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_206), .A2(n_232), .B(n_467), .C(n_468), .Y(n_466) );
OA21x2_ASAP7_75t_L g566 ( .A1(n_206), .A2(n_567), .B(n_574), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_209), .A2(n_517), .B(n_523), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_210), .B(n_280), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_210), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_214), .Y(n_211) );
AND2x2_ASAP7_75t_L g305 ( .A(n_212), .B(n_280), .Y(n_305) );
AND2x2_ASAP7_75t_L g323 ( .A(n_212), .B(n_215), .Y(n_323) );
INVx1_ASAP7_75t_L g343 ( .A(n_212), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_212), .B(n_279), .Y(n_388) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_212), .Y(n_430) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_213), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_214), .B(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_214), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_214), .A2(n_275), .B(n_336), .C(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g342 ( .A(n_214), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g351 ( .A(n_214), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g355 ( .A(n_214), .B(n_279), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_214), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g370 ( .A(n_214), .B(n_280), .Y(n_370) );
AND2x2_ASAP7_75t_L g420 ( .A(n_214), .B(n_421), .Y(n_420) );
INVx5_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx2_ASAP7_75t_L g284 ( .A(n_215), .Y(n_284) );
AND2x2_ASAP7_75t_L g325 ( .A(n_215), .B(n_278), .Y(n_325) );
AND2x2_ASAP7_75t_L g337 ( .A(n_215), .B(n_312), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_215), .B(n_366), .Y(n_384) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_224), .Y(n_215) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_251), .Y(n_226) );
INVx1_ASAP7_75t_L g273 ( .A(n_227), .Y(n_273) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_243), .Y(n_227) );
OR2x2_ASAP7_75t_L g275 ( .A(n_228), .B(n_243), .Y(n_275) );
NAND3xp33_ASAP7_75t_L g281 ( .A(n_228), .B(n_282), .C(n_283), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_228), .B(n_253), .Y(n_292) );
OR2x2_ASAP7_75t_L g307 ( .A(n_228), .B(n_295), .Y(n_307) );
AND2x2_ASAP7_75t_L g313 ( .A(n_228), .B(n_262), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_228), .B(n_444), .Y(n_443) );
INVx5_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_229), .B(n_253), .Y(n_310) );
AND2x2_ASAP7_75t_L g349 ( .A(n_229), .B(n_263), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_229), .B(n_262), .Y(n_377) );
OR2x2_ASAP7_75t_L g380 ( .A(n_229), .B(n_262), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_232), .A2(n_500), .B(n_501), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_232), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_237), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_237), .A2(n_268), .B(n_270), .Y(n_267) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g488 ( .A(n_242), .Y(n_488) );
INVx5_ASAP7_75t_SL g295 ( .A(n_243), .Y(n_295) );
OR2x2_ASAP7_75t_L g301 ( .A(n_243), .B(n_252), .Y(n_301) );
AND2x2_ASAP7_75t_L g317 ( .A(n_243), .B(n_318), .Y(n_317) );
AOI321xp33_ASAP7_75t_L g324 ( .A1(n_243), .A2(n_325), .A3(n_326), .B1(n_327), .B2(n_333), .C(n_335), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_243), .B(n_251), .Y(n_334) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_243), .Y(n_347) );
OR2x2_ASAP7_75t_L g394 ( .A(n_243), .B(n_292), .Y(n_394) );
AND2x2_ASAP7_75t_L g416 ( .A(n_243), .B(n_313), .Y(n_416) );
AND2x2_ASAP7_75t_L g435 ( .A(n_243), .B(n_253), .Y(n_435) );
OR2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_250), .Y(n_243) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_262), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_253), .B(n_262), .Y(n_276) );
AND2x2_ASAP7_75t_L g285 ( .A(n_253), .B(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g312 ( .A(n_253), .Y(n_312) );
AND2x2_ASAP7_75t_L g318 ( .A(n_253), .B(n_313), .Y(n_318) );
INVxp67_ASAP7_75t_L g348 ( .A(n_253), .Y(n_348) );
OR2x2_ASAP7_75t_L g390 ( .A(n_253), .B(n_295), .Y(n_390) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_261), .Y(n_253) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_254), .A2(n_475), .B(n_482), .Y(n_474) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_254), .A2(n_527), .B(n_534), .Y(n_526) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_254), .A2(n_536), .B(n_542), .Y(n_535) );
OR2x2_ASAP7_75t_L g272 ( .A(n_262), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_SL g286 ( .A(n_262), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_262), .B(n_275), .Y(n_319) );
AND2x2_ASAP7_75t_L g368 ( .A(n_262), .B(n_312), .Y(n_368) );
AND2x2_ASAP7_75t_L g406 ( .A(n_262), .B(n_295), .Y(n_406) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_263), .B(n_295), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_274), .B(n_277), .C(n_281), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_272), .A2(n_274), .B1(n_399), .B2(n_401), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_274), .A2(n_297), .B1(n_352), .B2(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_SL g426 ( .A(n_275), .Y(n_426) );
INVx1_ASAP7_75t_SL g326 ( .A(n_276), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_278), .B(n_298), .Y(n_328) );
AOI222xp33_ASAP7_75t_L g339 ( .A1(n_278), .A2(n_319), .B1(n_326), .B2(n_340), .C1(n_344), .C2(n_350), .Y(n_339) );
AND2x2_ASAP7_75t_L g429 ( .A(n_278), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_L g304 ( .A(n_279), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_279), .B(n_299), .Y(n_374) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_279), .Y(n_411) );
AND2x2_ASAP7_75t_L g414 ( .A(n_279), .B(n_323), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_279), .B(n_430), .Y(n_440) );
INVx1_ASAP7_75t_L g331 ( .A(n_280), .Y(n_331) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_280), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g422 ( .A1(n_282), .A2(n_423), .B(n_424), .C(n_427), .Y(n_422) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND3xp33_ASAP7_75t_L g345 ( .A(n_284), .B(n_346), .C(n_349), .Y(n_345) );
OR2x2_ASAP7_75t_L g373 ( .A(n_284), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_284), .B(n_300), .Y(n_401) );
OR2x2_ASAP7_75t_L g306 ( .A(n_286), .B(n_307), .Y(n_306) );
AOI211xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B(n_296), .C(n_308), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_289), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g395 ( .A(n_290), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_291), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g309 ( .A(n_294), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_295), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g363 ( .A(n_295), .B(n_313), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_295), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_295), .B(n_312), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_301), .B1(n_302), .B2(n_306), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_298), .B(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_300), .B(n_342), .Y(n_341) );
OAI221xp5_ASAP7_75t_SL g364 ( .A1(n_301), .A2(n_365), .B1(n_367), .B2(n_369), .C(n_371), .Y(n_364) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x2_ASAP7_75t_L g419 ( .A(n_304), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g432 ( .A(n_304), .B(n_421), .Y(n_432) );
INVx1_ASAP7_75t_L g352 ( .A(n_305), .Y(n_352) );
INVx1_ASAP7_75t_L g423 ( .A(n_306), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_307), .A2(n_390), .B(n_413), .Y(n_412) );
AOI21xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B(n_314), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI21xp5_ASAP7_75t_SL g316 ( .A1(n_317), .A2(n_319), .B(n_320), .Y(n_316) );
INVx1_ASAP7_75t_L g356 ( .A(n_317), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_318), .A2(n_404), .B1(n_407), .B2(n_409), .C(n_412), .Y(n_403) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_326), .A2(n_416), .B1(n_417), .B2(n_419), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g392 ( .A(n_328), .Y(n_392) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR2xp67_ASAP7_75t_SL g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AND2x2_ASAP7_75t_L g396 ( .A(n_332), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g361 ( .A(n_337), .Y(n_361) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_342), .B(n_366), .Y(n_418) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_348), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g434 ( .A(n_349), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g441 ( .A(n_349), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI211xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_356), .B(n_357), .C(n_391), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI211xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B(n_364), .C(n_383), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g444 ( .A(n_368), .Y(n_444) );
AND2x2_ASAP7_75t_L g381 ( .A(n_370), .B(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B1(n_379), .B2(n_381), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
OR2x2_ASAP7_75t_L g389 ( .A(n_377), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g442 ( .A(n_378), .Y(n_442) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI31xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .A3(n_386), .B(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI211xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_395), .C(n_398), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
NAND5xp2_ASAP7_75t_L g402 ( .A(n_403), .B(n_415), .C(n_422), .D(n_436), .E(n_439), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_414), .A2(n_440), .B1(n_441), .B2(n_443), .Y(n_439) );
INVx1_ASAP7_75t_SL g438 ( .A(n_416), .Y(n_438) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_431), .B(n_433), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_454), .B1(n_457), .B2(n_720), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g733 ( .A(n_455), .Y(n_733) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR3x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_631), .C(n_678), .Y(n_458) );
NAND3xp33_ASAP7_75t_SL g459 ( .A(n_460), .B(n_577), .C(n_602), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_515), .B1(n_543), .B2(n_546), .C(n_554), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_483), .B(n_508), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_463), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_463), .B(n_559), .Y(n_675) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
AND2x2_ASAP7_75t_L g545 ( .A(n_464), .B(n_514), .Y(n_545) );
AND2x2_ASAP7_75t_L g595 ( .A(n_464), .B(n_513), .Y(n_595) );
AND2x2_ASAP7_75t_L g616 ( .A(n_464), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g621 ( .A(n_464), .B(n_588), .Y(n_621) );
OR2x2_ASAP7_75t_L g629 ( .A(n_464), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g701 ( .A(n_464), .B(n_497), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_464), .B(n_650), .Y(n_715) );
INVx3_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g560 ( .A(n_465), .B(n_474), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_465), .B(n_497), .Y(n_561) );
AND2x4_ASAP7_75t_L g583 ( .A(n_465), .B(n_514), .Y(n_583) );
AND2x2_ASAP7_75t_L g613 ( .A(n_465), .B(n_485), .Y(n_613) );
AND2x2_ASAP7_75t_L g622 ( .A(n_465), .B(n_612), .Y(n_622) );
AND2x2_ASAP7_75t_L g638 ( .A(n_465), .B(n_498), .Y(n_638) );
OR2x2_ASAP7_75t_L g647 ( .A(n_465), .B(n_630), .Y(n_647) );
AND2x2_ASAP7_75t_L g653 ( .A(n_465), .B(n_588), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_465), .B(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g667 ( .A(n_465), .B(n_510), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_465), .B(n_556), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_465), .B(n_617), .Y(n_706) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_472), .Y(n_465) );
INVx2_ASAP7_75t_L g514 ( .A(n_474), .Y(n_514) );
AND2x2_ASAP7_75t_L g612 ( .A(n_474), .B(n_497), .Y(n_612) );
AND2x2_ASAP7_75t_L g617 ( .A(n_474), .B(n_498), .Y(n_617) );
INVx1_ASAP7_75t_L g673 ( .A(n_474), .Y(n_673) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g582 ( .A(n_484), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_497), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_485), .B(n_545), .Y(n_544) );
BUFx3_ASAP7_75t_L g559 ( .A(n_485), .Y(n_559) );
OR2x2_ASAP7_75t_L g630 ( .A(n_485), .B(n_497), .Y(n_630) );
OR2x2_ASAP7_75t_L g691 ( .A(n_485), .B(n_598), .Y(n_691) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_489), .B(n_496), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_487), .A2(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g511 ( .A(n_489), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_496), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_497), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g650 ( .A(n_497), .B(n_510), .Y(n_650) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g589 ( .A(n_498), .Y(n_589) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_509), .A2(n_695), .B1(n_699), .B2(n_702), .C(n_703), .Y(n_694) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_513), .Y(n_509) );
INVx1_ASAP7_75t_SL g557 ( .A(n_510), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_510), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g689 ( .A(n_510), .B(n_545), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_513), .B(n_559), .Y(n_681) );
AND2x2_ASAP7_75t_L g588 ( .A(n_514), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g592 ( .A(n_515), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_515), .B(n_598), .Y(n_628) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .Y(n_515) );
AND2x2_ASAP7_75t_L g553 ( .A(n_516), .B(n_526), .Y(n_553) );
INVx4_ASAP7_75t_L g565 ( .A(n_516), .Y(n_565) );
BUFx3_ASAP7_75t_L g608 ( .A(n_516), .Y(n_608) );
AND3x2_ASAP7_75t_L g623 ( .A(n_516), .B(n_624), .C(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g705 ( .A(n_525), .B(n_619), .Y(n_705) );
AND2x2_ASAP7_75t_L g713 ( .A(n_525), .B(n_598), .Y(n_713) );
INVx1_ASAP7_75t_SL g718 ( .A(n_525), .Y(n_718) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_535), .Y(n_525) );
INVx1_ASAP7_75t_SL g576 ( .A(n_526), .Y(n_576) );
AND2x2_ASAP7_75t_L g599 ( .A(n_526), .B(n_565), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_526), .B(n_549), .Y(n_601) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_526), .Y(n_641) );
OR2x2_ASAP7_75t_L g646 ( .A(n_526), .B(n_565), .Y(n_646) );
INVx2_ASAP7_75t_L g551 ( .A(n_535), .Y(n_551) );
AND2x2_ASAP7_75t_L g586 ( .A(n_535), .B(n_566), .Y(n_586) );
OR2x2_ASAP7_75t_L g606 ( .A(n_535), .B(n_566), .Y(n_606) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_535), .Y(n_626) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_544), .A2(n_585), .B(n_677), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g712 ( .A1(n_546), .A2(n_556), .A3(n_583), .B1(n_713), .B2(n_714), .C1(n_716), .C2(n_719), .Y(n_712) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_548), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_549), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g575 ( .A(n_550), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g643 ( .A(n_551), .B(n_565), .Y(n_643) );
AND2x2_ASAP7_75t_L g710 ( .A(n_551), .B(n_566), .Y(n_710) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g651 ( .A(n_553), .B(n_605), .Y(n_651) );
AOI31xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .A3(n_561), .B(n_562), .Y(n_554) );
AND2x2_ASAP7_75t_L g610 ( .A(n_556), .B(n_588), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_556), .B(n_580), .Y(n_692) );
AND2x2_ASAP7_75t_L g711 ( .A(n_556), .B(n_616), .Y(n_711) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_559), .B(n_588), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g634 ( .A(n_559), .B(n_617), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_559), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_559), .B(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_560), .B(n_617), .Y(n_649) );
INVx1_ASAP7_75t_L g693 ( .A(n_560), .Y(n_693) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_575), .Y(n_563) );
INVxp67_ASAP7_75t_L g645 ( .A(n_564), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_565), .B(n_576), .Y(n_581) );
INVx1_ASAP7_75t_L g687 ( .A(n_565), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_565), .B(n_664), .Y(n_698) );
BUFx3_ASAP7_75t_L g598 ( .A(n_566), .Y(n_598) );
AND2x2_ASAP7_75t_L g624 ( .A(n_566), .B(n_576), .Y(n_624) );
INVx2_ASAP7_75t_L g664 ( .A(n_566), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_575), .B(n_697), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_582), .B(n_584), .C(n_593), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_579), .A2(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_580), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_580), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g660 ( .A(n_581), .B(n_606), .Y(n_660) );
INVx3_ASAP7_75t_L g591 ( .A(n_583), .Y(n_591) );
OAI22xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_587), .B1(n_590), .B2(n_592), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_586), .A2(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g635 ( .A(n_586), .B(n_599), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_586), .B(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g590 ( .A(n_589), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g659 ( .A(n_589), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g603 ( .A1(n_590), .A2(n_604), .B(n_609), .Y(n_603) );
OAI22xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_596), .B1(n_600), .B2(n_601), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_595), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g619 ( .A(n_598), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_598), .B(n_641), .Y(n_640) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_614), .C(n_627), .Y(n_602) );
OAI22xp5_ASAP7_75t_SL g669 ( .A1(n_604), .A2(n_670), .B1(n_674), .B2(n_675), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g674 ( .A(n_606), .B(n_607), .Y(n_674) );
AND2x2_ASAP7_75t_L g682 ( .A(n_607), .B(n_663), .Y(n_682) );
CKINVDCx16_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_SL g690 ( .A1(n_608), .A2(n_691), .B(n_692), .C(n_693), .Y(n_690) );
OR2x2_ASAP7_75t_L g717 ( .A(n_608), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_618), .B(n_620), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_616), .A2(n_653), .B(n_654), .C(n_657), .Y(n_652) );
OAI21xp33_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_622), .B(n_623), .Y(n_620) );
AND2x2_ASAP7_75t_L g685 ( .A(n_624), .B(n_643), .Y(n_685) );
INVxp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g663 ( .A(n_626), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g668 ( .A(n_628), .Y(n_668) );
NAND3xp33_ASAP7_75t_SL g631 ( .A(n_632), .B(n_652), .C(n_665), .Y(n_631) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_636), .C(n_644), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g702 ( .A(n_639), .Y(n_702) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g662 ( .A(n_641), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_641), .B(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B(n_647), .C(n_648), .Y(n_644) );
INVx2_ASAP7_75t_SL g656 ( .A(n_646), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_647), .A2(n_658), .B1(n_660), .B2(n_661), .Y(n_657) );
OAI21xp33_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_650), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B(n_669), .C(n_676), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVxp33_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g719 ( .A(n_673), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_694), .C(n_707), .D(n_712), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_682), .B(n_683), .C(n_690), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B(n_688), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g703 ( .A1(n_684), .A2(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_691), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .Y(n_707) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g735 ( .A(n_720), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_725), .Y(n_731) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx3_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
endmodule