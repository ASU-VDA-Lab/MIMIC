module real_jpeg_16597_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_1),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_1),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_1),
.B(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_1),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_1),
.B(n_446),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_19),
.B(n_20),
.Y(n_18)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_3),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_4),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_5),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_5),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_5),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_5),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_5),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_5),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_5),
.B(n_88),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_6),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_6),
.A2(n_11),
.B1(n_119),
.B2(n_122),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_6),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_6),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_6),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_6),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_7),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_7),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_7),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_7),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_7),
.B(n_361),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_7),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_7),
.B(n_413),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_8),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_8),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_8),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_8),
.B(n_121),
.Y(n_180)
);

NAND2x1p5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_8),
.B(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_8),
.B(n_105),
.Y(n_296)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_9),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_9),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_9),
.Y(n_143)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_10),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_10),
.Y(n_225)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_11),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_11),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_11),
.B(n_101),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_11),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_11),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_11),
.B(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_11),
.B(n_476),
.Y(n_475)
);

NAND2x1_ASAP7_75t_SL g501 ( 
.A(n_11),
.B(n_502),
.Y(n_501)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_12),
.Y(n_265)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_12),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_13),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_13),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_13),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_13),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_13),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_14),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_15),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_15),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_15),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_15),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_15),
.B(n_360),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_15),
.B(n_65),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_15),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_15),
.B(n_399),
.Y(n_417)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_16),
.Y(n_111)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g448 ( 
.A(n_17),
.Y(n_448)
);

A2O1A1O1Ixp25_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_429),
.B(n_521),
.C(n_528),
.D(n_530),
.Y(n_21)
);

NAND2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_320),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_233),
.B(n_282),
.C(n_283),
.D(n_319),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_204),
.B(n_232),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g321 ( 
.A(n_25),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_156),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_26),
.B(n_156),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_102),
.C(n_127),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_27),
.B(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_67),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_45),
.Y(n_28)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_29),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_32),
.B(n_40),
.C(n_41),
.Y(n_182)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_34),
.Y(n_170)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_34),
.Y(n_458)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_35),
.A2(n_40),
.B1(n_57),
.B2(n_130),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_35),
.A2(n_40),
.B1(n_192),
.B2(n_197),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_35),
.B(n_130),
.C(n_504),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_38),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_40),
.B(n_197),
.C(n_312),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_41),
.A2(n_42),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_42),
.B(n_312),
.C(n_318),
.Y(n_459)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_45),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_56),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_47),
.A2(n_51),
.B(n_56),
.C(n_201),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_49),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_49),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_50),
.B(n_55),
.Y(n_201)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.C(n_64),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_57),
.A2(n_64),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_57),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_57),
.A2(n_100),
.B1(n_130),
.B2(n_216),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_57),
.B(n_216),
.C(n_456),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_60),
.B(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_62),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_64),
.B(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_67),
.B(n_158),
.C(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_83),
.C(n_93),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_68),
.B(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_75),
.C(n_79),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_77),
.Y(n_397)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_78),
.Y(n_343)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_78),
.Y(n_369)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_83),
.A2(n_84),
.B1(n_93),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_89),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_90),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_90),
.Y(n_179)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_93),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.C(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_94),
.A2(n_100),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_94),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_96),
.B(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_99),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_100),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_100),
.A2(n_146),
.B1(n_216),
.B2(n_267),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_100),
.B(n_267),
.C(n_304),
.Y(n_460)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_101),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_101),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_102),
.B(n_127),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_115),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_103),
.B(n_117),
.C(n_126),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_104),
.B(n_108),
.C(n_112),
.Y(n_198)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g468 ( 
.A(n_105),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_114),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_110),
.Y(n_416)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_112),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_114),
.B(n_146),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_126),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_133),
.B(n_139),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_144),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_128),
.B(n_132),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_131),
.B(n_272),
.C(n_279),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_134),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_134),
.B(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_144),
.B(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_152),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_145),
.B(n_333),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_146),
.A2(n_180),
.B1(n_181),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_146),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_146),
.B(n_181),
.C(n_262),
.Y(n_297)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_333)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_157),
.B(n_185),
.C(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_185),
.B2(n_186),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_174),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_163),
.B(n_182),
.C(n_183),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_164),
.B(n_169),
.C(n_171),
.Y(n_257)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_171),
.A2(n_439),
.B1(n_440),
.B2(n_441),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_171),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_171),
.B(n_440),
.C(n_445),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_174)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_176),
.B(n_179),
.C(n_181),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_180),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_180),
.B(n_342),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_181),
.B(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_198),
.B2(n_199),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_192),
.A2(n_197),
.B1(n_262),
.B2(n_517),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_L g529 ( 
.A(n_192),
.B(n_445),
.C(n_517),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_194),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_197),
.C(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_198),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_230),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_205),
.B(n_230),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.C(n_212),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_206),
.B(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_212),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.C(n_218),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_213),
.B(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_217),
.B(n_218),
.Y(n_331)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.C(n_226),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_219),
.B(n_226),
.Y(n_376)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_223),
.B(n_376),
.Y(n_375)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND4xp25_ASAP7_75t_SL g320 ( 
.A(n_233),
.B(n_283),
.C(n_321),
.D(n_323),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_236),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.C(n_240),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_260),
.B1(n_280),
.B2(n_281),
.Y(n_241)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_259),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_246),
.C(n_258),
.Y(n_287)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_248),
.B2(n_258),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_248),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_257),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_253),
.C(n_257),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_253),
.A2(n_254),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_253),
.B(n_472),
.C(n_475),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_254),
.B(n_299),
.C(n_451),
.Y(n_450)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_280),
.C(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_269),
.C(n_270),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_262),
.Y(n_517)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_275),
.B2(n_279),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_275),
.Y(n_279)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_286),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_287),
.B(n_289),
.C(n_301),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_301),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_300),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_290),
.B(n_293),
.C(n_294),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

AO22x1_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_295),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_296),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_297),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_309),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_302),
.B(n_310),
.C(n_311),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_305),
.B(n_457),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_305),
.B(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_312),
.B(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI21x1_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_344),
.B(n_428),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_325),
.B(n_328),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.C(n_334),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_329),
.A2(n_330),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_332),
.B(n_334),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.C(n_341),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_335),
.A2(n_336),
.B1(n_337),
.B2(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_335),
.Y(n_379)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_341),
.B(n_378),
.Y(n_377)
);

AOI21x1_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_422),
.B(n_427),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_380),
.B(n_421),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_372),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_347),
.B(n_372),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_363),
.C(n_370),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_348),
.A2(n_349),
.B1(n_388),
.B2(n_390),
.Y(n_387)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_359),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_356),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_356),
.C(n_359),
.Y(n_374)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_363),
.A2(n_370),
.B1(n_371),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_364),
.A2(n_365),
.B1(n_366),
.B2(n_367),
.Y(n_383)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_377),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_374),
.B(n_375),
.C(n_377),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_391),
.B(n_420),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_387),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_382),
.B(n_387),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.C(n_386),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_384),
.A2(n_385),
.B1(n_386),
.B2(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_386),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_388),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_392),
.A2(n_405),
.B(n_419),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_402),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_393),
.B(n_402),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_398),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_398),
.Y(n_410)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_411),
.B(n_418),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_410),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_407),
.B(n_410),
.Y(n_418)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_417),
.Y(n_411)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_423),
.B(n_424),
.Y(n_427)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NOR3xp33_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_491),
.C(n_510),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_487),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_432),
.A2(n_524),
.B(n_525),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_481),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_433),
.B(n_481),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_452),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_434),
.B(n_453),
.C(n_461),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.C(n_450),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_435),
.B(n_483),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_436),
.B(n_450),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_445),
.B2(n_449),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_445),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_445),
.A2(n_449),
.B1(n_516),
.B2(n_518),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_447),
.Y(n_502)
);

INVx8_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_451),
.A2(n_514),
.B(n_529),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_461),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_459),
.C(n_460),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_485),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_460),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_470),
.B2(n_471),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_464),
.B(n_465),
.C(n_470),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_466),
.Y(n_504)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.C(n_486),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_484),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_486),
.B(n_489),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_490),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_488),
.B(n_490),
.Y(n_524)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

A2O1A1O1Ixp25_ASAP7_75t_L g522 ( 
.A1(n_492),
.A2(n_511),
.B(n_523),
.C(n_526),
.D(n_527),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_493),
.B(n_509),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_493),
.B(n_509),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_494),
.B(n_496),
.C(n_508),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_497),
.B1(n_507),
.B2(n_508),
.Y(n_495)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_496),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_500),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_503),
.C(n_505),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_503),
.B1(n_505),
.B2(n_506),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_501),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_503),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_520),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_512),
.B(n_520),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_519),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_516),
.Y(n_518)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_529),
.Y(n_528)
);


endmodule