module real_aes_1391_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_961, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_960, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_959, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_961;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_960;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_959;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_865;
wire n_666;
wire n_551;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_550;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_936;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_867;
wire n_722;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_702;
wire n_954;
wire n_912;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_713;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_653;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_922;
wire n_633;
wire n_679;
wire n_926;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_0), .A2(n_292), .B1(n_581), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_1), .A2(n_184), .B1(n_484), .B2(n_485), .Y(n_832) );
AOI22xp33_ASAP7_75t_SL g754 ( .A1(n_2), .A2(n_103), .B1(n_517), .B2(n_545), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_3), .A2(n_89), .B1(n_484), .B2(n_485), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_4), .A2(n_213), .B1(n_577), .B2(n_578), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_5), .A2(n_20), .B1(n_517), .B2(n_947), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_6), .A2(n_80), .B1(n_546), .B2(n_670), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_7), .A2(n_145), .B1(n_480), .B2(n_481), .Y(n_633) );
AOI222xp33_ASAP7_75t_SL g446 ( .A1(n_8), .A2(n_31), .B1(n_125), .B2(n_447), .C1(n_450), .C2(n_452), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_9), .A2(n_295), .B1(n_505), .B2(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g755 ( .A1(n_10), .A2(n_109), .B1(n_426), .B2(n_551), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_11), .Y(n_645) );
AOI222xp33_ASAP7_75t_L g753 ( .A1(n_12), .A2(n_142), .B1(n_165), .B2(n_548), .C1(n_553), .C2(n_687), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_13), .A2(n_150), .B1(n_517), .B2(n_670), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_14), .A2(n_203), .B1(n_467), .B2(n_468), .Y(n_466) );
AOI222xp33_ASAP7_75t_L g878 ( .A1(n_15), .A2(n_102), .B1(n_261), .B2(n_734), .C1(n_835), .C2(n_879), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_16), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_17), .A2(n_65), .B1(n_519), .B2(n_520), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g834 ( .A1(n_18), .A2(n_314), .B1(n_339), .B2(n_426), .C1(n_513), .C2(n_835), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_19), .A2(n_28), .B1(n_423), .B2(n_426), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_21), .B(n_784), .Y(n_783) );
AOI222xp33_ASAP7_75t_L g479 ( .A1(n_22), .A2(n_83), .B1(n_154), .B2(n_480), .C1(n_481), .C2(n_482), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_23), .A2(n_215), .B1(n_538), .B2(n_539), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_24), .A2(n_134), .B1(n_539), .B2(n_569), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_25), .A2(n_216), .B1(n_481), .B2(n_520), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_26), .A2(n_224), .B1(n_805), .B2(n_853), .Y(n_852) );
INVx1_ASAP7_75t_SL g382 ( .A(n_27), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_27), .B(n_36), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_29), .A2(n_49), .B1(n_467), .B2(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_30), .A2(n_330), .B1(n_411), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_32), .A2(n_270), .B1(n_516), .B2(n_546), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_33), .A2(n_74), .B1(n_627), .B2(n_652), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_34), .A2(n_351), .B1(n_360), .B2(n_899), .C(n_913), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_35), .A2(n_50), .B1(n_444), .B2(n_496), .Y(n_891) );
AO22x2_ASAP7_75t_L g385 ( .A1(n_36), .A2(n_328), .B1(n_374), .B2(n_386), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_37), .A2(n_234), .B1(n_444), .B2(n_617), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g928 ( .A1(n_38), .A2(n_262), .B1(n_426), .B2(n_551), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_39), .A2(n_190), .B1(n_420), .B2(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_40), .A2(n_335), .B1(n_670), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_41), .A2(n_324), .B1(n_433), .B2(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g383 ( .A(n_42), .Y(n_383) );
AO22x1_ASAP7_75t_L g698 ( .A1(n_43), .A2(n_140), .B1(n_699), .B2(n_700), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_44), .A2(n_212), .B1(n_419), .B2(n_619), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_45), .A2(n_230), .B1(n_476), .B2(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_46), .B(n_482), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_47), .A2(n_96), .B1(n_519), .B2(n_520), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_48), .A2(n_113), .B1(n_742), .B2(n_820), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_51), .A2(n_52), .B1(n_665), .B2(n_666), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_53), .A2(n_915), .B1(n_916), .B2(n_930), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_53), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_54), .A2(n_329), .B1(n_538), .B2(n_539), .Y(n_826) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_55), .A2(n_191), .B1(n_225), .B2(n_593), .C1(n_666), .C2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_56), .A2(n_220), .B1(n_401), .B2(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_57), .B(n_559), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_58), .A2(n_126), .B1(n_410), .B2(n_718), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_59), .A2(n_346), .B1(n_804), .B2(n_805), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_60), .A2(n_238), .B1(n_578), .B2(n_613), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_61), .A2(n_105), .B1(n_506), .B2(n_541), .Y(n_757) );
AO22x2_ASAP7_75t_L g373 ( .A1(n_62), .A2(n_161), .B1(n_374), .B2(n_375), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_63), .A2(n_342), .B1(n_444), .B2(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_64), .A2(n_278), .B1(n_778), .B2(n_779), .Y(n_777) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_66), .A2(n_325), .B1(n_496), .B2(n_497), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_67), .A2(n_237), .B1(n_538), .B2(n_697), .Y(n_696) );
XOR2xp5_ASAP7_75t_L g706 ( .A(n_68), .B(n_707), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_69), .A2(n_558), .B(n_560), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_70), .A2(n_149), .B1(n_470), .B2(n_471), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g948 ( .A1(n_71), .A2(n_204), .B1(n_513), .B2(n_666), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_72), .B(n_553), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_73), .A2(n_112), .B1(n_619), .B2(n_771), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g949 ( .A1(n_75), .A2(n_348), .B1(n_519), .B2(n_520), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_76), .A2(n_231), .B1(n_474), .B2(n_598), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_77), .A2(n_316), .B1(n_542), .B2(n_715), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_78), .A2(n_258), .B1(n_388), .B2(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_79), .A2(n_245), .B1(n_811), .B2(n_813), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_81), .A2(n_127), .B1(n_497), .B2(n_569), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_82), .A2(n_135), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_84), .A2(n_317), .B1(n_470), .B2(n_471), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_85), .B(n_409), .Y(n_408) );
XOR2x2_ASAP7_75t_L g528 ( .A(n_86), .B(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_87), .A2(n_176), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_88), .A2(n_302), .B1(n_420), .B2(n_503), .Y(n_502) );
OA22x2_ASAP7_75t_L g841 ( .A1(n_90), .A2(n_842), .B1(n_843), .B2(n_863), .Y(n_841) );
INVx1_ASAP7_75t_L g863 ( .A(n_90), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_91), .A2(n_233), .B1(n_410), .B2(n_652), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_92), .A2(n_253), .B1(n_487), .B2(n_488), .Y(n_637) );
AOI22x1_ASAP7_75t_L g647 ( .A1(n_93), .A2(n_648), .B1(n_672), .B2(n_673), .Y(n_647) );
CKINVDCx14_ASAP7_75t_R g673 ( .A(n_93), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_94), .A2(n_151), .B1(n_470), .B2(n_471), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_95), .A2(n_180), .B1(n_426), .B2(n_513), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_97), .A2(n_321), .B1(n_415), .B2(n_418), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_98), .A2(n_286), .B1(n_781), .B2(n_782), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_99), .A2(n_331), .B1(n_411), .B2(n_468), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_100), .A2(n_185), .B1(n_541), .B2(n_542), .Y(n_540) );
AO22x2_ASAP7_75t_L g377 ( .A1(n_101), .A2(n_276), .B1(n_374), .B2(n_378), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_104), .A2(n_336), .B1(n_535), .B2(n_718), .Y(n_717) );
OA22x2_ASAP7_75t_L g866 ( .A1(n_106), .A2(n_867), .B1(n_868), .B2(n_880), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_106), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_107), .A2(n_250), .B1(n_401), .B2(n_627), .Y(n_626) );
AOI222xp33_ASAP7_75t_L g845 ( .A1(n_108), .A2(n_211), .B1(n_257), .B2(n_846), .C1(n_848), .C2(n_850), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_110), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_110), .B(n_566), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_110), .A2(n_583), .B(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_111), .A2(n_248), .B1(n_488), .B2(n_734), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_114), .A2(n_275), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_115), .A2(n_283), .B1(n_700), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_116), .A2(n_186), .B1(n_720), .B2(n_721), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_117), .A2(n_334), .B1(n_516), .B2(n_546), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_118), .A2(n_239), .B1(n_426), .B2(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_119), .A2(n_169), .B1(n_484), .B2(n_485), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_120), .A2(n_207), .B1(n_399), .B2(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_121), .A2(n_148), .B1(n_503), .B2(n_818), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_122), .A2(n_267), .B1(n_415), .B2(n_418), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_123), .A2(n_189), .B1(n_484), .B2(n_485), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_124), .A2(n_227), .B1(n_474), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_128), .A2(n_288), .B1(n_470), .B2(n_471), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_129), .A2(n_293), .B1(n_568), .B2(n_570), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_130), .A2(n_229), .B1(n_426), .B2(n_551), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_131), .A2(n_264), .B1(n_715), .B2(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_132), .A2(n_307), .B1(n_467), .B2(n_468), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_133), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_136), .A2(n_195), .B1(n_433), .B2(n_535), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_137), .A2(n_196), .B1(n_394), .B2(n_399), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_138), .A2(n_326), .B1(n_481), .B2(n_520), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g854 ( .A1(n_139), .A2(n_166), .B1(n_855), .B2(n_857), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_141), .A2(n_268), .B1(n_452), .B2(n_548), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_143), .A2(n_194), .B1(n_487), .B2(n_488), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_144), .A2(n_147), .B1(n_516), .B2(n_517), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_146), .A2(n_172), .B1(n_417), .B2(n_419), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_152), .A2(n_284), .B1(n_401), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_153), .A2(n_155), .B1(n_720), .B2(n_922), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_156), .A2(n_300), .B1(n_388), .B2(n_670), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_157), .A2(n_309), .B1(n_519), .B2(n_520), .Y(n_518) );
OA22x2_ASAP7_75t_L g727 ( .A1(n_158), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_158), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_159), .A2(n_305), .B1(n_759), .B2(n_812), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_160), .A2(n_173), .B1(n_505), .B2(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g907 ( .A(n_161), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_162), .A2(n_303), .B1(n_476), .B2(n_477), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_163), .A2(n_242), .B1(n_487), .B2(n_488), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_164), .A2(n_298), .B1(n_470), .B2(n_471), .Y(n_596) );
INVx1_ASAP7_75t_L g750 ( .A(n_167), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_168), .A2(n_349), .B1(n_570), .B2(n_617), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_170), .A2(n_219), .B1(n_811), .B2(n_813), .Y(n_810) );
OA22x2_ASAP7_75t_L g765 ( .A1(n_171), .A2(n_766), .B1(n_767), .B2(n_785), .Y(n_765) );
INVx1_ASAP7_75t_L g785 ( .A(n_171), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_174), .A2(n_263), .B1(n_532), .B2(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_175), .A2(n_205), .B1(n_418), .B2(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g407 ( .A(n_177), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_177), .A2(n_178), .B(n_432), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_177), .A2(n_438), .B1(n_457), .B2(n_961), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_178), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_179), .A2(n_244), .B1(n_467), .B2(n_563), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_181), .A2(n_256), .B1(n_440), .B2(n_444), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_182), .A2(n_235), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_183), .A2(n_251), .B1(n_759), .B2(n_812), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_187), .A2(n_197), .B1(n_538), .B2(n_721), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_188), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_192), .B(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_193), .A2(n_265), .B1(n_419), .B2(n_541), .Y(n_769) );
INVx1_ASAP7_75t_L g682 ( .A(n_198), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_199), .A2(n_285), .B1(n_415), .B2(n_418), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_200), .A2(n_236), .B1(n_444), .B2(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g356 ( .A(n_201), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_202), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_206), .A2(n_287), .B1(n_548), .B2(n_612), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_208), .A2(n_260), .B1(n_474), .B2(n_598), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_209), .A2(n_345), .B1(n_516), .B2(n_546), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_210), .A2(n_218), .B1(n_666), .B2(n_807), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_214), .A2(n_337), .B1(n_426), .B2(n_513), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_217), .A2(n_311), .B1(n_548), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_221), .A2(n_226), .B1(n_419), .B2(n_505), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_222), .A2(n_322), .B1(n_419), .B2(n_503), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_223), .A2(n_259), .B1(n_563), .B2(n_771), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_228), .A2(n_271), .B1(n_426), .B2(n_551), .Y(n_550) );
XNOR2x1_ASAP7_75t_L g608 ( .A(n_232), .B(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_240), .A2(n_289), .B1(n_476), .B2(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_241), .B(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_243), .A2(n_304), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_246), .A2(n_280), .B1(n_388), .B2(n_670), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_247), .B(n_447), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_249), .A2(n_344), .B1(n_368), .B2(n_387), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_252), .A2(n_315), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_254), .A2(n_269), .B1(n_423), .B2(n_426), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_255), .Y(n_511) );
OA22x2_ASAP7_75t_L g935 ( .A1(n_266), .A2(n_936), .B1(n_937), .B2(n_950), .Y(n_935) );
INVx1_ASAP7_75t_L g950 ( .A(n_266), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_272), .A2(n_318), .B1(n_467), .B2(n_468), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_273), .A2(n_327), .B1(n_539), .B2(n_568), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_274), .A2(n_299), .B1(n_541), .B2(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_276), .B(n_906), .Y(n_905) );
OA22x2_ASAP7_75t_L g882 ( .A1(n_277), .A2(n_883), .B1(n_894), .B2(n_895), .Y(n_882) );
INVx1_ASAP7_75t_L g894 ( .A(n_277), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_279), .A2(n_323), .B1(n_410), .B2(n_619), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_281), .B(n_553), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_282), .A2(n_320), .B1(n_563), .B2(n_742), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_290), .A2(n_310), .B1(n_548), .B2(n_549), .Y(n_547) );
INVx3_ASAP7_75t_L g374 ( .A(n_291), .Y(n_374) );
XNOR2x2_ASAP7_75t_L g586 ( .A(n_294), .B(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_296), .A2(n_313), .B1(n_467), .B2(n_468), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_297), .B(n_558), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_301), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_306), .B(n_447), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_308), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_312), .B(n_559), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_319), .A2(n_347), .B1(n_467), .B2(n_468), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_332), .A2(n_341), .B1(n_578), .B2(n_613), .Y(n_710) );
AND2x4_ASAP7_75t_L g358 ( .A(n_333), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g903 ( .A(n_333), .Y(n_903) );
AO21x1_ASAP7_75t_L g956 ( .A1(n_333), .A2(n_354), .B(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g359 ( .A(n_338), .Y(n_359) );
AND2x2_ASAP7_75t_R g932 ( .A(n_338), .B(n_903), .Y(n_932) );
INVxp67_ASAP7_75t_L g355 ( .A(n_340), .Y(n_355) );
NAND2xp33_ASAP7_75t_SL g808 ( .A(n_343), .B(n_387), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_357), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_359), .B(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g957 ( .A(n_359), .Y(n_957) );
OAI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_702), .B1(n_789), .B2(n_790), .C(n_791), .Y(n_360) );
INVx1_ASAP7_75t_L g789 ( .A(n_361), .Y(n_789) );
NAND3xp33_ASAP7_75t_L g909 ( .A(n_361), .B(n_790), .C(n_910), .Y(n_909) );
XNOR2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_604), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_524), .B1(n_525), .B2(n_603), .Y(n_362) );
INVx3_ASAP7_75t_L g603 ( .A(n_363), .Y(n_603) );
OA22x2_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_460), .B1(n_461), .B2(n_523), .Y(n_363) );
INVx2_ASAP7_75t_SL g523 ( .A(n_364), .Y(n_523) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_429), .Y(n_364) );
OAI222xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_407), .B1(n_408), .B2(n_413), .C1(n_959), .C2(n_960), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_366), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_393), .Y(n_366) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVxp33_ASAP7_75t_L g801 ( .A(n_369), .Y(n_801) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g545 ( .A(n_370), .Y(n_545) );
INVx4_ASAP7_75t_L g947 ( .A(n_370), .Y(n_947) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_371), .Y(n_516) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_371), .Y(n_670) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_379), .Y(n_371) );
AND2x4_ASAP7_75t_L g396 ( .A(n_372), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g443 ( .A(n_372), .B(n_403), .Y(n_443) );
AND2x6_ASAP7_75t_L g467 ( .A(n_372), .B(n_397), .Y(n_467) );
AND2x2_ASAP7_75t_SL g473 ( .A(n_372), .B(n_403), .Y(n_473) );
AND2x4_ASAP7_75t_L g485 ( .A(n_372), .B(n_379), .Y(n_485) );
AND2x2_ASAP7_75t_L g598 ( .A(n_372), .B(n_403), .Y(n_598) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
INVx2_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
AND2x2_ASAP7_75t_L g421 ( .A(n_373), .B(n_377), .Y(n_421) );
INVx1_ASAP7_75t_L g375 ( .A(n_374), .Y(n_375) );
INVx2_ASAP7_75t_L g378 ( .A(n_374), .Y(n_378) );
OAI22x1_ASAP7_75t_L g380 ( .A1(n_374), .A2(n_381), .B1(n_382), .B2(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_374), .Y(n_381) );
INVx1_ASAP7_75t_L g386 ( .A(n_374), .Y(n_386) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_376), .Y(n_392) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g405 ( .A(n_377), .Y(n_405) );
AND2x4_ASAP7_75t_L g412 ( .A(n_377), .B(n_406), .Y(n_412) );
AND2x4_ASAP7_75t_L g417 ( .A(n_379), .B(n_404), .Y(n_417) );
AND2x2_ASAP7_75t_L g425 ( .A(n_379), .B(n_412), .Y(n_425) );
AND2x2_ASAP7_75t_L g470 ( .A(n_379), .B(n_404), .Y(n_470) );
AND2x4_ASAP7_75t_L g488 ( .A(n_379), .B(n_412), .Y(n_488) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_384), .Y(n_379) );
AND2x2_ASAP7_75t_L g390 ( .A(n_380), .B(n_385), .Y(n_390) );
INVx2_ASAP7_75t_L g398 ( .A(n_380), .Y(n_398) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_380), .Y(n_428) );
AND2x4_ASAP7_75t_L g397 ( .A(n_384), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g403 ( .A(n_385), .B(n_398), .Y(n_403) );
BUFx2_ASAP7_75t_L g445 ( .A(n_385), .Y(n_445) );
BUFx6f_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_SL g517 ( .A(n_389), .Y(n_517) );
BUFx4f_ASAP7_75t_L g546 ( .A(n_389), .Y(n_546) );
INVx2_ASAP7_75t_L g691 ( .A(n_389), .Y(n_691) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AND2x2_ASAP7_75t_L g449 ( .A(n_390), .B(n_404), .Y(n_449) );
AND2x4_ASAP7_75t_L g454 ( .A(n_390), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g480 ( .A(n_390), .B(n_455), .Y(n_480) );
AND2x4_ASAP7_75t_L g482 ( .A(n_390), .B(n_404), .Y(n_482) );
AND2x2_ASAP7_75t_L g484 ( .A(n_390), .B(n_391), .Y(n_484) );
AND2x2_ASAP7_75t_L g520 ( .A(n_390), .B(n_455), .Y(n_520) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g532 ( .A(n_395), .Y(n_532) );
INVx2_ASAP7_75t_SL g581 ( .A(n_395), .Y(n_581) );
INVx2_ASAP7_75t_L g625 ( .A(n_395), .Y(n_625) );
INVx2_ASAP7_75t_SL g700 ( .A(n_395), .Y(n_700) );
INVx2_ASAP7_75t_L g759 ( .A(n_395), .Y(n_759) );
INVx2_ASAP7_75t_L g813 ( .A(n_395), .Y(n_813) );
INVx1_ASAP7_75t_SL g920 ( .A(n_395), .Y(n_920) );
INVx8_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g411 ( .A(n_397), .B(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g420 ( .A(n_397), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g435 ( .A(n_397), .B(n_404), .Y(n_435) );
AND2x4_ASAP7_75t_L g471 ( .A(n_397), .B(n_421), .Y(n_471) );
AND2x2_ASAP7_75t_L g476 ( .A(n_397), .B(n_412), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_397), .B(n_404), .Y(n_477) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g659 ( .A(n_402), .Y(n_659) );
BUFx2_ASAP7_75t_L g812 ( .A(n_402), .Y(n_812) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
AND2x4_ASAP7_75t_L g451 ( .A(n_403), .B(n_412), .Y(n_451) );
AND2x6_ASAP7_75t_L g468 ( .A(n_403), .B(n_404), .Y(n_468) );
AND2x2_ASAP7_75t_L g481 ( .A(n_403), .B(n_412), .Y(n_481) );
AND2x2_ASAP7_75t_L g519 ( .A(n_403), .B(n_412), .Y(n_519) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVxp67_ASAP7_75t_L g455 ( .A(n_406), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_408), .B(n_413), .C(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g507 ( .A(n_411), .Y(n_507) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_411), .Y(n_627) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_411), .Y(n_742) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_414), .B(n_422), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g534 ( .A(n_416), .Y(n_534) );
INVx3_ASAP7_75t_L g652 ( .A(n_416), .Y(n_652) );
INVx2_ASAP7_75t_L g718 ( .A(n_416), .Y(n_718) );
INVx6_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx3_ASAP7_75t_L g503 ( .A(n_417), .Y(n_503) );
BUFx3_ASAP7_75t_L g619 ( .A(n_417), .Y(n_619) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g536 ( .A(n_420), .Y(n_536) );
BUFx3_ASAP7_75t_L g656 ( .A(n_420), .Y(n_656) );
AND2x2_ASAP7_75t_L g427 ( .A(n_421), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g444 ( .A(n_421), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g474 ( .A(n_421), .B(n_445), .Y(n_474) );
AND2x2_ASAP7_75t_SL g487 ( .A(n_421), .B(n_428), .Y(n_487) );
AND2x2_ASAP7_75t_SL g734 ( .A(n_421), .B(n_428), .Y(n_734) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g781 ( .A(n_424), .Y(n_781) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx3_ASAP7_75t_L g513 ( .A(n_425), .Y(n_513) );
BUFx5_ASAP7_75t_L g551 ( .A(n_425), .Y(n_551) );
BUFx3_ASAP7_75t_L g665 ( .A(n_425), .Y(n_665) );
BUFx12f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g667 ( .A(n_427), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_436), .B(n_456), .Y(n_429) );
INVx1_ASAP7_75t_L g459 ( .A(n_432), .Y(n_459) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g505 ( .A(n_434), .Y(n_505) );
INVx2_ASAP7_75t_SL g541 ( .A(n_434), .Y(n_541) );
INVx3_ASAP7_75t_SL g563 ( .A(n_434), .Y(n_563) );
INVx4_ASAP7_75t_L g600 ( .A(n_434), .Y(n_600) );
INVx2_ASAP7_75t_L g820 ( .A(n_434), .Y(n_820) );
INVx8_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_446), .Y(n_438) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_441), .Y(n_720) );
INVx1_ASAP7_75t_L g816 ( .A(n_441), .Y(n_816) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g496 ( .A(n_442), .Y(n_496) );
INVx1_ASAP7_75t_L g617 ( .A(n_442), .Y(n_617) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_443), .Y(n_538) );
BUFx3_ASAP7_75t_L g569 ( .A(n_443), .Y(n_569) );
BUFx2_ASAP7_75t_L g497 ( .A(n_444), .Y(n_497) );
BUFx3_ASAP7_75t_L g539 ( .A(n_444), .Y(n_539) );
INVx5_ASAP7_75t_SL g571 ( .A(n_444), .Y(n_571) );
BUFx2_ASAP7_75t_L g922 ( .A(n_444), .Y(n_922) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g553 ( .A(n_448), .Y(n_553) );
INVx3_ASAP7_75t_SL g559 ( .A(n_448), .Y(n_559) );
INVx4_ASAP7_75t_SL g593 ( .A(n_448), .Y(n_593) );
BUFx2_ASAP7_75t_L g662 ( .A(n_448), .Y(n_662) );
INVx4_ASAP7_75t_SL g784 ( .A(n_448), .Y(n_784) );
INVx6_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx4f_ASAP7_75t_SL g577 ( .A(n_450), .Y(n_577) );
BUFx2_ASAP7_75t_L g804 ( .A(n_450), .Y(n_804) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx3_ASAP7_75t_L g548 ( .A(n_451), .Y(n_548) );
BUFx2_ASAP7_75t_L g613 ( .A(n_451), .Y(n_613) );
BUFx2_ASAP7_75t_L g778 ( .A(n_451), .Y(n_778) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g549 ( .A(n_453), .Y(n_549) );
INVx2_ASAP7_75t_SL g578 ( .A(n_453), .Y(n_578) );
INVx2_ASAP7_75t_L g612 ( .A(n_453), .Y(n_612) );
INVx2_ASAP7_75t_SL g687 ( .A(n_453), .Y(n_687) );
INVx2_ASAP7_75t_L g779 ( .A(n_453), .Y(n_779) );
INVx2_ASAP7_75t_L g805 ( .A(n_453), .Y(n_805) );
INVx6_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_490), .B(n_521), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g522 ( .A(n_463), .Y(n_522) );
XNOR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_489), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_478), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_466), .B(n_469), .C(n_472), .D(n_475), .Y(n_465) );
INVx1_ASAP7_75t_L g500 ( .A(n_468), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .C(n_486), .Y(n_478) );
INVx2_ASAP7_75t_SL g510 ( .A(n_482), .Y(n_510) );
BUFx2_ASAP7_75t_L g835 ( .A(n_482), .Y(n_835) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_488), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_490), .B(n_522), .Y(n_521) );
XNOR2x1_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_493), .B(n_508), .Y(n_492) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_494), .B(n_501), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g542 ( .A(n_507), .Y(n_542) );
INVx1_ASAP7_75t_L g771 ( .A(n_507), .Y(n_771) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .Y(n_508) );
OAI21xp5_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_509) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_513), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .Y(n_514) );
BUFx6f_ASAP7_75t_SL g853 ( .A(n_516), .Y(n_853) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_585), .B1(n_601), .B2(n_602), .Y(n_525) );
INVx1_ASAP7_75t_L g602 ( .A(n_526), .Y(n_602) );
XOR2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_554), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2xp67_ASAP7_75t_L g529 ( .A(n_530), .B(n_543), .Y(n_529) );
NAND4xp25_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .C(n_537), .D(n_540), .Y(n_530) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g924 ( .A(n_536), .Y(n_924) );
NAND4xp25_ASAP7_75t_L g543 ( .A(n_544), .B(n_547), .C(n_550), .D(n_552), .Y(n_543) );
INVx1_ASAP7_75t_L g851 ( .A(n_548), .Y(n_851) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_572), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B(n_564), .C(n_565), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_556), .B(n_557), .C(n_580), .Y(n_579) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g847 ( .A(n_559), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_564), .B(n_567), .C(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g697 ( .A(n_571), .Y(n_697) );
INVx3_ASAP7_75t_L g721 ( .A(n_571), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_579), .B(n_582), .Y(n_572) );
INVx1_ASAP7_75t_L g584 ( .A(n_574), .Y(n_584) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g583 ( .A(n_580), .Y(n_583) );
BUFx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g601 ( .A(n_586), .Y(n_601) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_594), .Y(n_587) );
NAND4xp25_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .C(n_591), .D(n_592), .Y(n_588) );
NAND4xp25_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .C(n_597), .D(n_599), .Y(n_594) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_600), .Y(n_713) );
AO22x2_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_678), .B2(n_701), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AO22x2_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_628), .B1(n_676), .B2(n_677), .Y(n_606) );
INVx1_ASAP7_75t_L g676 ( .A(n_607), .Y(n_676) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND4xp75_ASAP7_75t_L g609 ( .A(n_610), .B(n_615), .C(n_620), .D(n_623), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx2_ASAP7_75t_L g677 ( .A(n_628), .Y(n_677) );
OA22x2_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_646), .B1(n_647), .B2(n_674), .Y(n_628) );
AO22x2_ASAP7_75t_L g679 ( .A1(n_629), .A2(n_674), .B1(n_680), .B2(n_681), .Y(n_679) );
XOR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_645), .Y(n_629) );
XOR2x2_ASAP7_75t_L g675 ( .A(n_630), .B(n_645), .Y(n_675) );
NAND2x1_ASAP7_75t_SL g630 ( .A(n_631), .B(n_638), .Y(n_630) );
NOR2x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NOR2x1_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g672 ( .A(n_648), .Y(n_672) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_660), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_654), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g699 ( .A(n_659), .Y(n_699) );
INVx2_ASAP7_75t_SL g715 ( .A(n_659), .Y(n_715) );
INVx2_ASAP7_75t_L g773 ( .A(n_659), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_668), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_663), .B(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g724 ( .A(n_665), .Y(n_724) );
BUFx6f_ASAP7_75t_SL g807 ( .A(n_665), .Y(n_807) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g782 ( .A(n_667), .Y(n_782) );
INVx2_ASAP7_75t_L g856 ( .A(n_667), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g701 ( .A(n_678), .Y(n_701) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
XNOR2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_684), .B(n_692), .Y(n_683) );
AND4x1_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .C(n_688), .D(n_689), .Y(n_684) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g849 ( .A(n_691), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_698), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .C(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g790 ( .A(n_702), .Y(n_790) );
OAI22x1_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_745), .B1(n_746), .B2(n_788), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_705), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_725), .B1(n_726), .B2(n_744), .Y(n_705) );
INVx1_ASAP7_75t_L g744 ( .A(n_706), .Y(n_744) );
NAND4xp75_ASAP7_75t_SL g707 ( .A(n_708), .B(n_711), .C(n_716), .D(n_722), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AOI22x1_ASAP7_75t_SL g748 ( .A1(n_726), .A2(n_727), .B1(n_749), .B2(n_762), .Y(n_748) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NOR2x1_ASAP7_75t_L g730 ( .A(n_731), .B(n_737), .Y(n_730) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .C(n_735), .D(n_736), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_741), .C(n_743), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_742), .Y(n_818) );
INVx4_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OA22x2_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B1(n_763), .B2(n_786), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g762 ( .A(n_749), .Y(n_762) );
XNOR2x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
OR2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_756), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .C(n_755), .Y(n_752) );
NAND4xp25_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .C(n_760), .D(n_761), .Y(n_756) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
BUFx2_ASAP7_75t_L g787 ( .A(n_765), .Y(n_787) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NOR2x1_ASAP7_75t_L g767 ( .A(n_768), .B(n_775), .Y(n_767) );
NAND4xp25_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .C(n_772), .D(n_774), .Y(n_768) );
NAND4xp25_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .C(n_780), .D(n_783), .Y(n_775) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_789), .B(n_912), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_790), .B(n_900), .Y(n_912) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OAI211xp5_ASAP7_75t_L g899 ( .A1(n_792), .A2(n_900), .B(n_909), .C(n_911), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_838), .B1(n_839), .B2(n_898), .Y(n_792) );
INVx1_ASAP7_75t_L g898 ( .A(n_793), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_821), .B1(n_822), .B2(n_837), .Y(n_793) );
INVx2_ASAP7_75t_L g837 ( .A(n_794), .Y(n_837) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
XNOR2x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
OR2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_809), .Y(n_797) );
NAND4xp25_ASAP7_75t_L g798 ( .A(n_799), .B(n_803), .C(n_806), .D(n_808), .Y(n_798) );
OA21x2_ASAP7_75t_SL g799 ( .A1(n_800), .A2(n_801), .B(n_802), .Y(n_799) );
NAND4xp25_ASAP7_75t_L g809 ( .A(n_810), .B(n_814), .C(n_817), .D(n_819), .Y(n_809) );
BUFx3_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
XOR2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_836), .Y(n_823) );
NAND4xp75_ASAP7_75t_L g824 ( .A(n_825), .B(n_828), .C(n_831), .D(n_834), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AO22x2_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_864), .B1(n_896), .B2(n_897), .Y(n_840) );
INVx1_ASAP7_75t_L g896 ( .A(n_841), .Y(n_896) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
OR2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_858), .Y(n_843) );
NAND3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_852), .C(n_854), .Y(n_844) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
BUFx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NAND4xp25_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .C(n_861), .D(n_862), .Y(n_858) );
INVx1_ASAP7_75t_L g897 ( .A(n_864), .Y(n_897) );
AO22x1_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_866), .B1(n_881), .B2(n_882), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g880 ( .A(n_868), .Y(n_880) );
NAND4xp75_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .C(n_875), .D(n_878), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
AND2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
AND2x2_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g895 ( .A(n_883), .Y(n_895) );
NOR2x1_ASAP7_75t_L g883 ( .A(n_884), .B(n_889), .Y(n_883) );
NAND4xp25_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .C(n_887), .D(n_888), .Y(n_884) );
NAND4xp25_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .C(n_892), .D(n_893), .Y(n_889) );
INVx1_ASAP7_75t_L g910 ( .A(n_900), .Y(n_910) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_902), .B(n_905), .Y(n_953) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
OAI222xp33_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_931), .B1(n_933), .B2(n_950), .C1(n_951), .C2(n_954), .Y(n_913) );
INVxp67_ASAP7_75t_SL g915 ( .A(n_916), .Y(n_915) );
OR2x2_ASAP7_75t_L g916 ( .A(n_917), .B(n_925), .Y(n_916) );
NAND4xp25_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .C(n_921), .D(n_923), .Y(n_917) );
NAND4xp25_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .C(n_928), .D(n_929), .Y(n_925) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
NOR2xp67_ASAP7_75t_L g937 ( .A(n_938), .B(n_944), .Y(n_937) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_942), .C(n_943), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .Y(n_939) );
NAND4xp25_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .C(n_948), .D(n_949), .Y(n_944) );
INVx1_ASAP7_75t_SL g951 ( .A(n_952), .Y(n_951) );
CKINVDCx6p67_ASAP7_75t_R g952 ( .A(n_953), .Y(n_952) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_955), .Y(n_954) );
CKINVDCx20_ASAP7_75t_R g955 ( .A(n_956), .Y(n_955) );
endmodule