module fake_aes_860_n_630 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_630);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_630;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_12), .Y(n_76) );
BUFx2_ASAP7_75t_L g77 ( .A(n_39), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_38), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_53), .Y(n_79) );
BUFx2_ASAP7_75t_L g80 ( .A(n_3), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_3), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_42), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_33), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_73), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_24), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_74), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_35), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_40), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_20), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_1), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_8), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_27), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_57), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_64), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_68), .Y(n_95) );
NOR2xp33_ASAP7_75t_L g96 ( .A(n_48), .B(n_51), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_17), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_45), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_70), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_46), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_0), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_30), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_55), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_50), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_36), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_60), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_75), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_26), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_59), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_9), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_69), .Y(n_112) );
NOR2xp67_ASAP7_75t_L g113 ( .A(n_11), .B(n_65), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_41), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_56), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_43), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_62), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_17), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_54), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_10), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_16), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_72), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g123 ( .A(n_77), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_121), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_87), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_85), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_87), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_121), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_80), .B(n_1), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_77), .B(n_2), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_121), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_85), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_80), .Y(n_134) );
NAND2xp33_ASAP7_75t_R g135 ( .A(n_89), .B(n_47), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_78), .A2(n_67), .B(n_66), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_120), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_117), .B(n_2), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_107), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_104), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_119), .B(n_4), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_118), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_105), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_118), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_88), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_120), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_76), .B(n_4), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_107), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_76), .B(n_5), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_78), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_107), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_114), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_81), .B(n_5), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_79), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_114), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_79), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_82), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_122), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_109), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_81), .B(n_6), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_122), .Y(n_163) );
NAND3xp33_ASAP7_75t_L g164 ( .A(n_134), .B(n_90), .C(n_97), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_148), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_153), .B(n_99), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_125), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_134), .B(n_99), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_130), .B(n_129), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_126), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_144), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
AO22x2_ASAP7_75t_L g178 ( .A1(n_130), .A2(n_95), .B1(n_94), .B2(n_93), .Y(n_178) );
NAND3xp33_ASAP7_75t_L g179 ( .A(n_160), .B(n_90), .C(n_97), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
NOR2x1p5_ASAP7_75t_L g181 ( .A(n_140), .B(n_91), .Y(n_181) );
AND2x6_ASAP7_75t_L g182 ( .A(n_130), .B(n_82), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_125), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_133), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_148), .A2(n_101), .B1(n_111), .B2(n_118), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_146), .B(n_102), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_132), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_129), .B(n_101), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_163), .A2(n_111), .B1(n_118), .B2(n_108), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_129), .A2(n_118), .B1(n_116), .B2(n_115), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_127), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_127), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_150), .B(n_118), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_150), .Y(n_199) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_150), .B(n_116), .Y(n_200) );
INVxp67_ASAP7_75t_SL g201 ( .A(n_141), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_136), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_133), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_141), .A2(n_84), .B1(n_98), .B2(n_112), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_154), .B(n_115), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_154), .B(n_100), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_154), .Y(n_207) );
NAND2x1p5_ASAP7_75t_L g208 ( .A(n_151), .B(n_98), .Y(n_208) );
AND2x6_ASAP7_75t_L g209 ( .A(n_151), .B(n_100), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_155), .B(n_83), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_139), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_139), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_127), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_139), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_139), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_139), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_155), .B(n_102), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_152), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_152), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_201), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_198), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_172), .B(n_158), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_198), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_207), .B(n_183), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_182), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_182), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_172), .B(n_123), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_172), .B(n_138), .Y(n_229) );
INVx5_ASAP7_75t_L g230 ( .A(n_182), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_182), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_207), .B(n_159), .Y(n_232) );
INVx4_ASAP7_75t_L g233 ( .A(n_182), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_209), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_176), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_189), .Y(n_237) );
OR2x6_ASAP7_75t_L g238 ( .A(n_200), .B(n_162), .Y(n_238) );
AO22x1_ASAP7_75t_L g239 ( .A1(n_173), .A2(n_143), .B1(n_162), .B2(n_158), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_208), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_206), .B(n_159), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_199), .B(n_113), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_208), .B(n_109), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_206), .B(n_124), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_209), .Y(n_245) );
BUFx12f_ASAP7_75t_L g246 ( .A(n_173), .Y(n_246) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_196), .A2(n_136), .B(n_128), .Y(n_247) );
NOR3xp33_ASAP7_75t_SL g248 ( .A(n_190), .B(n_135), .C(n_93), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_189), .B(n_128), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_182), .Y(n_250) );
NAND3xp33_ASAP7_75t_SL g251 ( .A(n_190), .B(n_94), .C(n_92), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_181), .Y(n_252) );
NOR2xp33_ASAP7_75t_R g253 ( .A(n_182), .B(n_131), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_174), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_191), .B(n_137), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_200), .B(n_131), .Y(n_256) );
AND2x6_ASAP7_75t_L g257 ( .A(n_165), .B(n_83), .Y(n_257) );
NAND3xp33_ASAP7_75t_SL g258 ( .A(n_204), .B(n_86), .C(n_92), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_209), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_191), .B(n_137), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_191), .B(n_113), .Y(n_261) );
BUFx10_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
OR2x6_ASAP7_75t_L g263 ( .A(n_200), .B(n_86), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_205), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_208), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_205), .Y(n_266) );
NOR3xp33_ASAP7_75t_L g267 ( .A(n_179), .B(n_95), .C(n_112), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_171), .B(n_145), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_205), .A2(n_156), .B1(n_152), .B2(n_145), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_170), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_189), .B(n_161), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_170), .Y(n_272) );
AND2x6_ASAP7_75t_SL g273 ( .A(n_218), .B(n_147), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_205), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_184), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_205), .B(n_147), .Y(n_276) );
NAND2xp33_ASAP7_75t_SL g277 ( .A(n_166), .B(n_103), .Y(n_277) );
AOI21xp33_ASAP7_75t_L g278 ( .A1(n_178), .A2(n_103), .B(n_106), .Y(n_278) );
NOR3xp33_ASAP7_75t_SL g279 ( .A(n_164), .B(n_106), .C(n_110), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_174), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_205), .B(n_156), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_243), .A2(n_167), .B(n_202), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_221), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_234), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_225), .B(n_188), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_228), .A2(n_178), .B1(n_209), .B2(n_168), .Y(n_286) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_247), .A2(n_196), .B(n_202), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_241), .B(n_178), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_270), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_278), .A2(n_220), .B(n_219), .C(n_194), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_266), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_268), .B(n_178), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_243), .A2(n_202), .B(n_196), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_271), .A2(n_169), .B(n_210), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_226), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_229), .B(n_192), .Y(n_296) );
BUFx5_ASAP7_75t_L g297 ( .A(n_262), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_255), .B(n_218), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_238), .B(n_197), .Y(n_299) );
INVx3_ASAP7_75t_SL g300 ( .A(n_263), .Y(n_300) );
O2A1O1Ixp5_ASAP7_75t_L g301 ( .A1(n_277), .A2(n_193), .B(n_197), .C(n_184), .Y(n_301) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_226), .B(n_220), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_266), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_234), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_272), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_263), .A2(n_209), .B1(n_186), .B2(n_168), .Y(n_306) );
AND2x2_ASAP7_75t_SL g307 ( .A(n_266), .B(n_136), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_260), .B(n_209), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_228), .A2(n_209), .B1(n_197), .B2(n_187), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_263), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_222), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_223), .B(n_219), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_236), .B(n_194), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_235), .B(n_187), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_232), .B(n_214), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_238), .B(n_214), .Y(n_316) );
AND2x4_ASAP7_75t_SL g317 ( .A(n_238), .B(n_156), .Y(n_317) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_226), .B(n_136), .Y(n_318) );
CKINVDCx6p67_ASAP7_75t_R g319 ( .A(n_238), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_240), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_224), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_244), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_265), .B(n_110), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_275), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_274), .Y(n_325) );
AND3x1_ASAP7_75t_SL g326 ( .A(n_246), .B(n_6), .C(n_7), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_262), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_233), .B(n_7), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_233), .B(n_8), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_283), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_300), .B(n_239), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_311), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_300), .A2(n_246), .B1(n_229), .B2(n_228), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_322), .B(n_233), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_316), .B(n_250), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_285), .B(n_273), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_305), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_319), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_289), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_298), .A2(n_258), .B1(n_242), .B2(n_261), .C(n_252), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_316), .A2(n_229), .B1(n_264), .B2(n_252), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_296), .B(n_261), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_310), .B(n_250), .Y(n_343) );
AOI21x1_ASAP7_75t_L g344 ( .A1(n_287), .A2(n_242), .B(n_213), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_292), .A2(n_286), .B1(n_319), .B2(n_288), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_316), .B(n_250), .Y(n_346) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_310), .A2(n_264), .B1(n_274), .B2(n_227), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_293), .A2(n_281), .B(n_276), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_SL g349 ( .A1(n_290), .A2(n_271), .B(n_256), .C(n_251), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_313), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_321), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_328), .A2(n_277), .B1(n_257), .B2(n_267), .Y(n_352) );
NOR2x1_ASAP7_75t_SL g353 ( .A(n_320), .B(n_230), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_306), .A2(n_269), .B1(n_231), .B2(n_227), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_302), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_289), .Y(n_357) );
OAI211xp5_ASAP7_75t_SL g358 ( .A1(n_313), .A2(n_314), .B(n_248), .C(n_279), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_294), .A2(n_301), .B(n_305), .C(n_324), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
AOI222xp33_ASAP7_75t_L g361 ( .A1(n_355), .A2(n_261), .B1(n_242), .B2(n_323), .C1(n_315), .C2(n_329), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_339), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_337), .B(n_320), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_342), .A2(n_323), .B1(n_312), .B2(n_299), .C(n_269), .Y(n_364) );
OAI22xp5_ASAP7_75t_SL g365 ( .A1(n_338), .A2(n_329), .B1(n_328), .B2(n_326), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_356), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_350), .A2(n_299), .B1(n_328), .B2(n_329), .C(n_249), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_336), .A2(n_358), .B1(n_340), .B2(n_345), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
INVxp67_ASAP7_75t_L g370 ( .A(n_331), .Y(n_370) );
OA21x2_ASAP7_75t_L g371 ( .A1(n_344), .A2(n_290), .B(n_282), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_356), .B(n_331), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_334), .A2(n_257), .B1(n_317), .B2(n_308), .Y(n_373) );
INVx4_ASAP7_75t_L g374 ( .A(n_356), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_332), .A2(n_249), .B1(n_317), .B2(n_309), .C(n_237), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_352), .A2(n_302), .B1(n_291), .B2(n_303), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_357), .A2(n_302), .B1(n_291), .B2(n_303), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g378 ( .A1(n_338), .A2(n_257), .B1(n_253), .B2(n_307), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_357), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_334), .A2(n_257), .B1(n_325), .B2(n_295), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_337), .A2(n_257), .B1(n_325), .B2(n_295), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_344), .A2(n_295), .B(n_212), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_359), .A2(n_307), .B(n_318), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_360), .B(n_237), .Y(n_384) );
OAI211xp5_ASAP7_75t_L g385 ( .A1(n_333), .A2(n_253), .B(n_139), .C(n_149), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_356), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_356), .A2(n_318), .B1(n_231), .B2(n_262), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_367), .A2(n_341), .B1(n_360), .B2(n_351), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_368), .A2(n_330), .B1(n_349), .B2(n_354), .C(n_161), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_379), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_369), .B(n_346), .Y(n_391) );
AOI21x1_ASAP7_75t_L g392 ( .A1(n_382), .A2(n_383), .B(n_371), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_386), .Y(n_393) );
OAI22xp5_ASAP7_75t_SL g394 ( .A1(n_365), .A2(n_343), .B1(n_96), .B2(n_353), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_365), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_367), .A2(n_378), .B1(n_363), .B2(n_377), .Y(n_396) );
OAI211xp5_ASAP7_75t_SL g397 ( .A1(n_370), .A2(n_142), .B(n_185), .C(n_195), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_369), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_362), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_382), .A2(n_348), .B(n_215), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_383), .A2(n_377), .B(n_376), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_362), .B(n_346), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_361), .A2(n_335), .B1(n_343), .B2(n_347), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_362), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_363), .Y(n_406) );
OAI21xp33_ASAP7_75t_L g407 ( .A1(n_361), .A2(n_149), .B(n_161), .Y(n_407) );
OAI211xp5_ASAP7_75t_SL g408 ( .A1(n_372), .A2(n_142), .B(n_185), .C(n_195), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_374), .Y(n_409) );
AOI222xp33_ASAP7_75t_L g410 ( .A1(n_364), .A2(n_343), .B1(n_335), .B2(n_353), .C1(n_161), .C2(n_149), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_386), .B(n_348), .Y(n_411) );
NAND3xp33_ASAP7_75t_SL g412 ( .A(n_364), .B(n_203), .C(n_211), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_374), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_363), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_363), .B(n_149), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_366), .Y(n_416) );
INVx3_ASAP7_75t_SL g417 ( .A(n_374), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_384), .B(n_149), .Y(n_418) );
AOI33xp33_ASAP7_75t_L g419 ( .A1(n_384), .A2(n_203), .A3(n_211), .B1(n_212), .B2(n_213), .B3(n_215), .Y(n_419) );
INVx5_ASAP7_75t_L g420 ( .A(n_366), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_366), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_399), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_399), .B(n_366), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_398), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_403), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_405), .B(n_366), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_409), .B(n_366), .Y(n_427) );
AND2x4_ASAP7_75t_SL g428 ( .A(n_403), .B(n_380), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_411), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_405), .B(n_371), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_411), .Y(n_431) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_414), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_409), .B(n_371), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_401), .B(n_371), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_421), .B(n_149), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_390), .B(n_376), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_421), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_402), .B(n_149), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_413), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_413), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_416), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_416), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_407), .A2(n_385), .B(n_375), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_393), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_402), .B(n_161), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_417), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_420), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_388), .A2(n_161), .B1(n_142), .B2(n_373), .C(n_381), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_392), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_392), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_417), .B(n_161), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_418), .B(n_9), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_407), .B(n_410), .C(n_419), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_396), .A2(n_387), .B1(n_230), .B2(n_304), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_400), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_418), .B(n_10), .Y(n_456) );
OR2x6_ASAP7_75t_L g457 ( .A(n_406), .B(n_304), .Y(n_457) );
AO21x1_ASAP7_75t_L g458 ( .A1(n_404), .A2(n_11), .B(n_12), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_417), .B(n_13), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_394), .A2(n_284), .B1(n_237), .B2(n_175), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_415), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_415), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_391), .B(n_13), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_391), .B(n_14), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_395), .A2(n_142), .B1(n_175), .B2(n_177), .C(n_180), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_400), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_420), .B(n_14), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_395), .A2(n_175), .B1(n_177), .B2(n_180), .C(n_216), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_463), .B(n_404), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g470 ( .A(n_453), .B(n_389), .C(n_397), .D(n_408), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_424), .B(n_15), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_444), .B(n_15), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_463), .B(n_420), .Y(n_473) );
NAND2xp33_ASAP7_75t_SL g474 ( .A(n_446), .B(n_420), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_458), .A2(n_412), .B1(n_420), .B2(n_175), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_444), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_464), .B(n_16), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_453), .B(n_18), .C(n_19), .D(n_20), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g479 ( .A(n_459), .B(n_18), .C(n_19), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_425), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_425), .Y(n_481) );
NOR2xp67_ASAP7_75t_SL g482 ( .A(n_459), .B(n_420), .Y(n_482) );
OR2x6_ASAP7_75t_L g483 ( .A(n_447), .B(n_284), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_452), .B(n_21), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_437), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_452), .B(n_21), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_429), .B(n_22), .Y(n_487) );
AND2x2_ASAP7_75t_SL g488 ( .A(n_436), .B(n_259), .Y(n_488) );
NOR3xp33_ASAP7_75t_SL g489 ( .A(n_454), .B(n_22), .C(n_23), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_452), .B(n_23), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_464), .B(n_25), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_456), .B(n_28), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_467), .Y(n_493) );
INVx6_ASAP7_75t_L g494 ( .A(n_467), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_456), .B(n_29), .Y(n_495) );
NOR4xp25_ASAP7_75t_SL g496 ( .A(n_468), .B(n_31), .C(n_32), .D(n_34), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_456), .B(n_37), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_458), .A2(n_216), .B1(n_175), .B2(n_180), .Y(n_498) );
OAI211xp5_ASAP7_75t_SL g499 ( .A1(n_460), .A2(n_448), .B(n_443), .C(n_436), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_439), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_439), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_429), .B(n_216), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_440), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_440), .B(n_216), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_447), .B(n_234), .Y(n_505) );
NAND2x1p5_ASAP7_75t_L g506 ( .A(n_467), .B(n_230), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_437), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_422), .B(n_44), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_461), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_462), .B(n_217), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_462), .B(n_49), .Y(n_511) );
CKINVDCx8_ASAP7_75t_R g512 ( .A(n_427), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_437), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_431), .B(n_52), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_438), .B(n_58), .Y(n_515) );
OR2x6_ASAP7_75t_L g516 ( .A(n_457), .B(n_327), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_431), .B(n_61), .Y(n_517) );
AOI21xp33_ASAP7_75t_SL g518 ( .A1(n_479), .A2(n_451), .B(n_457), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_476), .Y(n_519) );
AO22x2_ASAP7_75t_L g520 ( .A1(n_480), .A2(n_431), .B1(n_434), .B2(n_432), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_509), .B(n_434), .Y(n_521) );
NAND4xp25_ASAP7_75t_L g522 ( .A(n_478), .B(n_434), .C(n_465), .D(n_433), .Y(n_522) );
NAND4xp25_ASAP7_75t_L g523 ( .A(n_498), .B(n_465), .C(n_433), .D(n_438), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_493), .B(n_427), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_477), .B(n_428), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_500), .B(n_430), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_501), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_503), .Y(n_528) );
AND3x1_ASAP7_75t_L g529 ( .A(n_489), .B(n_423), .C(n_449), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_489), .A2(n_451), .B(n_445), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_484), .A2(n_445), .B1(n_450), .B2(n_435), .C(n_430), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_473), .B(n_423), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_472), .A2(n_435), .B(n_450), .C(n_449), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_485), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_474), .B(n_428), .Y(n_535) );
XNOR2x2_ASAP7_75t_L g536 ( .A(n_486), .B(n_423), .Y(n_536) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_498), .A2(n_475), .B(n_491), .Y(n_537) );
AOI32xp33_ASAP7_75t_L g538 ( .A1(n_490), .A2(n_435), .A3(n_426), .B1(n_449), .B2(n_466), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_469), .B(n_426), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_494), .B(n_442), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_487), .B(n_441), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_492), .Y(n_542) );
OAI322xp33_ASAP7_75t_L g543 ( .A1(n_471), .A2(n_441), .A3(n_442), .B1(n_455), .B2(n_216), .C1(n_217), .C2(n_180), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_494), .B(n_442), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_494), .B(n_441), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_487), .B(n_457), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_491), .B(n_457), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_483), .Y(n_548) );
OAI32xp33_ASAP7_75t_L g549 ( .A1(n_480), .A2(n_455), .A3(n_457), .B1(n_63), .B2(n_327), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_485), .B(n_455), .Y(n_550) );
AO32x1_ASAP7_75t_L g551 ( .A1(n_495), .A2(n_280), .A3(n_254), .B1(n_217), .B2(n_177), .Y(n_551) );
AOI21xp33_ASAP7_75t_L g552 ( .A1(n_482), .A2(n_177), .B(n_180), .Y(n_552) );
AO22x2_ASAP7_75t_L g553 ( .A1(n_481), .A2(n_297), .B1(n_280), .B2(n_254), .Y(n_553) );
NOR2xp33_ASAP7_75t_R g554 ( .A(n_512), .B(n_230), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_499), .B(n_177), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_497), .Y(n_556) );
AOI322xp5_ASAP7_75t_L g557 ( .A1(n_488), .A2(n_217), .A3(n_234), .B1(n_245), .B2(n_259), .C1(n_297), .C2(n_481), .Y(n_557) );
AOI222xp33_ASAP7_75t_L g558 ( .A1(n_499), .A2(n_217), .B1(n_245), .B2(n_259), .C1(n_297), .C2(n_488), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_519), .B(n_507), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_527), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_528), .Y(n_561) );
AOI21xp33_ASAP7_75t_L g562 ( .A1(n_533), .A2(n_508), .B(n_516), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_539), .B(n_513), .Y(n_563) );
NOR4xp25_ASAP7_75t_SL g564 ( .A(n_518), .B(n_505), .C(n_516), .D(n_506), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_542), .B(n_470), .Y(n_565) );
XNOR2x2_ASAP7_75t_L g566 ( .A(n_536), .B(n_517), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_550), .Y(n_567) );
OAI322xp33_ASAP7_75t_L g568 ( .A1(n_521), .A2(n_514), .A3(n_502), .B1(n_510), .B2(n_504), .C1(n_506), .C2(n_511), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_531), .B(n_516), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_556), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_532), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_529), .B(n_505), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_520), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_529), .B(n_496), .C(n_515), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_526), .B(n_483), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_534), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_541), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_538), .B(n_483), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_537), .B(n_245), .Y(n_579) );
NOR3xp33_ASAP7_75t_SL g580 ( .A(n_535), .B(n_297), .C(n_245), .Y(n_580) );
NOR2x1_ASAP7_75t_L g581 ( .A(n_543), .B(n_259), .Y(n_581) );
AOI21xp33_ASAP7_75t_L g582 ( .A1(n_548), .A2(n_297), .B(n_555), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_522), .B(n_297), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_522), .A2(n_525), .B1(n_547), .B2(n_546), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_554), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_520), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_540), .B(n_544), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_545), .B(n_524), .Y(n_588) );
NAND2x1_ASAP7_75t_SL g589 ( .A(n_586), .B(n_553), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_573), .A2(n_543), .B1(n_549), .B2(n_530), .C(n_553), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_565), .A2(n_557), .B(n_558), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_588), .B(n_557), .Y(n_592) );
XNOR2x1_ASAP7_75t_L g593 ( .A(n_566), .B(n_523), .Y(n_593) );
OA22x2_ASAP7_75t_L g594 ( .A1(n_578), .A2(n_523), .B1(n_551), .B2(n_552), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_560), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_561), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_573), .B(n_551), .C(n_565), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_SL g598 ( .A1(n_564), .A2(n_551), .B(n_579), .C(n_584), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_572), .A2(n_578), .B(n_579), .Y(n_599) );
AOI221x1_ASAP7_75t_L g600 ( .A1(n_574), .A2(n_582), .B1(n_569), .B2(n_583), .C(n_562), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_588), .B(n_587), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_572), .A2(n_585), .B1(n_570), .B2(n_566), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_577), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_581), .B(n_580), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_559), .B(n_576), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_592), .B(n_571), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_602), .A2(n_568), .B(n_575), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_605), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_592), .B(n_567), .Y(n_609) );
OAI311xp33_ASAP7_75t_L g610 ( .A1(n_591), .A2(n_563), .A3(n_587), .B1(n_590), .C1(n_597), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_593), .B(n_603), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_593), .A2(n_594), .B1(n_604), .B2(n_605), .Y(n_612) );
AOI21xp33_ASAP7_75t_SL g613 ( .A1(n_594), .A2(n_604), .B(n_601), .Y(n_613) );
OAI22xp5_ASAP7_75t_SL g614 ( .A1(n_598), .A2(n_600), .B1(n_595), .B2(n_596), .Y(n_614) );
AO22x2_ASAP7_75t_L g615 ( .A1(n_589), .A2(n_593), .B1(n_586), .B2(n_600), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_598), .A2(n_593), .B1(n_602), .B2(n_592), .Y(n_616) );
AOI211x1_ASAP7_75t_L g617 ( .A1(n_602), .A2(n_599), .B(n_591), .C(n_597), .Y(n_617) );
INVxp33_ASAP7_75t_SL g618 ( .A(n_599), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_616), .B(n_617), .Y(n_619) );
NAND3xp33_ASAP7_75t_SL g620 ( .A(n_612), .B(n_613), .C(n_607), .Y(n_620) );
AOI22xp33_ASAP7_75t_R g621 ( .A1(n_608), .A2(n_610), .B1(n_615), .B2(n_618), .Y(n_621) );
CKINVDCx12_ASAP7_75t_R g622 ( .A(n_614), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_619), .Y(n_623) );
XOR2xp5_ASAP7_75t_L g624 ( .A(n_620), .B(n_615), .Y(n_624) );
XNOR2xp5_ASAP7_75t_L g625 ( .A(n_621), .B(n_611), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_624), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_623), .Y(n_627) );
INVx2_ASAP7_75t_SL g628 ( .A(n_627), .Y(n_628) );
AOI22xp5_ASAP7_75t_SL g629 ( .A1(n_628), .A2(n_626), .B1(n_625), .B2(n_622), .Y(n_629) );
AO21x2_ASAP7_75t_L g630 ( .A1(n_629), .A2(n_606), .B(n_609), .Y(n_630) );
endmodule