module fake_jpeg_3843_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_14),
.A2(n_2),
.B(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_35),
.Y(n_62)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_17),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_1),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_45),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_18),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_57),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_52),
.B1(n_36),
.B2(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_16),
.B1(n_20),
.B2(n_28),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_55),
.B1(n_61),
.B2(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_58),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_16),
.B1(n_20),
.B2(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_16),
.B1(n_20),
.B2(n_28),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_16),
.B(n_17),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_46),
.B1(n_55),
.B2(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_67),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_78),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_20),
.B1(n_36),
.B2(n_38),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_35),
.B1(n_52),
.B2(n_31),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_20),
.B1(n_35),
.B2(n_36),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_56),
.B1(n_57),
.B2(n_48),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_85),
.B(n_48),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_87),
.A2(n_91),
.B1(n_39),
.B2(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_88),
.B(n_67),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_44),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_90),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_53),
.B(n_41),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_49),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_93),
.B(n_97),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_103),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_76),
.C(n_68),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_72),
.C(n_76),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_99),
.A2(n_101),
.B1(n_70),
.B2(n_88),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_48),
.B1(n_42),
.B2(n_62),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_60),
.B1(n_35),
.B2(n_31),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_62),
.C(n_33),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_114),
.Y(n_154)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_71),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_99),
.A3(n_97),
.B1(n_74),
.B2(n_90),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_107),
.A2(n_76),
.B1(n_80),
.B2(n_74),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_128),
.B1(n_129),
.B2(n_86),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_74),
.B(n_83),
.C(n_42),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_106),
.B(n_34),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_27),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_54),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_54),
.B1(n_71),
.B2(n_66),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_60),
.B1(n_39),
.B2(n_33),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_34),
.B(n_15),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_23),
.B(n_21),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_100),
.B1(n_23),
.B2(n_92),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_106),
.C(n_94),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_139),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_106),
.C(n_94),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_150),
.B(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_129),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_157),
.B(n_23),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_84),
.B1(n_100),
.B2(n_104),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_149),
.B1(n_111),
.B2(n_122),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_47),
.B1(n_66),
.B2(n_27),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_152),
.B1(n_120),
.B2(n_148),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_100),
.B1(n_86),
.B2(n_92),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_21),
.B(n_24),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_81),
.C(n_73),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_158),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_113),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_169),
.B1(n_177),
.B2(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_123),
.B1(n_130),
.B2(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_109),
.B1(n_116),
.B2(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_151),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_178),
.B(n_179),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_119),
.B1(n_130),
.B2(n_131),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_25),
.B(n_24),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_73),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_24),
.B1(n_25),
.B2(n_95),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_81),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_148),
.B1(n_153),
.B2(n_134),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_137),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_187),
.A2(n_184),
.B(n_172),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_154),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_192),
.C(n_200),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_158),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_181),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_139),
.C(n_141),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_136),
.C(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_135),
.C(n_95),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_27),
.Y(n_208)
);

BUFx12_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_213),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_165),
.B1(n_171),
.B2(n_179),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_220),
.B1(n_224),
.B2(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_221),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_217),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_168),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_222),
.B(n_228),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_176),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_227),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_167),
.B1(n_183),
.B2(n_162),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_163),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_174),
.B(n_182),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_225),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_172),
.B1(n_166),
.B2(n_161),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_192),
.C(n_200),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_230),
.C(n_237),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_190),
.C(n_199),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_186),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_240),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_244),
.B(n_224),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_204),
.C(n_206),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_208),
.C(n_189),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_237),
.C(n_230),
.Y(n_260)
);

XOR2x2_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_193),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_245),
.B(n_1),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_194),
.B1(n_25),
.B2(n_47),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_13),
.B1(n_12),
.B2(n_27),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_135),
.B(n_13),
.C(n_12),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_27),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_214),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_238),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_210),
.B1(n_223),
.B2(n_215),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_253),
.B1(n_248),
.B2(n_260),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_233),
.Y(n_263)
);

OAI321xp33_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_210),
.A3(n_26),
.B1(n_19),
.B2(n_13),
.C(n_12),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_47),
.B1(n_82),
.B2(n_26),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_1),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_2),
.B(n_3),
.Y(n_265)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_259),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_29),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_245),
.B(n_2),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_229),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_26),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_261),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_265),
.B(n_252),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_273),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_255),
.B(n_26),
.C(n_19),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_273),
.C(n_268),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_253),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_240),
.Y(n_273)
);

OA21x2_ASAP7_75t_SL g276 ( 
.A1(n_263),
.A2(n_255),
.B(n_252),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_280),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_278),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_281),
.A2(n_283),
.B1(n_284),
.B2(n_3),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_26),
.B(n_19),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_265),
.A3(n_271),
.B1(n_272),
.B2(n_267),
.C1(n_19),
.C2(n_8),
.Y(n_285)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_19),
.B(n_27),
.Y(n_284)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_3),
.A3(n_6),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_29),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_27),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_289)
);

AOI332xp33_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_290),
.A3(n_291),
.B1(n_11),
.B2(n_29),
.B3(n_146),
.C1(n_54),
.C2(n_37),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_27),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_9),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_9),
.C2(n_10),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_275),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_11),
.C(n_29),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_296),
.Y(n_297)
);

AOI32xp33_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_29),
.A3(n_287),
.B1(n_295),
.B2(n_298),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_299),
.Y(n_300)
);


endmodule