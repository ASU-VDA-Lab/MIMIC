module fake_aes_8953_n_670 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_670);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_670;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_63), .Y(n_74) );
INVxp67_ASAP7_75t_SL g75 ( .A(n_49), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_37), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_33), .Y(n_77) );
INVx1_ASAP7_75t_SL g78 ( .A(n_21), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_11), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_61), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_56), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_24), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_8), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_67), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_25), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_71), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_50), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_23), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_7), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_46), .Y(n_90) );
INVx1_ASAP7_75t_SL g91 ( .A(n_25), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_21), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_31), .Y(n_93) );
CKINVDCx14_ASAP7_75t_R g94 ( .A(n_41), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_20), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_19), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_23), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_28), .Y(n_98) );
HB1xp67_ASAP7_75t_L g99 ( .A(n_36), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_51), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_64), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_73), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_38), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_35), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_65), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_40), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_45), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_18), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_30), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_43), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_39), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_57), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_18), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_7), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_15), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_59), .Y(n_119) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_11), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_54), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_70), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_86), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_99), .B(n_0), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_92), .B(n_0), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_115), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_115), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_79), .B(n_1), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_115), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_74), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_74), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_79), .B(n_85), .Y(n_132) );
NOR2xp33_ASAP7_75t_R g133 ( .A(n_94), .B(n_29), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_115), .Y(n_134) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_76), .A2(n_27), .B(n_68), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_77), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_77), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_80), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_80), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_115), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_105), .Y(n_141) );
NAND2xp33_ASAP7_75t_SL g142 ( .A(n_98), .B(n_1), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_76), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_107), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_87), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_85), .B(n_2), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_121), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_100), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_87), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_90), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_92), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_90), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_82), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_101), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_101), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_83), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_96), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_88), .B(n_89), .Y(n_158) );
INVx1_ASAP7_75t_SL g159 ( .A(n_118), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_103), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_88), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_120), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_89), .B(n_2), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_103), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_104), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_151), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_132), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_161), .B(n_95), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_155), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_155), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_128), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_159), .B(n_93), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_130), .B(n_84), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_132), .B(n_122), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
INVxp67_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_130), .B(n_97), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_161), .Y(n_184) );
AND2x6_ASAP7_75t_L g185 ( .A(n_128), .B(n_122), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_146), .A2(n_113), .B1(n_95), .B2(n_116), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_148), .B(n_119), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_123), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_162), .B(n_119), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_146), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_146), .A2(n_113), .B1(n_109), .B2(n_102), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_131), .B(n_106), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_153), .B(n_106), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_146), .B(n_104), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_158), .B(n_108), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_160), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_160), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_131), .B(n_108), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g202 ( .A1(n_141), .A2(n_117), .B1(n_78), .B2(n_91), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_136), .B(n_112), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_160), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_127), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_160), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_157), .B(n_112), .Y(n_208) );
AND2x2_ASAP7_75t_SL g209 ( .A(n_124), .B(n_111), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_158), .B(n_111), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_160), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_136), .B(n_110), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_125), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_137), .B(n_110), .Y(n_214) );
INVx4_ASAP7_75t_SL g215 ( .A(n_160), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_158), .B(n_114), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_125), .A2(n_81), .B1(n_75), .B2(n_5), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_137), .B(n_3), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_127), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_164), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_149), .B(n_3), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_164), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_149), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_127), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_164), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_150), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_170), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g232 ( .A(n_179), .B(n_144), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_184), .B(n_165), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_230), .Y(n_234) );
OR2x6_ASAP7_75t_L g235 ( .A(n_184), .B(n_124), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_230), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_227), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_196), .B(n_165), .Y(n_238) );
BUFx12f_ASAP7_75t_L g239 ( .A(n_206), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_206), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_216), .A2(n_142), .B1(n_154), .B2(n_152), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_227), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_172), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_225), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_225), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_196), .B(n_145), .Y(n_247) );
NAND2x1p5_ASAP7_75t_L g248 ( .A(n_195), .B(n_149), .Y(n_248) );
INVxp67_ASAP7_75t_SL g249 ( .A(n_170), .Y(n_249) );
NAND2xp33_ASAP7_75t_SL g250 ( .A(n_176), .B(n_147), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_195), .B(n_133), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_196), .B(n_145), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_174), .B(n_154), .Y(n_253) );
NOR2xp33_ASAP7_75t_SL g254 ( .A(n_195), .B(n_163), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_186), .A2(n_163), .B1(n_152), .B2(n_138), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_168), .B(n_139), .Y(n_256) );
INVx3_ASAP7_75t_SL g257 ( .A(n_216), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_196), .B(n_139), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_210), .B(n_138), .Y(n_259) );
NAND2xp33_ASAP7_75t_R g260 ( .A(n_188), .B(n_135), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_210), .B(n_135), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_213), .Y(n_262) );
NAND3xp33_ASAP7_75t_SL g263 ( .A(n_166), .B(n_150), .C(n_143), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_202), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_170), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_225), .Y(n_266) );
INVx4_ASAP7_75t_L g267 ( .A(n_225), .Y(n_267) );
NOR3xp33_ASAP7_75t_SL g268 ( .A(n_202), .B(n_4), .C(n_5), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_172), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_207), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_216), .A2(n_149), .B1(n_150), .B2(n_143), .Y(n_271) );
NOR2xp33_ASAP7_75t_R g272 ( .A(n_171), .B(n_47), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_181), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_216), .Y(n_274) );
NAND3xp33_ASAP7_75t_L g275 ( .A(n_191), .B(n_143), .C(n_140), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_181), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_216), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_210), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_210), .B(n_135), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_168), .B(n_4), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_216), .B(n_6), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_209), .B(n_140), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_181), .Y(n_283) );
INVxp67_ASAP7_75t_L g284 ( .A(n_175), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_176), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_207), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_176), .B(n_129), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_209), .B(n_140), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_185), .Y(n_289) );
NOR2xp33_ASAP7_75t_R g290 ( .A(n_171), .B(n_42), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_209), .B(n_134), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_167), .B(n_134), .Y(n_292) );
NOR2xp33_ASAP7_75t_R g293 ( .A(n_171), .B(n_44), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_167), .B(n_134), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_219), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_183), .B(n_126), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_185), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_208), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_171), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_280), .B(n_176), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_258), .B(n_185), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_239), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_257), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_254), .A2(n_185), .B1(n_189), .B2(n_187), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_279), .A2(n_173), .B(n_190), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_261), .A2(n_173), .B(n_190), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_258), .B(n_185), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_253), .A2(n_173), .B(n_190), .C(n_214), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_257), .Y(n_309) );
NOR3xp33_ASAP7_75t_L g310 ( .A(n_240), .B(n_217), .C(n_193), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_239), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_248), .A2(n_185), .B1(n_173), .B2(n_190), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_258), .B(n_185), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_235), .Y(n_314) );
OR2x6_ASAP7_75t_L g315 ( .A(n_248), .B(n_221), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_281), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_297), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_280), .B(n_177), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_250), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_281), .A2(n_221), .B1(n_212), .B2(n_201), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_278), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_278), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_273), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_231), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_234), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_280), .B(n_192), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_256), .B(n_203), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_257), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_245), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_262), .B(n_6), .Y(n_330) );
BUFx2_ASAP7_75t_SL g331 ( .A(n_281), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_256), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_235), .B(n_215), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_248), .B(n_8), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_284), .B(n_9), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_298), .B(n_235), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_235), .B(n_215), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_242), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_273), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_250), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_233), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_261), .A2(n_229), .B(n_169), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_289), .B(n_215), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_299), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_234), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_299), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_296), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g349 ( .A(n_289), .B(n_198), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_297), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_236), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_332), .A2(n_264), .B1(n_232), .B2(n_255), .C1(n_247), .C2(n_238), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_341), .B(n_241), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g355 ( .A1(n_314), .A2(n_264), .B1(n_242), .B2(n_277), .Y(n_355) );
INVx5_ASAP7_75t_SL g356 ( .A(n_333), .Y(n_356) );
NAND2xp33_ASAP7_75t_SL g357 ( .A(n_314), .B(n_297), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_348), .Y(n_358) );
INVx6_ASAP7_75t_L g359 ( .A(n_300), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_300), .B(n_277), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_331), .A2(n_267), .B1(n_246), .B2(n_266), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_326), .A2(n_263), .B1(n_246), .B2(n_266), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_302), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g364 ( .A(n_303), .B(n_267), .Y(n_364) );
NAND2xp33_ASAP7_75t_R g365 ( .A(n_333), .B(n_261), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_326), .A2(n_271), .B1(n_252), .B2(n_259), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_319), .A2(n_267), .B1(n_274), .B2(n_245), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_300), .B(n_265), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_326), .A2(n_245), .B1(n_241), .B2(n_236), .Y(n_370) );
NAND2xp33_ASAP7_75t_L g371 ( .A(n_317), .B(n_245), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_310), .A2(n_268), .B1(n_275), .B2(n_251), .C(n_282), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_315), .A2(n_245), .B1(n_249), .B2(n_265), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_333), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_325), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_327), .B(n_231), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
OR2x6_ASAP7_75t_L g378 ( .A(n_315), .B(n_283), .Y(n_378) );
NOR3xp33_ASAP7_75t_SL g379 ( .A(n_302), .B(n_311), .C(n_340), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_315), .A2(n_283), .B1(n_288), .B2(n_291), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_334), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_336), .A2(n_275), .B1(n_231), .B2(n_276), .C(n_292), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_318), .B(n_276), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_311), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_352), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_352), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_358), .B(n_315), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_353), .A2(n_319), .B1(n_318), .B2(n_316), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_375), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_365), .A2(n_340), .B1(n_260), .B2(n_304), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_381), .A2(n_334), .B1(n_318), .B2(n_351), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_354), .B(n_345), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_360), .B(n_345), .Y(n_393) );
AOI21xp33_ASAP7_75t_L g394 ( .A1(n_370), .A2(n_335), .B(n_305), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_378), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_369), .A2(n_308), .B1(n_320), .B2(n_323), .C(n_339), .Y(n_396) );
OAI222xp33_ASAP7_75t_L g397 ( .A1(n_378), .A2(n_337), .B1(n_312), .B2(n_344), .C1(n_338), .C2(n_346), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_372), .A2(n_346), .B1(n_337), .B2(n_321), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_365), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_377), .A2(n_306), .B1(n_322), .B2(n_307), .C(n_301), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_360), .B(n_337), .Y(n_401) );
OAI221xp5_ASAP7_75t_SL g402 ( .A1(n_366), .A2(n_313), .B1(n_328), .B2(n_309), .C(n_324), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_378), .A2(n_366), .B1(n_380), .B2(n_362), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_376), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_374), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_383), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_359), .Y(n_407) );
OA21x2_ASAP7_75t_L g408 ( .A1(n_382), .A2(n_342), .B(n_126), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_362), .A2(n_324), .B1(n_329), .B2(n_276), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_368), .B(n_324), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_363), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_355), .B(n_347), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_356), .B(n_309), .Y(n_413) );
AOI221xp5_ASAP7_75t_SL g414 ( .A1(n_403), .A2(n_361), .B1(n_373), .B2(n_371), .C(n_126), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_403), .A2(n_359), .B1(n_368), .B2(n_374), .Y(n_415) );
AO21x2_ASAP7_75t_L g416 ( .A1(n_394), .A2(n_272), .B(n_290), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_385), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_391), .A2(n_359), .B1(n_384), .B2(n_356), .C1(n_357), .C2(n_328), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_386), .Y(n_419) );
AO21x1_ASAP7_75t_SL g420 ( .A1(n_399), .A2(n_356), .B(n_364), .Y(n_420) );
NOR2xp33_ASAP7_75t_R g421 ( .A(n_411), .B(n_303), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_388), .A2(n_391), .B1(n_398), .B2(n_396), .C(n_400), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_388), .A2(n_367), .B1(n_379), .B2(n_364), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_385), .Y(n_425) );
OAI33xp33_ASAP7_75t_L g426 ( .A1(n_390), .A2(n_197), .A3(n_169), .B1(n_178), .B2(n_229), .B3(n_180), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_390), .A2(n_350), .B(n_317), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_402), .A2(n_303), .B1(n_379), .B2(n_350), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_389), .B(n_9), .Y(n_430) );
OAI31xp33_ASAP7_75t_SL g431 ( .A1(n_387), .A2(n_343), .A3(n_12), .B(n_13), .Y(n_431) );
AOI33xp33_ASAP7_75t_L g432 ( .A1(n_398), .A2(n_194), .A3(n_178), .B1(n_180), .B2(n_223), .B3(n_182), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_399), .A2(n_293), .B1(n_347), .B2(n_317), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_389), .B(n_10), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_386), .A2(n_350), .B(n_317), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_404), .Y(n_436) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_394), .A2(n_194), .B(n_197), .Y(n_437) );
INVx6_ASAP7_75t_L g438 ( .A(n_393), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_405), .Y(n_439) );
AOI211xp5_ASAP7_75t_L g440 ( .A1(n_402), .A2(n_294), .B(n_287), .C(n_127), .Y(n_440) );
OAI33xp33_ASAP7_75t_L g441 ( .A1(n_406), .A2(n_182), .A3(n_199), .B1(n_200), .B2(n_204), .B3(n_211), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_393), .B(n_10), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_396), .A2(n_237), .B1(n_243), .B2(n_349), .C(n_285), .Y(n_443) );
AOI33xp33_ASAP7_75t_L g444 ( .A1(n_387), .A2(n_199), .A3(n_200), .B1(n_204), .B2(n_211), .B3(n_218), .Y(n_444) );
OA21x2_ASAP7_75t_L g445 ( .A1(n_400), .A2(n_218), .B(n_223), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_387), .A2(n_317), .B1(n_350), .B2(n_237), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_404), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_409), .B(n_127), .C(n_129), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_404), .A2(n_350), .B1(n_349), .B2(n_285), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_436), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_436), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_447), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g453 ( .A1(n_431), .A2(n_395), .B1(n_407), .B2(n_410), .C(n_406), .Y(n_453) );
OAI21xp33_ASAP7_75t_L g454 ( .A1(n_431), .A2(n_409), .B(n_404), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_417), .B(n_395), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_417), .B(n_395), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_419), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_419), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_447), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_430), .B(n_397), .C(n_395), .Y(n_460) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_422), .A2(n_412), .B1(n_397), .B2(n_407), .C1(n_392), .C2(n_405), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_447), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_425), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_425), .B(n_405), .Y(n_464) );
AND2x6_ASAP7_75t_SL g465 ( .A(n_442), .B(n_430), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_434), .B(n_410), .C(n_413), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_423), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_423), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_427), .B(n_392), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_439), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_437), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_440), .B(n_127), .C(n_129), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_440), .B(n_127), .C(n_129), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_434), .B(n_408), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_437), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_415), .B(n_408), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_445), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_429), .B(n_408), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_437), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_445), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_445), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_424), .A2(n_408), .B(n_412), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_437), .Y(n_483) );
OA332x1_ASAP7_75t_L g484 ( .A1(n_429), .A2(n_12), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_16), .C1(n_17), .C2(n_19), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_438), .B(n_408), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_445), .B(n_408), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_424), .B(n_412), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_438), .Y(n_489) );
AND2x4_ASAP7_75t_SL g490 ( .A(n_420), .B(n_401), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_449), .B(n_448), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_438), .B(n_401), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_438), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_418), .B(n_401), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_418), .B(n_413), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_416), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_432), .Y(n_497) );
NAND3xp33_ASAP7_75t_SL g498 ( .A(n_472), .B(n_421), .C(n_444), .Y(n_498) );
OAI211xp5_ASAP7_75t_SL g499 ( .A1(n_470), .A2(n_413), .B(n_446), .C(n_433), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_461), .B(n_414), .C(n_129), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_452), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_469), .B(n_463), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_488), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_450), .B(n_428), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_487), .B(n_420), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_466), .B(n_20), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
NAND2xp33_ASAP7_75t_SL g508 ( .A(n_488), .B(n_416), .Y(n_508) );
CKINVDCx6p67_ASAP7_75t_R g509 ( .A(n_490), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_465), .B(n_426), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_452), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_465), .B(n_22), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_451), .B(n_448), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_462), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_464), .B(n_22), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_455), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_489), .B(n_435), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_455), .B(n_24), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_456), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_494), .B(n_441), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_490), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_456), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g524 ( .A(n_497), .B(n_343), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_495), .B(n_416), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_459), .Y(n_526) );
AND2x2_ASAP7_75t_SL g527 ( .A(n_490), .B(n_416), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_459), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_457), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_467), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_460), .B(n_129), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_457), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_474), .B(n_443), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_474), .B(n_219), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_485), .B(n_26), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_487), .B(n_32), .Y(n_536) );
NAND2xp33_ASAP7_75t_SL g537 ( .A(n_491), .B(n_343), .Y(n_537) );
OAI33xp33_ASAP7_75t_L g538 ( .A1(n_497), .A2(n_226), .A3(n_224), .B1(n_220), .B2(n_53), .B3(n_55), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_493), .B(n_224), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_458), .B(n_34), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_472), .B(n_220), .C(n_226), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_468), .B(n_48), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_493), .B(n_52), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_468), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_489), .B(n_58), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_489), .B(n_60), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_492), .B(n_62), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_504), .B(n_485), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_507), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_502), .B(n_476), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_516), .B(n_482), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_509), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_509), .Y(n_553) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_512), .B(n_453), .C(n_473), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_510), .A2(n_454), .B1(n_473), .B2(n_484), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_520), .B(n_454), .Y(n_556) );
OAI21xp33_ASAP7_75t_L g557 ( .A1(n_510), .A2(n_478), .B(n_496), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_511), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_526), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_522), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_523), .B(n_477), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_528), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_522), .Y(n_563) );
CKINVDCx16_ASAP7_75t_R g564 ( .A(n_503), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_504), .B(n_478), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_498), .A2(n_491), .B(n_496), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_530), .Y(n_567) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_521), .A2(n_496), .B1(n_481), .B2(n_477), .C(n_480), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_521), .A2(n_476), .B1(n_481), .B2(n_480), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_529), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_529), .Y(n_571) );
OA21x2_ASAP7_75t_L g572 ( .A1(n_525), .A2(n_479), .B(n_483), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g573 ( .A1(n_506), .A2(n_496), .B1(n_481), .B2(n_483), .C(n_479), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_505), .Y(n_574) );
OAI21xp33_ASAP7_75t_L g575 ( .A1(n_531), .A2(n_486), .B(n_481), .Y(n_575) );
NOR2x2_ASAP7_75t_L g576 ( .A(n_501), .B(n_475), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_511), .B(n_486), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_500), .A2(n_475), .B1(n_471), .B2(n_349), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_504), .B(n_471), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_501), .B(n_66), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_515), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_532), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_532), .Y(n_584) );
OAI32xp33_ASAP7_75t_L g585 ( .A1(n_537), .A2(n_69), .A3(n_198), .B1(n_243), .B2(n_269), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_527), .B(n_205), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_536), .Y(n_587) );
NOR2x1p5_ASAP7_75t_L g588 ( .A(n_533), .B(n_205), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_499), .A2(n_198), .B1(n_205), .B2(n_222), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_544), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_541), .A2(n_269), .B(n_295), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_513), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_527), .A2(n_205), .B1(n_222), .B2(n_228), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_569), .B(n_514), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_L g595 ( .A1(n_554), .A2(n_524), .B(n_543), .C(n_534), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_549), .Y(n_596) );
OAI31xp33_ASAP7_75t_L g597 ( .A1(n_553), .A2(n_508), .A3(n_535), .B(n_513), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_574), .B(n_517), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_564), .A2(n_535), .B1(n_513), .B2(n_517), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_550), .B(n_544), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_559), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_548), .B(n_518), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_562), .Y(n_603) );
XNOR2x2_ASAP7_75t_L g604 ( .A(n_586), .B(n_540), .Y(n_604) );
NOR2xp33_ASAP7_75t_R g605 ( .A(n_552), .B(n_547), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_558), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_570), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_579), .B(n_568), .Y(n_608) );
INVxp33_ASAP7_75t_SL g609 ( .A(n_560), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_582), .B(n_556), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_576), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_551), .B(n_518), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_567), .B(n_518), .Y(n_613) );
NOR4xp25_ASAP7_75t_SL g614 ( .A(n_586), .B(n_538), .C(n_542), .D(n_545), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_558), .B(n_539), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_561), .Y(n_616) );
XOR2x2_ASAP7_75t_L g617 ( .A(n_555), .B(n_546), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_570), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_577), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_566), .A2(n_538), .B(n_270), .C(n_286), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_571), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_548), .B(n_205), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_563), .Y(n_623) );
AOI32xp33_ASAP7_75t_L g624 ( .A1(n_552), .A2(n_270), .A3(n_295), .B1(n_286), .B2(n_244), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_557), .A2(n_222), .B(n_228), .Y(n_625) );
AOI21xp5_ASAP7_75t_SL g626 ( .A1(n_599), .A2(n_588), .B(n_578), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_609), .B(n_587), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_608), .B(n_573), .C(n_589), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_614), .A2(n_585), .B(n_575), .Y(n_629) );
INVxp67_ASAP7_75t_L g630 ( .A(n_606), .Y(n_630) );
AOI321xp33_ASAP7_75t_L g631 ( .A1(n_599), .A2(n_565), .A3(n_580), .B1(n_592), .B2(n_593), .C(n_581), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_623), .Y(n_632) );
XOR2xp5_ASAP7_75t_L g633 ( .A(n_623), .B(n_580), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_616), .B(n_619), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_597), .A2(n_592), .B1(n_572), .B2(n_584), .C(n_583), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_610), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_594), .A2(n_580), .B1(n_590), .B2(n_584), .C(n_583), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_SL g638 ( .A1(n_609), .A2(n_576), .B(n_571), .C(n_590), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_612), .B(n_572), .Y(n_639) );
XOR2x2_ASAP7_75t_L g640 ( .A(n_617), .B(n_591), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_596), .B(n_222), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_626), .A2(n_605), .B(n_624), .C(n_625), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_640), .A2(n_617), .B1(n_628), .B2(n_636), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_634), .Y(n_644) );
AOI221xp5_ASAP7_75t_SL g645 ( .A1(n_635), .A2(n_602), .B1(n_595), .B2(n_603), .C(n_601), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g646 ( .A(n_633), .B(n_604), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_627), .A2(n_613), .B1(n_622), .B2(n_615), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g648 ( .A(n_629), .B(n_620), .C(n_621), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_627), .A2(n_598), .B1(n_600), .B2(n_605), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_637), .B(n_639), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_631), .B(n_604), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g652 ( .A1(n_632), .A2(n_618), .B1(n_607), .B2(n_228), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_638), .A2(n_244), .B(n_222), .C(n_228), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_630), .B(n_228), .Y(n_654) );
OA22x2_ASAP7_75t_L g655 ( .A1(n_641), .A2(n_626), .B1(n_633), .B2(n_611), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_632), .Y(n_656) );
OAI21xp33_ASAP7_75t_L g657 ( .A1(n_640), .A2(n_626), .B(n_635), .Y(n_657) );
NAND5xp2_ASAP7_75t_L g658 ( .A(n_657), .B(n_642), .C(n_643), .D(n_645), .E(n_648), .Y(n_658) );
XNOR2x1_ASAP7_75t_L g659 ( .A(n_655), .B(n_646), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_656), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_654), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_650), .B(n_644), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_658), .B(n_642), .C(n_651), .Y(n_663) );
AO21x1_ASAP7_75t_L g664 ( .A1(n_659), .A2(n_653), .B(n_649), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_660), .A2(n_655), .B(n_656), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_663), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_664), .A2(n_661), .B1(n_660), .B2(n_662), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_666), .B(n_665), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_667), .B1(n_652), .B2(n_647), .Y(n_669) );
UNKNOWN g670 ( );
endmodule