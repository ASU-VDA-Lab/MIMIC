module fake_netlist_1_4871_n_58 (n_11, n_1, n_2, n_13, n_16, n_12, n_6, n_4, n_3, n_9, n_17, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_58);
input n_11;
input n_1;
input n_2;
input n_13;
input n_16;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_17;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_58;
wire n_53;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_54;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_46;
wire n_48;
wire n_57;
wire n_25;
wire n_26;
wire n_30;
wire n_33;
wire n_50;
wire n_52;
wire n_49;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_55;
wire n_56;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_51;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
INVxp33_ASAP7_75t_SL g18 ( .A(n_3), .Y(n_18) );
INVx5_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_10), .B(n_11), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_16), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_8), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_15), .B(n_6), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_3), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_8), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_10), .B(n_7), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_20), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_19), .B(n_0), .Y(n_29) );
AO21x1_ASAP7_75t_L g30 ( .A1(n_21), .A2(n_0), .B(n_1), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_19), .B(n_1), .Y(n_31) );
AOI31xp67_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_22), .A3(n_26), .B(n_25), .Y(n_32) );
AOI21xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_27), .B(n_21), .Y(n_33) );
OAI21x1_ASAP7_75t_L g34 ( .A1(n_28), .A2(n_23), .B(n_27), .Y(n_34) );
INVxp67_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
HB1xp67_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
INVxp67_ASAP7_75t_SL g37 ( .A(n_35), .Y(n_37) );
AND2x2_ASAP7_75t_L g38 ( .A(n_36), .B(n_33), .Y(n_38) );
NOR2xp33_ASAP7_75t_L g39 ( .A(n_35), .B(n_18), .Y(n_39) );
AND2x4_ASAP7_75t_SL g40 ( .A(n_38), .B(n_28), .Y(n_40) );
NAND2x1p5_ASAP7_75t_L g41 ( .A(n_38), .B(n_19), .Y(n_41) );
AND2x2_ASAP7_75t_L g42 ( .A(n_38), .B(n_30), .Y(n_42) );
AOI31xp33_ASAP7_75t_SL g43 ( .A1(n_40), .A2(n_24), .A3(n_39), .B(n_30), .Y(n_43) );
AOI222xp33_ASAP7_75t_L g44 ( .A1(n_42), .A2(n_37), .B1(n_4), .B2(n_5), .C1(n_6), .C2(n_7), .Y(n_44) );
OAI21xp5_ASAP7_75t_SL g45 ( .A1(n_40), .A2(n_37), .B(n_4), .Y(n_45) );
AOI21xp33_ASAP7_75t_L g46 ( .A1(n_42), .A2(n_32), .B(n_5), .Y(n_46) );
NAND2xp5_ASAP7_75t_SL g47 ( .A(n_46), .B(n_41), .Y(n_47) );
XOR2xp5_ASAP7_75t_L g48 ( .A(n_43), .B(n_41), .Y(n_48) );
O2A1O1Ixp5_ASAP7_75t_SL g49 ( .A1(n_45), .A2(n_17), .B(n_9), .C(n_11), .Y(n_49) );
NOR3xp33_ASAP7_75t_L g50 ( .A(n_45), .B(n_2), .C(n_9), .Y(n_50) );
AND2x2_ASAP7_75t_L g51 ( .A(n_50), .B(n_44), .Y(n_51) );
NOR2xp33_ASAP7_75t_L g52 ( .A(n_48), .B(n_2), .Y(n_52) );
NAND3xp33_ASAP7_75t_SL g53 ( .A(n_49), .B(n_12), .C(n_13), .Y(n_53) );
NOR3xp33_ASAP7_75t_L g54 ( .A(n_47), .B(n_13), .C(n_14), .Y(n_54) );
NAND2xp5_ASAP7_75t_L g55 ( .A(n_51), .B(n_47), .Y(n_55) );
INVx1_ASAP7_75t_L g56 ( .A(n_53), .Y(n_56) );
OAI22xp33_ASAP7_75t_L g57 ( .A1(n_55), .A2(n_52), .B1(n_54), .B2(n_14), .Y(n_57) );
AOI22x1_ASAP7_75t_L g58 ( .A1(n_57), .A2(n_16), .B1(n_56), .B2(n_48), .Y(n_58) );
endmodule