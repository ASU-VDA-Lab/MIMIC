module fake_netlist_6_2893_n_1069 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1069);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1069;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_989;
wire n_843;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_939;
wire n_819;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_982;
wire n_831;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_249;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_882;
wire n_811;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_122),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_104),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_141),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_116),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_55),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_52),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_144),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_17),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_1),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_29),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_95),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_71),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_48),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_80),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_27),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_28),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_176),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_67),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_108),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_42),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_7),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_129),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_107),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_74),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_81),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_9),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_32),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_75),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_178),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_124),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_150),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_89),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_57),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_37),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_38),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_96),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_15),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_59),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_82),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_126),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_174),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_17),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_167),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_62),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_33),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_54),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_31),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_164),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_19),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_70),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_24),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_190),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_163),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_171),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_203),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_50),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_243),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_216),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_247),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_217),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_226),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_231),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_232),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_240),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_265),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_210),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_215),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_243),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_246),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_219),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_221),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_225),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_227),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_262),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_260),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_236),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_206),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_238),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_245),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_248),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_260),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_255),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_250),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_270),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_252),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_261),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_266),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_214),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_298),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_207),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_294),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

CKINVDCx11_ASAP7_75t_R g337 ( 
.A(n_298),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_273),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_325),
.B(n_246),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_208),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_274),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_281),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_323),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_305),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_289),
.B(n_272),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_277),
.B(n_209),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_297),
.B(n_212),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_285),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_290),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_286),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_305),
.B(n_213),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_290),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_291),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_291),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_278),
.B(n_220),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g366 ( 
.A(n_287),
.B(n_222),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_325),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_223),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_300),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_295),
.B(n_228),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_301),
.B(n_229),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_303),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_309),
.B(n_230),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_287),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_304),
.B(n_234),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_307),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_318),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_292),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_337),
.Y(n_380)
);

AO22x2_ASAP7_75t_L g381 ( 
.A1(n_328),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.Y(n_381)
);

BUFx10_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_369),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_327),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_378),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_375),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_319),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_379),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_282),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_373),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_379),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_320),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_R g394 ( 
.A(n_371),
.B(n_318),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_373),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_373),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_352),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_374),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_361),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_332),
.B(n_315),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_R g401 ( 
.A(n_366),
.B(n_321),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_368),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_R g403 ( 
.A(n_341),
.B(n_306),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_368),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_344),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_344),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_354),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_332),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_341),
.B(n_235),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_357),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_354),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_365),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_327),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_331),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_365),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_327),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_376),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_376),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_355),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_355),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_362),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_327),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_331),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_336),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_288),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_372),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_372),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_336),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_331),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_326),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_R g438 ( 
.A(n_353),
.B(n_306),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_326),
.B(n_272),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_326),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_326),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_362),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_340),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_340),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_340),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_336),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_340),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_439),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_414),
.A2(n_353),
.B1(n_345),
.B2(n_367),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_367),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_383),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_403),
.B(n_276),
.Y(n_453)
);

AO22x2_ASAP7_75t_L g454 ( 
.A1(n_414),
.A2(n_345),
.B1(n_363),
.B2(n_364),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_345),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_415),
.B(n_345),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_386),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_399),
.B(n_367),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_402),
.B(n_367),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_426),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_404),
.B(n_422),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_398),
.B(n_276),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_364),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_448),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_388),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_419),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_393),
.B(n_347),
.Y(n_470)
);

NAND3xp33_ASAP7_75t_L g471 ( 
.A(n_432),
.B(n_393),
.C(n_423),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_411),
.B(n_237),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_416),
.B(n_211),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_347),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_390),
.B(n_370),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_412),
.B(n_370),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_437),
.B(n_347),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_428),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_440),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_443),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_444),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_387),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_447),
.B(n_347),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_417),
.B(n_359),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_428),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_420),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_421),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_421),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_406),
.B(n_224),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_381),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_433),
.B(n_359),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_400),
.B(n_370),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_410),
.B(n_239),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_381),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_434),
.B(n_359),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_438),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_385),
.Y(n_501)
);

AND2x2_ASAP7_75t_SL g502 ( 
.A(n_446),
.B(n_377),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_381),
.B(n_377),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_430),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_418),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_435),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_R g509 ( 
.A(n_380),
.B(n_242),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_391),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_395),
.B(n_396),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_SL g514 ( 
.A(n_403),
.B(n_244),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_430),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_389),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_382),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_413),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_382),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_394),
.A2(n_249),
.B1(n_253),
.B2(n_254),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_436),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_397),
.B(n_377),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_392),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_401),
.B(n_359),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_401),
.B(n_348),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_464),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_468),
.B(n_360),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_466),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_459),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_348),
.Y(n_532)
);

OAI22xp33_ASAP7_75t_L g533 ( 
.A1(n_451),
.A2(n_394),
.B1(n_258),
.B2(n_259),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_465),
.B(n_263),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_491),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_524),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_467),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_466),
.Y(n_538)
);

AO22x2_ASAP7_75t_L g539 ( 
.A1(n_498),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_455),
.Y(n_540)
);

NAND3x1_ASAP7_75t_L g541 ( 
.A(n_492),
.B(n_360),
.C(n_334),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_468),
.A2(n_360),
.B1(n_329),
.B2(n_334),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_504),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_474),
.B(n_360),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_471),
.B(n_264),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_462),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_462),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_527),
.B(n_268),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_473),
.B(n_275),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_456),
.A2(n_329),
.B1(n_342),
.B2(n_346),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_470),
.B(n_349),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_475),
.B(n_356),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_501),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_509),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_524),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_501),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_495),
.B(n_356),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_502),
.B(n_349),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_502),
.B(n_349),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_507),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_513),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_503),
.A2(n_350),
.B1(n_342),
.B2(n_346),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_449),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_516),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_473),
.B(n_0),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_507),
.Y(n_567)
);

OAI221xp5_ASAP7_75t_L g568 ( 
.A1(n_493),
.A2(n_358),
.B1(n_343),
.B2(n_346),
.C(n_342),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_450),
.B(n_350),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_517),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_449),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_493),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_450),
.B(n_350),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_456),
.A2(n_346),
.B1(n_342),
.B2(n_343),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_460),
.B(n_350),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_500),
.B(n_358),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_460),
.B(n_350),
.Y(n_577)
);

NAND2x1p5_ASAP7_75t_L g578 ( 
.A(n_521),
.B(n_338),
.Y(n_578)
);

OAI221xp5_ASAP7_75t_L g579 ( 
.A1(n_485),
.A2(n_339),
.B1(n_335),
.B2(n_333),
.C(n_350),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_519),
.B(n_30),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_457),
.B(n_34),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_457),
.B(n_35),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_489),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_489),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_476),
.B(n_333),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_492),
.B(n_2),
.Y(n_586)
);

AO22x2_ASAP7_75t_L g587 ( 
.A1(n_461),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_461),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_588)
);

CKINVDCx10_ASAP7_75t_R g589 ( 
.A(n_531),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_552),
.B(n_494),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_558),
.B(n_549),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_540),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_534),
.B(n_499),
.Y(n_593)
);

AOI21x1_ASAP7_75t_L g594 ( 
.A1(n_575),
.A2(n_512),
.B(n_454),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_529),
.A2(n_486),
.B(n_478),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_504),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_543),
.B(n_463),
.Y(n_597)
);

AO21x1_ASAP7_75t_L g598 ( 
.A1(n_566),
.A2(n_526),
.B(n_514),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_529),
.A2(n_486),
.B(n_478),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_586),
.A2(n_463),
.B1(n_488),
.B2(n_480),
.Y(n_600)
);

O2A1O1Ixp5_ASAP7_75t_L g601 ( 
.A1(n_545),
.A2(n_514),
.B(n_477),
.C(n_484),
.Y(n_601)
);

CKINVDCx8_ASAP7_75t_R g602 ( 
.A(n_554),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_551),
.A2(n_496),
.B(n_458),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_551),
.A2(n_496),
.B(n_458),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_544),
.A2(n_505),
.B(n_476),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_533),
.A2(n_453),
.B1(n_481),
.B2(n_482),
.Y(n_606)
);

O2A1O1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_571),
.A2(n_472),
.B(n_497),
.C(n_479),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_537),
.B(n_469),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_546),
.B(n_527),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_548),
.A2(n_505),
.B(n_510),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_581),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_536),
.B(n_518),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_547),
.B(n_527),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_535),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_569),
.A2(n_454),
.B1(n_523),
.B2(n_525),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_571),
.B(n_452),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_556),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_564),
.B(n_497),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_530),
.A2(n_522),
.B(n_472),
.C(n_506),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_555),
.B(n_538),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_569),
.A2(n_454),
.B1(n_505),
.B2(n_515),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_562),
.B(n_527),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_573),
.A2(n_487),
.B1(n_490),
.B2(n_508),
.Y(n_623)
);

AOI21xp33_ASAP7_75t_L g624 ( 
.A1(n_528),
.A2(n_483),
.B(n_520),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_565),
.B(n_527),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_581),
.B(n_333),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_582),
.B(n_509),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_572),
.B(n_6),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_585),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_582),
.A2(n_532),
.B1(n_580),
.B2(n_541),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_553),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_532),
.B(n_36),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_570),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_580),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_575),
.B(n_335),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_583),
.B(n_338),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_559),
.B(n_339),
.Y(n_637)
);

O2A1O1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_568),
.A2(n_338),
.B(n_8),
.C(n_10),
.Y(n_638)
);

AO22x1_ASAP7_75t_L g639 ( 
.A1(n_584),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_577),
.A2(n_336),
.B(n_338),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_596),
.B(n_557),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_592),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_616),
.B(n_561),
.Y(n_643)
);

INVx6_ASAP7_75t_L g644 ( 
.A(n_611),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_611),
.B(n_567),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_618),
.B(n_587),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_617),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_611),
.B(n_577),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_602),
.B(n_578),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_600),
.B(n_578),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_593),
.A2(n_568),
.B(n_542),
.C(n_559),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_591),
.B(n_560),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_607),
.A2(n_550),
.B(n_574),
.C(n_560),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_597),
.A2(n_588),
.B1(n_587),
.B2(n_539),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_614),
.Y(n_655)
);

AO21x1_ASAP7_75t_L g656 ( 
.A1(n_615),
.A2(n_542),
.B(n_588),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_595),
.A2(n_579),
.B(n_563),
.Y(n_657)
);

AO32x2_ASAP7_75t_L g658 ( 
.A1(n_621),
.A2(n_588),
.A3(n_539),
.B1(n_579),
.B2(n_15),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_589),
.Y(n_659)
);

OA22x2_ASAP7_75t_L g660 ( 
.A1(n_606),
.A2(n_539),
.B1(n_13),
.B2(n_14),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_619),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_630),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_662)
);

BUFx4f_ASAP7_75t_L g663 ( 
.A(n_632),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_633),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_624),
.B(n_16),
.Y(n_665)
);

O2A1O1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_634),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_590),
.B(n_20),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_599),
.A2(n_40),
.B(n_39),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_608),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_627),
.B(n_21),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_601),
.A2(n_123),
.B(n_202),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_SL g672 ( 
.A1(n_628),
.A2(n_121),
.B(n_201),
.C(n_200),
.Y(n_672)
);

OAI21xp33_ASAP7_75t_L g673 ( 
.A1(n_612),
.A2(n_22),
.B(n_23),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_629),
.B(n_22),
.Y(n_674)
);

NAND2x1p5_ASAP7_75t_L g675 ( 
.A(n_632),
.B(n_41),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_605),
.A2(n_120),
.B(n_198),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_631),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_603),
.A2(n_118),
.B(n_196),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_620),
.Y(n_679)
);

OR2x6_ASAP7_75t_L g680 ( 
.A(n_639),
.B(n_43),
.Y(n_680)
);

A2O1A1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_622),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_681)
);

AOI21xp33_ASAP7_75t_L g682 ( 
.A1(n_625),
.A2(n_25),
.B(n_26),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_626),
.A2(n_26),
.B1(n_27),
.B2(n_44),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_604),
.A2(n_45),
.B(n_46),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_626),
.B(n_47),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_626),
.Y(n_686)
);

BUFx12f_ASAP7_75t_L g687 ( 
.A(n_636),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_610),
.A2(n_49),
.B(n_51),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_638),
.A2(n_53),
.B(n_56),
.C(n_58),
.Y(n_689)
);

OAI22x1_ASAP7_75t_L g690 ( 
.A1(n_594),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_690)
);

BUFx2_ASAP7_75t_SL g691 ( 
.A(n_598),
.Y(n_691)
);

NAND2x1p5_ASAP7_75t_L g692 ( 
.A(n_609),
.B(n_64),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_637),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_613),
.B(n_65),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_623),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_655),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_679),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_679),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_644),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_663),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_644),
.Y(n_701)
);

BUFx2_ASAP7_75t_SL g702 ( 
.A(n_659),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_687),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_645),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_646),
.B(n_641),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_645),
.B(n_640),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_667),
.B(n_66),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_669),
.Y(n_708)
);

BUFx4_ASAP7_75t_SL g709 ( 
.A(n_680),
.Y(n_709)
);

BUFx4f_ASAP7_75t_SL g710 ( 
.A(n_665),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_647),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_642),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_664),
.Y(n_713)
);

NAND2x1p5_ASAP7_75t_L g714 ( 
.A(n_686),
.B(n_635),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_677),
.Y(n_715)
);

CKINVDCx11_ASAP7_75t_R g716 ( 
.A(n_680),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_670),
.B(n_68),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_648),
.Y(n_718)
);

NAND2x1p5_ASAP7_75t_L g719 ( 
.A(n_650),
.B(n_635),
.Y(n_719)
);

CKINVDCx6p67_ASAP7_75t_R g720 ( 
.A(n_690),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_643),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_660),
.B(n_69),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_674),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_695),
.Y(n_724)
);

BUFx12f_ASAP7_75t_L g725 ( 
.A(n_675),
.Y(n_725)
);

BUFx2_ASAP7_75t_SL g726 ( 
.A(n_648),
.Y(n_726)
);

INVx8_ASAP7_75t_L g727 ( 
.A(n_649),
.Y(n_727)
);

NAND2x1p5_ASAP7_75t_L g728 ( 
.A(n_693),
.B(n_635),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_692),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_658),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_691),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_658),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_658),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_652),
.Y(n_734)
);

BUFx12f_ASAP7_75t_L g735 ( 
.A(n_683),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_685),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_662),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_656),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_694),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_666),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_654),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_676),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_661),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_671),
.Y(n_744)
);

BUFx4f_ASAP7_75t_SL g745 ( 
.A(n_672),
.Y(n_745)
);

BUFx6f_ASAP7_75t_SL g746 ( 
.A(n_673),
.Y(n_746)
);

AND2x6_ASAP7_75t_L g747 ( 
.A(n_681),
.B(n_72),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_653),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_682),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_668),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_678),
.Y(n_751)
);

INVx5_ASAP7_75t_SL g752 ( 
.A(n_688),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_684),
.Y(n_753)
);

INVx8_ASAP7_75t_L g754 ( 
.A(n_689),
.Y(n_754)
);

INVx5_ASAP7_75t_L g755 ( 
.A(n_651),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_657),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_698),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_699),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_756),
.A2(n_73),
.B(n_76),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_742),
.A2(n_77),
.B(n_78),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_734),
.B(n_79),
.Y(n_761)
);

OAI21x1_ASAP7_75t_L g762 ( 
.A1(n_742),
.A2(n_719),
.B(n_728),
.Y(n_762)
);

INVx6_ASAP7_75t_L g763 ( 
.A(n_700),
.Y(n_763)
);

AOI21xp33_ASAP7_75t_L g764 ( 
.A1(n_749),
.A2(n_83),
.B(n_84),
.Y(n_764)
);

OAI21x1_ASAP7_75t_L g765 ( 
.A1(n_719),
.A2(n_85),
.B(n_86),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_715),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_731),
.B(n_87),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_712),
.Y(n_768)
);

AO21x2_ASAP7_75t_L g769 ( 
.A1(n_744),
.A2(n_88),
.B(n_90),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_708),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_770)
);

AO21x2_ASAP7_75t_L g771 ( 
.A1(n_744),
.A2(n_94),
.B(n_97),
.Y(n_771)
);

OAI21x1_ASAP7_75t_L g772 ( 
.A1(n_728),
.A2(n_98),
.B(n_99),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_713),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_721),
.B(n_100),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_734),
.B(n_101),
.Y(n_775)
);

NOR2x1_ASAP7_75t_SL g776 ( 
.A(n_755),
.B(n_736),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_705),
.B(n_102),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_714),
.A2(n_103),
.B(n_105),
.Y(n_778)
);

OA21x2_ASAP7_75t_L g779 ( 
.A1(n_738),
.A2(n_106),
.B(n_109),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_724),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_702),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_R g782 ( 
.A(n_727),
.B(n_204),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_748),
.A2(n_756),
.B(n_743),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_714),
.A2(n_718),
.B(n_724),
.Y(n_784)
);

AO21x2_ASAP7_75t_L g785 ( 
.A1(n_738),
.A2(n_733),
.B(n_730),
.Y(n_785)
);

AO21x2_ASAP7_75t_L g786 ( 
.A1(n_732),
.A2(n_110),
.B(n_111),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_723),
.A2(n_112),
.B(n_113),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_708),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_746),
.A2(n_115),
.B1(n_117),
.B2(n_125),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_711),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_755),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_711),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_707),
.A2(n_127),
.B(n_128),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_752),
.A2(n_131),
.B(n_133),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_752),
.A2(n_134),
.B(n_135),
.Y(n_795)
);

AO32x2_ASAP7_75t_L g796 ( 
.A1(n_743),
.A2(n_136),
.A3(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_755),
.A2(n_140),
.B(n_142),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_721),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_731),
.B(n_149),
.Y(n_799)
);

INVx3_ASAP7_75t_SL g800 ( 
.A(n_727),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_711),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_741),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_696),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_726),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_710),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_805)
);

NOR2x1_ASAP7_75t_R g806 ( 
.A(n_716),
.B(n_154),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_701),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_749),
.B(n_155),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_737),
.A2(n_156),
.B(n_157),
.C(n_158),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_746),
.A2(n_195),
.B1(n_160),
.B2(n_161),
.Y(n_810)
);

OAI21x1_ASAP7_75t_L g811 ( 
.A1(n_752),
.A2(n_159),
.B(n_162),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_727),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_722),
.B(n_165),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_785),
.Y(n_814)
);

OAI221xp5_ASAP7_75t_SL g815 ( 
.A1(n_789),
.A2(n_717),
.B1(n_720),
.B2(n_739),
.C(n_709),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_768),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_773),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_788),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_785),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_780),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_800),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_783),
.B(n_754),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_791),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_766),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_784),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_786),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_791),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_783),
.B(n_755),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_800),
.Y(n_829)
);

AO21x1_ASAP7_75t_SL g830 ( 
.A1(n_797),
.A2(n_745),
.B(n_754),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_762),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_804),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_786),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_804),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_796),
.Y(n_835)
);

AO21x1_ASAP7_75t_SL g836 ( 
.A1(n_797),
.A2(n_745),
.B(n_754),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_796),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_779),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_796),
.B(n_706),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_779),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_772),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_802),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_765),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_769),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_760),
.A2(n_750),
.B(n_751),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_790),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_769),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_778),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_771),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_803),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_792),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_812),
.B(n_751),
.Y(n_852)
);

OR2x6_ASAP7_75t_L g853 ( 
.A(n_767),
.B(n_725),
.Y(n_853)
);

NOR2x1_ASAP7_75t_SL g854 ( 
.A(n_771),
.B(n_770),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_794),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_801),
.Y(n_856)
);

BUFx12f_ASAP7_75t_L g857 ( 
.A(n_758),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_850),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_854),
.A2(n_753),
.B(n_776),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_820),
.B(n_781),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_829),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_834),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_829),
.B(n_812),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_834),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_823),
.B(n_827),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_857),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_816),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_R g868 ( 
.A(n_853),
.B(n_782),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_857),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_832),
.Y(n_870)
);

NOR3xp33_ASAP7_75t_SL g871 ( 
.A(n_815),
.B(n_805),
.C(n_798),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_SL g872 ( 
.A(n_844),
.B(n_805),
.C(n_798),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_818),
.B(n_757),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_850),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_842),
.B(n_818),
.Y(n_875)
);

OR2x6_ASAP7_75t_L g876 ( 
.A(n_822),
.B(n_767),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_821),
.Y(n_877)
);

AO31x2_ASAP7_75t_L g878 ( 
.A1(n_854),
.A2(n_770),
.A3(n_759),
.B(n_761),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_830),
.A2(n_735),
.B1(n_747),
.B2(n_710),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_828),
.B(n_807),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_824),
.B(n_761),
.Y(n_881)
);

INVx8_ASAP7_75t_L g882 ( 
.A(n_853),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_828),
.B(n_799),
.Y(n_883)
);

BUFx4f_ASAP7_75t_SL g884 ( 
.A(n_821),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_816),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_837),
.A2(n_789),
.B1(n_810),
.B2(n_799),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_852),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_837),
.A2(n_810),
.B(n_759),
.C(n_809),
.Y(n_888)
);

AO31x2_ASAP7_75t_L g889 ( 
.A1(n_838),
.A2(n_775),
.A3(n_774),
.B(n_709),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_822),
.B(n_795),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_853),
.A2(n_793),
.B(n_809),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_817),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_817),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_R g894 ( 
.A(n_853),
.B(n_808),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_867),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_887),
.B(n_839),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_870),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_865),
.B(n_839),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_885),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_865),
.B(n_837),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_884),
.B(n_829),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_861),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_881),
.B(n_852),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_861),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_858),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_875),
.B(n_824),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_888),
.A2(n_822),
.B(n_764),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_862),
.B(n_825),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_864),
.B(n_814),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_878),
.B(n_825),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_883),
.B(n_851),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_892),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_893),
.B(n_880),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_860),
.B(n_837),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_889),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_873),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_873),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_889),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_897),
.B(n_889),
.Y(n_919)
);

AOI21xp33_ASAP7_75t_L g920 ( 
.A1(n_907),
.A2(n_894),
.B(n_886),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_909),
.Y(n_921)
);

OAI21x1_ASAP7_75t_L g922 ( 
.A1(n_915),
.A2(n_859),
.B(n_918),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_901),
.A2(n_891),
.B(n_876),
.Y(n_923)
);

OAI211xp5_ASAP7_75t_L g924 ( 
.A1(n_918),
.A2(n_872),
.B(n_871),
.C(n_879),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_905),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_900),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_905),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_906),
.A2(n_903),
.B(n_863),
.Y(n_928)
);

NAND4xp25_ASAP7_75t_L g929 ( 
.A(n_910),
.B(n_774),
.C(n_868),
.D(n_775),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_899),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_900),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_914),
.A2(n_830),
.B1(n_836),
.B2(n_837),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_909),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_925),
.B(n_882),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_930),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_926),
.B(n_898),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_925),
.Y(n_937)
);

AOI221xp5_ASAP7_75t_L g938 ( 
.A1(n_920),
.A2(n_914),
.B1(n_910),
.B2(n_913),
.C(n_911),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_921),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_921),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_922),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_931),
.Y(n_942)
);

NOR3xp33_ASAP7_75t_L g943 ( 
.A(n_924),
.B(n_806),
.C(n_866),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_929),
.B(n_910),
.C(n_764),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_937),
.B(n_928),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_935),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_937),
.B(n_919),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_939),
.B(n_933),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_934),
.B(n_936),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_942),
.B(n_933),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_934),
.B(n_916),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_939),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_947),
.B(n_940),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_952),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_949),
.B(n_943),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_945),
.B(n_927),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_946),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_951),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_950),
.B(n_944),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_954),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_956),
.B(n_938),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_954),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_957),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_953),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_955),
.B(n_948),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_958),
.B(n_948),
.Y(n_966)
);

INVxp67_ASAP7_75t_SL g967 ( 
.A(n_959),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_956),
.B(n_941),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_956),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_956),
.B(n_923),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_967),
.B(n_898),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_967),
.B(n_916),
.Y(n_972)
);

OAI322xp33_ASAP7_75t_L g973 ( 
.A1(n_963),
.A2(n_835),
.A3(n_849),
.B1(n_847),
.B2(n_844),
.C1(n_838),
.C2(n_877),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_969),
.B(n_869),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_960),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_960),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_962),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_965),
.B(n_874),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_975),
.A2(n_961),
.B(n_964),
.C(n_963),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_978),
.B(n_966),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_978),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_SL g982 ( 
.A1(n_974),
.A2(n_970),
.B(n_968),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_976),
.B(n_917),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_971),
.A2(n_972),
.B(n_977),
.Y(n_984)
);

OR2x6_ASAP7_75t_L g985 ( 
.A(n_973),
.B(n_703),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_983),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_979),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_981),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_980),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_984),
.B(n_917),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_988),
.B(n_982),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_989),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_990),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_986),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_987),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_988),
.B(n_985),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_993),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_991),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_996),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_995),
.B(n_910),
.Y(n_1000)
);

NAND4xp25_ASAP7_75t_L g1001 ( 
.A(n_992),
.B(n_994),
.C(n_932),
.D(n_813),
.Y(n_1001)
);

NAND4xp25_ASAP7_75t_SL g1002 ( 
.A(n_996),
.B(n_932),
.C(n_896),
.D(n_777),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_1002),
.A2(n_697),
.B(n_876),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_998),
.A2(n_703),
.B(n_882),
.Y(n_1004)
);

NOR2x1_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_703),
.Y(n_1005)
);

OAI32xp33_ASAP7_75t_L g1006 ( 
.A1(n_1000),
.A2(n_849),
.A3(n_847),
.B1(n_899),
.B2(n_843),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_SL g1007 ( 
.A(n_1004),
.B(n_997),
.C(n_1001),
.Y(n_1007)
);

AOI211xp5_ASAP7_75t_L g1008 ( 
.A1(n_1003),
.A2(n_700),
.B(n_811),
.C(n_904),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_SL g1009 ( 
.A1(n_1005),
.A2(n_895),
.B(n_912),
.C(n_169),
.Y(n_1009)
);

NOR2x1_ASAP7_75t_L g1010 ( 
.A(n_1006),
.B(n_700),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_1005),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1005),
.Y(n_1012)
);

OAI221xp5_ASAP7_75t_SL g1013 ( 
.A1(n_1003),
.A2(n_904),
.B1(n_902),
.B2(n_890),
.C(n_822),
.Y(n_1013)
);

OAI211xp5_ASAP7_75t_SL g1014 ( 
.A1(n_1005),
.A2(n_753),
.B(n_843),
.C(n_851),
.Y(n_1014)
);

OAI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_1011),
.A2(n_763),
.B1(n_902),
.B2(n_890),
.Y(n_1015)
);

XOR2xp5_ASAP7_75t_L g1016 ( 
.A(n_1007),
.B(n_166),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_1012),
.B(n_896),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_L g1018 ( 
.A(n_1009),
.B(n_1010),
.C(n_1008),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1013),
.B(n_912),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_1014),
.B(n_763),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_1011),
.Y(n_1021)
);

AOI311xp33_ASAP7_75t_L g1022 ( 
.A1(n_1009),
.A2(n_833),
.A3(n_826),
.B(n_820),
.C(n_819),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_1012),
.A2(n_704),
.B(n_895),
.C(n_843),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1011),
.Y(n_1024)
);

AO22x2_ASAP7_75t_L g1025 ( 
.A1(n_1024),
.A2(n_840),
.B1(n_856),
.B2(n_833),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1017),
.B(n_908),
.Y(n_1026)
);

AND3x4_ASAP7_75t_L g1027 ( 
.A(n_1016),
.B(n_763),
.C(n_729),
.Y(n_1027)
);

OAI221xp5_ASAP7_75t_L g1028 ( 
.A1(n_1018),
.A2(n_855),
.B1(n_841),
.B2(n_848),
.C(n_856),
.Y(n_1028)
);

AOI32xp33_ASAP7_75t_L g1029 ( 
.A1(n_1020),
.A2(n_787),
.A3(n_908),
.B1(n_841),
.B2(n_846),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_L g1030 ( 
.A(n_1019),
.B(n_841),
.C(n_846),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_1021),
.B(n_908),
.Y(n_1031)
);

OAI311xp33_ASAP7_75t_L g1032 ( 
.A1(n_1023),
.A2(n_846),
.A3(n_836),
.B1(n_740),
.C1(n_878),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1021),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_L g1034 ( 
.A(n_1015),
.B(n_168),
.C(n_170),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_1022),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_1021),
.B(n_908),
.Y(n_1036)
);

AOI221xp5_ASAP7_75t_SL g1037 ( 
.A1(n_1024),
.A2(n_855),
.B1(n_848),
.B2(n_831),
.C(n_826),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_1031),
.Y(n_1038)
);

CKINVDCx16_ASAP7_75t_R g1039 ( 
.A(n_1033),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1026),
.Y(n_1040)
);

AO22x2_ASAP7_75t_L g1041 ( 
.A1(n_1027),
.A2(n_840),
.B1(n_740),
.B2(n_831),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_1035),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_1036),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_1034),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_L g1045 ( 
.A(n_1030),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1037),
.B(n_878),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_1038),
.Y(n_1047)
);

XOR2xp5_ASAP7_75t_L g1048 ( 
.A(n_1039),
.B(n_1044),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1042),
.A2(n_1028),
.B1(n_1029),
.B2(n_1025),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1040),
.B(n_1025),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1043),
.Y(n_1051)
);

OA21x2_ASAP7_75t_L g1052 ( 
.A1(n_1046),
.A2(n_1032),
.B(n_845),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_1045),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_1047),
.Y(n_1054)
);

OA21x2_ASAP7_75t_L g1055 ( 
.A1(n_1050),
.A2(n_1051),
.B(n_1049),
.Y(n_1055)
);

AO21x1_ASAP7_75t_L g1056 ( 
.A1(n_1048),
.A2(n_1041),
.B(n_175),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1054),
.Y(n_1057)
);

AOI22x1_ASAP7_75t_L g1058 ( 
.A1(n_1057),
.A2(n_1053),
.B1(n_1041),
.B2(n_1055),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1058),
.Y(n_1059)
);

OAI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1059),
.A2(n_1052),
.B1(n_1056),
.B2(n_855),
.Y(n_1060)
);

AOI211xp5_ASAP7_75t_L g1061 ( 
.A1(n_1059),
.A2(n_173),
.B(n_177),
.C(n_179),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1060),
.A2(n_747),
.B(n_181),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1061),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1063),
.A2(n_855),
.B1(n_848),
.B2(n_747),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1062),
.A2(n_855),
.B1(n_747),
.B2(n_848),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_1065),
.A2(n_848),
.B1(n_182),
.B2(n_184),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1064),
.A2(n_180),
.B(n_185),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_SL g1068 ( 
.A1(n_1067),
.A2(n_1066),
.B1(n_187),
.B2(n_188),
.Y(n_1068)
);

AOI211xp5_ASAP7_75t_L g1069 ( 
.A1(n_1068),
.A2(n_186),
.B(n_189),
.C(n_191),
.Y(n_1069)
);


endmodule