module real_aes_6953_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g432 ( .A(n_0), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_1), .A2(n_136), .B(n_139), .C(n_142), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_2), .A2(n_162), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g548 ( .A(n_3), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_4), .B(n_185), .Y(n_208) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_5), .A2(n_162), .B(n_476), .Y(n_475) );
AND2x6_ASAP7_75t_L g136 ( .A(n_6), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g169 ( .A(n_7), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_8), .B(n_43), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_9), .A2(n_216), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_10), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g480 ( .A(n_11), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_12), .B(n_191), .Y(n_519) );
INVx1_ASAP7_75t_L g128 ( .A(n_13), .Y(n_128) );
INVx1_ASAP7_75t_L g531 ( .A(n_14), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_15), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_16), .A2(n_170), .B(n_180), .C(n_183), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_17), .B(n_185), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_18), .A2(n_451), .B1(n_452), .B2(n_453), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_18), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_19), .B(n_487), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_20), .B(n_162), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_21), .B(n_226), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_22), .A2(n_191), .B(n_192), .C(n_194), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_23), .B(n_185), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_24), .B(n_148), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_25), .A2(n_182), .B(n_183), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_26), .B(n_148), .Y(n_235) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_27), .Y(n_244) );
INVx1_ASAP7_75t_L g234 ( .A(n_28), .Y(n_234) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_29), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_30), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_31), .B(n_148), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g111 ( .A1(n_32), .A2(n_66), .B1(n_112), .B2(n_113), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_32), .Y(n_113) );
INVx1_ASAP7_75t_L g221 ( .A(n_33), .Y(n_221) );
INVx1_ASAP7_75t_L g470 ( .A(n_34), .Y(n_470) );
AOI222xp33_ASAP7_75t_SL g446 ( .A1(n_35), .A2(n_447), .B1(n_448), .B2(n_457), .C1(n_731), .C2(n_734), .Y(n_446) );
INVx2_ASAP7_75t_L g134 ( .A(n_36), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_37), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_38), .A2(n_191), .B(n_204), .C(n_206), .Y(n_203) );
INVxp67_ASAP7_75t_L g223 ( .A(n_39), .Y(n_223) );
CKINVDCx14_ASAP7_75t_R g202 ( .A(n_40), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_41), .A2(n_139), .B(n_233), .C(n_237), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_42), .A2(n_136), .B(n_139), .C(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g469 ( .A(n_44), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_45), .A2(n_150), .B(n_167), .C(n_168), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_46), .B(n_148), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_47), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_48), .Y(n_218) );
INVx1_ASAP7_75t_L g189 ( .A(n_49), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_50), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_51), .B(n_162), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_52), .A2(n_139), .B1(n_194), .B2(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_53), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_54), .Y(n_545) );
CKINVDCx14_ASAP7_75t_R g164 ( .A(n_55), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g109 ( .A1(n_56), .A2(n_110), .B1(n_111), .B2(n_114), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_56), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_57), .A2(n_167), .B(n_206), .C(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g477 ( .A(n_58), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_59), .Y(n_511) );
INVx1_ASAP7_75t_L g137 ( .A(n_60), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_61), .A2(n_79), .B1(n_454), .B2(n_455), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_61), .Y(n_455) );
INVx1_ASAP7_75t_L g127 ( .A(n_62), .Y(n_127) );
INVx1_ASAP7_75t_SL g205 ( .A(n_63), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_64), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_65), .B(n_185), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_66), .Y(n_112) );
INVx1_ASAP7_75t_L g247 ( .A(n_67), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_SL g486 ( .A1(n_68), .A2(n_206), .B(n_487), .C(n_488), .Y(n_486) );
INVxp67_ASAP7_75t_L g489 ( .A(n_69), .Y(n_489) );
INVx1_ASAP7_75t_L g444 ( .A(n_70), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_71), .A2(n_162), .B(n_163), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_72), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_73), .A2(n_162), .B(n_177), .Y(n_176) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_74), .A2(n_104), .B1(n_437), .B2(n_445), .C1(n_738), .C2(n_743), .Y(n_103) );
OAI22xp33_ASAP7_75t_SL g106 ( .A1(n_74), .A2(n_107), .B1(n_108), .B2(n_426), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_74), .Y(n_426) );
INVx1_ASAP7_75t_L g505 ( .A(n_75), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_76), .A2(n_216), .B(n_217), .Y(n_215) );
INVx1_ASAP7_75t_L g178 ( .A(n_77), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_78), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_79), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_80), .A2(n_136), .B(n_139), .C(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_81), .A2(n_162), .B(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g181 ( .A(n_82), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_83), .B(n_222), .Y(n_499) );
INVx2_ASAP7_75t_L g125 ( .A(n_84), .Y(n_125) );
INVx1_ASAP7_75t_L g143 ( .A(n_85), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_86), .B(n_487), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_87), .A2(n_136), .B(n_139), .C(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g429 ( .A(n_88), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g729 ( .A(n_88), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_88), .B(n_431), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_89), .A2(n_139), .B(n_246), .C(n_249), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_90), .B(n_124), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_91), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_92), .A2(n_136), .B(n_139), .C(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_93), .Y(n_523) );
INVx1_ASAP7_75t_L g485 ( .A(n_94), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_95), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_96), .B(n_222), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_97), .B(n_155), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_98), .B(n_155), .Y(n_532) );
INVx2_ASAP7_75t_L g193 ( .A(n_99), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_100), .B(n_444), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_101), .A2(n_162), .B(n_484), .Y(n_483) );
OAI22xp5_ASAP7_75t_SL g448 ( .A1(n_102), .A2(n_449), .B1(n_450), .B2(n_456), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_102), .Y(n_456) );
INVxp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_427), .B(n_434), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
XNOR2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_115), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_115), .A2(n_458), .B1(n_726), .B2(n_730), .Y(n_457) );
INVx2_ASAP7_75t_L g735 ( .A(n_115), .Y(n_735) );
OR2x2_ASAP7_75t_SL g115 ( .A(n_116), .B(n_381), .Y(n_115) );
NAND5xp2_ASAP7_75t_L g116 ( .A(n_117), .B(n_293), .C(n_331), .D(n_352), .E(n_369), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_265), .C(n_286), .Y(n_117) );
OAI221xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_197), .B1(n_228), .B2(n_252), .C(n_256), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_157), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_121), .B(n_254), .Y(n_273) );
OR2x2_ASAP7_75t_L g300 ( .A(n_121), .B(n_174), .Y(n_300) );
AND2x2_ASAP7_75t_L g314 ( .A(n_121), .B(n_174), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_121), .B(n_160), .Y(n_328) );
AND2x2_ASAP7_75t_L g366 ( .A(n_121), .B(n_330), .Y(n_366) );
AND2x2_ASAP7_75t_L g395 ( .A(n_121), .B(n_305), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_121), .B(n_277), .Y(n_412) );
INVx4_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g292 ( .A(n_122), .B(n_173), .Y(n_292) );
BUFx3_ASAP7_75t_L g317 ( .A(n_122), .Y(n_317) );
AND2x2_ASAP7_75t_L g346 ( .A(n_122), .B(n_174), .Y(n_346) );
AND3x2_ASAP7_75t_L g359 ( .A(n_122), .B(n_360), .C(n_361), .Y(n_359) );
AO21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_129), .B(n_152), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_123), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_123), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_123), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_124), .A2(n_161), .B(n_172), .Y(n_160) );
INVx2_ASAP7_75t_L g227 ( .A(n_124), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_124), .A2(n_131), .B(n_231), .C(n_232), .Y(n_230) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_124), .A2(n_526), .B(n_532), .Y(n_525) );
AND2x2_ASAP7_75t_SL g124 ( .A(n_125), .B(n_126), .Y(n_124) );
AND2x2_ASAP7_75t_L g156 ( .A(n_125), .B(n_126), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
OAI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_138), .Y(n_129) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_131), .A2(n_244), .B(n_245), .Y(n_243) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_131), .A2(n_171), .B1(n_467), .B2(n_471), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_131), .A2(n_505), .B(n_506), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_131), .A2(n_545), .B(n_546), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
AND2x4_ASAP7_75t_L g162 ( .A(n_132), .B(n_136), .Y(n_162) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g224 ( .A(n_133), .Y(n_224) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
INVx1_ASAP7_75t_L g195 ( .A(n_134), .Y(n_195) );
INVx1_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_135), .Y(n_146) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
INVx3_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
INVx1_ASAP7_75t_L g487 ( .A(n_135), .Y(n_487) );
INVx4_ASAP7_75t_SL g171 ( .A(n_136), .Y(n_171) );
BUFx3_ASAP7_75t_L g237 ( .A(n_136), .Y(n_237) );
INVx5_ASAP7_75t_L g165 ( .A(n_139), .Y(n_165) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx3_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_140), .Y(n_207) );
O2A1O1Ixp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_147), .C(n_149), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_144), .A2(n_149), .B(n_247), .C(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g468 ( .A1(n_145), .A2(n_146), .B1(n_469), .B2(n_470), .Y(n_468) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx4_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
INVx2_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
INVx4_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_149), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_149), .A2(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
INVx3_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_154), .B(n_239), .Y(n_238) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_154), .A2(n_243), .B(n_250), .Y(n_242) );
NOR2xp33_ASAP7_75t_SL g501 ( .A(n_154), .B(n_502), .Y(n_501) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_155), .A2(n_483), .B(n_490), .Y(n_482) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g214 ( .A(n_156), .Y(n_214) );
INVx1_ASAP7_75t_L g282 ( .A(n_157), .Y(n_282) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_173), .Y(n_157) );
AOI32xp33_ASAP7_75t_L g337 ( .A1(n_158), .A2(n_289), .A3(n_338), .B1(n_341), .B2(n_342), .Y(n_337) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g264 ( .A(n_159), .B(n_173), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_159), .B(n_292), .Y(n_335) );
AND2x2_ASAP7_75t_L g342 ( .A(n_159), .B(n_314), .Y(n_342) );
OR2x2_ASAP7_75t_L g348 ( .A(n_159), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_159), .B(n_303), .Y(n_373) );
OR2x2_ASAP7_75t_L g391 ( .A(n_159), .B(n_210), .Y(n_391) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g255 ( .A(n_160), .B(n_186), .Y(n_255) );
INVx2_ASAP7_75t_L g277 ( .A(n_160), .Y(n_277) );
OR2x2_ASAP7_75t_L g299 ( .A(n_160), .B(n_186), .Y(n_299) );
AND2x2_ASAP7_75t_L g304 ( .A(n_160), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_160), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g360 ( .A(n_160), .B(n_254), .Y(n_360) );
BUFx2_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_SL g163 ( .A1(n_164), .A2(n_165), .B(n_166), .C(n_171), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_SL g177 ( .A1(n_165), .A2(n_171), .B(n_178), .C(n_179), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g188 ( .A1(n_165), .A2(n_171), .B(n_189), .C(n_190), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_165), .A2(n_171), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_SL g217 ( .A1(n_165), .A2(n_171), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_165), .A2(n_171), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_165), .A2(n_171), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_165), .A2(n_171), .B(n_528), .C(n_529), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVx5_ASAP7_75t_L g222 ( .A(n_170), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_170), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_170), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g249 ( .A(n_171), .Y(n_249) );
INVx1_ASAP7_75t_SL g411 ( .A(n_173), .Y(n_411) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_186), .Y(n_173) );
INVx1_ASAP7_75t_SL g254 ( .A(n_174), .Y(n_254) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_174), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_174), .B(n_340), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_174), .B(n_277), .C(n_395), .Y(n_406) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_184), .Y(n_174) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_175), .A2(n_187), .B(n_196), .Y(n_186) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_175), .A2(n_200), .B(n_208), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_182), .B(n_193), .Y(n_192) );
OAI22xp33_ASAP7_75t_L g220 ( .A1(n_182), .A2(n_221), .B1(n_222), .B2(n_223), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_182), .B(n_531), .Y(n_530) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_185), .A2(n_475), .B(n_481), .Y(n_474) );
INVx2_ASAP7_75t_L g305 ( .A(n_186), .Y(n_305) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_186), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_191), .B(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g550 ( .A(n_194), .Y(n_550) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_209), .Y(n_197) );
INVx1_ASAP7_75t_L g341 ( .A(n_198), .Y(n_341) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g259 ( .A(n_199), .B(n_241), .Y(n_259) );
INVx2_ASAP7_75t_L g276 ( .A(n_199), .Y(n_276) );
AND2x2_ASAP7_75t_L g281 ( .A(n_199), .B(n_242), .Y(n_281) );
AND2x2_ASAP7_75t_L g296 ( .A(n_199), .B(n_229), .Y(n_296) );
AND2x2_ASAP7_75t_L g308 ( .A(n_199), .B(n_280), .Y(n_308) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_207), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_209), .B(n_324), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_209), .B(n_281), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_209), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_209), .B(n_275), .Y(n_403) );
BUFx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g240 ( .A(n_210), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_210), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g285 ( .A(n_210), .B(n_229), .Y(n_285) );
AND2x2_ASAP7_75t_L g311 ( .A(n_210), .B(n_241), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_210), .B(n_351), .Y(n_350) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_215), .B(n_225), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_212), .A2(n_270), .B(n_271), .Y(n_269) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_212), .A2(n_504), .B(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AOI21xp5_ASAP7_75t_SL g495 ( .A1(n_213), .A2(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_214), .A2(n_466), .B(n_472), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_214), .B(n_426), .Y(n_472) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_214), .A2(n_544), .B(n_551), .Y(n_543) );
INVx1_ASAP7_75t_L g270 ( .A(n_215), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_220), .B(n_224), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_222), .A2(n_234), .B(n_235), .C(n_236), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_222), .A2(n_548), .B(n_549), .C(n_550), .Y(n_547) );
INVx2_ASAP7_75t_L g236 ( .A(n_224), .Y(n_236) );
INVx1_ASAP7_75t_L g271 ( .A(n_225), .Y(n_271) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_227), .B(n_251), .Y(n_250) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_227), .A2(n_515), .B(n_522), .Y(n_514) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_240), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_229), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g275 ( .A(n_229), .B(n_276), .Y(n_275) );
INVx3_ASAP7_75t_SL g280 ( .A(n_229), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_229), .B(n_267), .Y(n_333) );
OR2x2_ASAP7_75t_L g343 ( .A(n_229), .B(n_269), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_229), .B(n_311), .Y(n_371) );
OR2x2_ASAP7_75t_L g401 ( .A(n_229), .B(n_241), .Y(n_401) );
AND2x2_ASAP7_75t_L g405 ( .A(n_229), .B(n_242), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_229), .B(n_281), .Y(n_418) );
AND2x2_ASAP7_75t_L g425 ( .A(n_229), .B(n_307), .Y(n_425) );
OR2x6_ASAP7_75t_L g229 ( .A(n_230), .B(n_238), .Y(n_229) );
INVx1_ASAP7_75t_SL g368 ( .A(n_240), .Y(n_368) );
AND2x2_ASAP7_75t_L g307 ( .A(n_241), .B(n_269), .Y(n_307) );
AND2x2_ASAP7_75t_L g321 ( .A(n_241), .B(n_276), .Y(n_321) );
AND2x2_ASAP7_75t_L g324 ( .A(n_241), .B(n_280), .Y(n_324) );
INVx1_ASAP7_75t_L g351 ( .A(n_241), .Y(n_351) );
INVx2_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_L g263 ( .A(n_242), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g422 ( .A1(n_253), .A2(n_299), .B(n_423), .C(n_424), .Y(n_422) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g329 ( .A(n_254), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_255), .B(n_272), .Y(n_287) );
AND2x2_ASAP7_75t_L g313 ( .A(n_255), .B(n_314), .Y(n_313) );
OAI21xp5_ASAP7_75t_SL g256 ( .A1(n_257), .A2(n_260), .B(n_264), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_258), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g284 ( .A(n_259), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_259), .B(n_280), .Y(n_325) );
AND2x2_ASAP7_75t_L g416 ( .A(n_259), .B(n_267), .Y(n_416) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g289 ( .A(n_263), .B(n_276), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_263), .B(n_274), .Y(n_290) );
OAI322xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_273), .A3(n_274), .B1(n_277), .B2(n_278), .C1(n_282), .C2(n_283), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_272), .Y(n_266) );
AND2x2_ASAP7_75t_L g377 ( .A(n_267), .B(n_289), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_267), .B(n_341), .Y(n_423) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g320 ( .A(n_269), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g386 ( .A(n_273), .B(n_299), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_274), .B(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_275), .B(n_307), .Y(n_364) );
AND2x2_ASAP7_75t_L g310 ( .A(n_276), .B(n_280), .Y(n_310) );
AND2x2_ASAP7_75t_L g318 ( .A(n_277), .B(n_319), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_277), .A2(n_356), .B(n_416), .C(n_417), .Y(n_415) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_278), .A2(n_291), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_280), .B(n_307), .Y(n_347) );
AND2x2_ASAP7_75t_L g353 ( .A(n_280), .B(n_321), .Y(n_353) );
AND2x2_ASAP7_75t_L g387 ( .A(n_280), .B(n_289), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_281), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_SL g397 ( .A(n_281), .Y(n_397) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_285), .A2(n_313), .B1(n_315), .B2(n_320), .Y(n_312) );
OAI22xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_288), .B1(n_290), .B2(n_291), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g322 ( .A1(n_287), .A2(n_323), .B1(n_325), .B2(n_326), .Y(n_322) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_292), .A2(n_394), .B1(n_396), .B2(n_398), .C(n_402), .Y(n_393) );
AOI211xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B(n_301), .C(n_322), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
OR2x2_ASAP7_75t_L g363 ( .A(n_299), .B(n_316), .Y(n_363) );
INVx1_ASAP7_75t_L g414 ( .A(n_299), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g301 ( .A1(n_300), .A2(n_302), .B1(n_306), .B2(n_309), .C(n_312), .Y(n_301) );
INVx2_ASAP7_75t_SL g356 ( .A(n_300), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g421 ( .A(n_303), .Y(n_421) );
AND2x2_ASAP7_75t_L g345 ( .A(n_304), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g330 ( .A(n_305), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g392 ( .A(n_308), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_316), .B(n_418), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_317), .Y(n_316) );
INVxp67_ASAP7_75t_L g361 ( .A(n_319), .Y(n_361) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_320), .A2(n_332), .B(n_334), .C(n_336), .Y(n_331) );
INVx1_ASAP7_75t_L g409 ( .A(n_323), .Y(n_409) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_327), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g340 ( .A(n_330), .Y(n_340) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI222xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_343), .B1(n_344), .B2(n_347), .C1(n_348), .C2(n_350), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g376 ( .A(n_340), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_343), .B(n_397), .Y(n_396) );
NAND2xp33_ASAP7_75t_SL g374 ( .A(n_344), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g349 ( .A(n_346), .Y(n_349) );
AND2x2_ASAP7_75t_L g413 ( .A(n_346), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g379 ( .A(n_349), .B(n_376), .Y(n_379) );
INVx1_ASAP7_75t_L g408 ( .A(n_350), .Y(n_408) );
AOI211xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B(n_357), .C(n_362), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_356), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
AOI322xp5_ASAP7_75t_L g407 ( .A1(n_359), .A2(n_387), .A3(n_392), .B1(n_408), .B2(n_409), .C1(n_410), .C2(n_413), .Y(n_407) );
AND2x2_ASAP7_75t_L g394 ( .A(n_360), .B(n_395), .Y(n_394) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_365), .B2(n_367), .Y(n_362) );
INVxp33_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_372), .B1(n_374), .B2(n_377), .C(n_378), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NAND5xp2_ASAP7_75t_L g381 ( .A(n_382), .B(n_393), .C(n_407), .D(n_415), .E(n_419), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_387), .B(n_388), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVxp33_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g419 ( .A1(n_395), .A2(n_420), .B(n_421), .C(n_422), .Y(n_419) );
AOI31xp33_ASAP7_75t_L g402 ( .A1(n_397), .A2(n_403), .A3(n_404), .B(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g420 ( .A(n_418), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_429), .Y(n_436) );
INVx1_ASAP7_75t_SL g742 ( .A(n_429), .Y(n_742) );
BUFx2_ASAP7_75t_L g745 ( .A(n_429), .Y(n_745) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_430), .B(n_729), .Y(n_733) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g728 ( .A(n_431), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_SL g740 ( .A(n_441), .B(n_443), .Y(n_740) );
OA21x2_ASAP7_75t_L g744 ( .A1(n_441), .A2(n_442), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
CKINVDCx14_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_459), .A2(n_726), .B1(n_735), .B2(n_736), .Y(n_734) );
AND3x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_651), .C(n_700), .Y(n_459) );
NOR3xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_558), .C(n_596), .Y(n_460) );
OAI222xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_491), .B1(n_533), .B2(n_539), .C1(n_553), .C2(n_556), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_473), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_463), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_463), .B(n_601), .Y(n_692) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g569 ( .A(n_464), .B(n_482), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_464), .B(n_474), .Y(n_577) );
AND2x2_ASAP7_75t_L g612 ( .A(n_464), .B(n_589), .Y(n_612) );
OR2x2_ASAP7_75t_L g636 ( .A(n_464), .B(n_474), .Y(n_636) );
OR2x2_ASAP7_75t_L g644 ( .A(n_464), .B(n_543), .Y(n_644) );
AND2x2_ASAP7_75t_L g647 ( .A(n_464), .B(n_482), .Y(n_647) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g541 ( .A(n_465), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g555 ( .A(n_465), .B(n_482), .Y(n_555) );
AND2x2_ASAP7_75t_L g605 ( .A(n_465), .B(n_543), .Y(n_605) );
AND2x2_ASAP7_75t_L g618 ( .A(n_465), .B(n_474), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_465), .B(n_704), .Y(n_725) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_473), .A2(n_644), .B(n_645), .C(n_648), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_473), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_473), .B(n_588), .Y(n_710) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .Y(n_473) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_474), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g568 ( .A(n_474), .Y(n_568) );
AND2x2_ASAP7_75t_L g595 ( .A(n_474), .B(n_589), .Y(n_595) );
INVx1_ASAP7_75t_SL g603 ( .A(n_474), .Y(n_603) );
AND2x2_ASAP7_75t_L g626 ( .A(n_474), .B(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g704 ( .A(n_474), .Y(n_704) );
BUFx2_ASAP7_75t_L g540 ( .A(n_482), .Y(n_540) );
INVx1_ASAP7_75t_L g602 ( .A(n_482), .Y(n_602) );
INVx3_ASAP7_75t_L g627 ( .A(n_482), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_491), .B(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_512), .Y(n_491) );
INVx1_ASAP7_75t_L g623 ( .A(n_492), .Y(n_623) );
OAI32xp33_ASAP7_75t_L g629 ( .A1(n_492), .A2(n_568), .A3(n_630), .B1(n_631), .B2(n_632), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_492), .A2(n_634), .B1(n_637), .B2(n_642), .Y(n_633) );
INVx4_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g571 ( .A(n_493), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g649 ( .A(n_493), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g719 ( .A(n_493), .B(n_665), .Y(n_719) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
AND2x2_ASAP7_75t_L g534 ( .A(n_494), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g564 ( .A(n_494), .Y(n_564) );
INVx1_ASAP7_75t_L g583 ( .A(n_494), .Y(n_583) );
OR2x2_ASAP7_75t_L g591 ( .A(n_494), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g598 ( .A(n_494), .B(n_572), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_494), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g619 ( .A(n_494), .B(n_537), .Y(n_619) );
INVx3_ASAP7_75t_L g641 ( .A(n_494), .Y(n_641) );
AND2x2_ASAP7_75t_L g666 ( .A(n_494), .B(n_538), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_494), .B(n_631), .Y(n_714) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_501), .Y(n_494) );
INVx2_ASAP7_75t_L g538 ( .A(n_503), .Y(n_538) );
AND2x2_ASAP7_75t_L g670 ( .A(n_503), .B(n_513), .Y(n_670) );
INVx2_ASAP7_75t_L g712 ( .A(n_512), .Y(n_712) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .Y(n_512) );
INVx1_ASAP7_75t_L g557 ( .A(n_513), .Y(n_557) );
AND2x2_ASAP7_75t_L g584 ( .A(n_513), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_513), .B(n_538), .Y(n_592) );
AND2x2_ASAP7_75t_L g650 ( .A(n_513), .B(n_573), .Y(n_650) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g536 ( .A(n_514), .Y(n_536) );
AND2x2_ASAP7_75t_L g563 ( .A(n_514), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g572 ( .A(n_514), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_514), .B(n_538), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_521), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_524), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g585 ( .A(n_524), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_524), .B(n_538), .Y(n_631) );
AND2x2_ASAP7_75t_L g640 ( .A(n_524), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g665 ( .A(n_524), .Y(n_665) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g537 ( .A(n_525), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g573 ( .A(n_525), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_533), .A2(n_543), .B1(n_702), .B2(n_705), .Y(n_701) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
OAI21xp5_ASAP7_75t_SL g724 ( .A1(n_535), .A2(n_646), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_536), .B(n_641), .Y(n_658) );
INVx1_ASAP7_75t_L g683 ( .A(n_536), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_537), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g610 ( .A(n_537), .B(n_563), .Y(n_610) );
INVx2_ASAP7_75t_L g566 ( .A(n_538), .Y(n_566) );
INVx1_ASAP7_75t_L g616 ( .A(n_538), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_539), .A2(n_691), .B1(n_708), .B2(n_711), .C(n_713), .Y(n_707) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx1_ASAP7_75t_L g578 ( .A(n_540), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_540), .B(n_589), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_541), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g632 ( .A(n_541), .B(n_578), .Y(n_632) );
INVx3_ASAP7_75t_SL g673 ( .A(n_541), .Y(n_673) );
AND2x2_ASAP7_75t_L g617 ( .A(n_542), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g646 ( .A(n_542), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_542), .B(n_555), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_542), .B(n_601), .Y(n_687) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g589 ( .A(n_543), .Y(n_589) );
OAI322xp33_ASAP7_75t_L g684 ( .A1(n_543), .A2(n_615), .A3(n_637), .B1(n_685), .B2(n_687), .C1(n_688), .C2(n_689), .Y(n_684) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_554), .A2(n_557), .B(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_SL g634 ( .A(n_555), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g656 ( .A(n_555), .B(n_568), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_555), .B(n_595), .Y(n_671) );
INVxp67_ASAP7_75t_L g622 ( .A(n_557), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_557), .A2(n_629), .B(n_633), .C(n_643), .Y(n_628) );
OAI221xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_567), .B1(n_570), .B2(n_574), .C(n_579), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g582 ( .A(n_566), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g699 ( .A(n_566), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g715 ( .A1(n_567), .A2(n_716), .B1(n_721), .B2(n_722), .C(n_724), .Y(n_715) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_568), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g615 ( .A(n_568), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_568), .B(n_646), .Y(n_653) );
AND2x2_ASAP7_75t_L g695 ( .A(n_568), .B(n_673), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_569), .B(n_594), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_569), .A2(n_581), .B1(n_691), .B2(n_692), .Y(n_690) );
OR2x2_ASAP7_75t_L g721 ( .A(n_569), .B(n_589), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g698 ( .A(n_572), .Y(n_698) );
AND2x2_ASAP7_75t_L g723 ( .A(n_572), .B(n_666), .Y(n_723) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_SL g575 ( .A(n_576), .B(n_578), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g587 ( .A(n_577), .B(n_588), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_586), .B1(n_590), .B2(n_593), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
INVx1_ASAP7_75t_L g654 ( .A(n_582), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_582), .B(n_622), .Y(n_689) );
AOI322xp5_ASAP7_75t_L g613 ( .A1(n_584), .A2(n_614), .A3(n_616), .B1(n_617), .B2(n_619), .C1(n_620), .C2(n_624), .Y(n_613) );
INVxp67_ASAP7_75t_L g607 ( .A(n_585), .Y(n_607) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_587), .A2(n_592), .B1(n_609), .B2(n_611), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_588), .B(n_601), .Y(n_688) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_589), .B(n_627), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_589), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g685 ( .A(n_591), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
NAND3xp33_ASAP7_75t_SL g596 ( .A(n_597), .B(n_613), .C(n_628), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_604), .B2(n_606), .C(n_608), .Y(n_597) );
AND2x2_ASAP7_75t_L g604 ( .A(n_600), .B(n_605), .Y(n_604) );
INVx3_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g614 ( .A(n_605), .B(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_607), .Y(n_686) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_612), .B(n_626), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_615), .B(n_673), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_616), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g691 ( .A(n_619), .Y(n_691) );
AND2x2_ASAP7_75t_L g706 ( .A(n_619), .B(n_683), .Y(n_706) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g700 ( .A1(n_630), .A2(n_701), .B(n_707), .C(n_715), .Y(n_700) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g669 ( .A(n_640), .B(n_670), .Y(n_669) );
NAND2x1_ASAP7_75t_SL g711 ( .A(n_641), .B(n_712), .Y(n_711) );
CKINVDCx16_ASAP7_75t_R g681 ( .A(n_644), .Y(n_681) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g676 ( .A(n_650), .Y(n_676) );
AND2x2_ASAP7_75t_L g680 ( .A(n_650), .B(n_666), .Y(n_680) );
NOR5xp2_ASAP7_75t_L g651 ( .A(n_652), .B(n_667), .C(n_684), .D(n_690), .E(n_693), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B1(n_655), .B2(n_657), .C(n_659), .Y(n_652) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_656), .B(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g682 ( .A(n_666), .B(n_683), .Y(n_682) );
OAI221xp5_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_671), .B1(n_672), .B2(n_674), .C(n_677), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B1(n_681), .B2(n_682), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g720 ( .A(n_680), .Y(n_720) );
AOI211xp5_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_696), .B(n_698), .C(n_699), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
CKINVDCx14_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g737 ( .A(n_730), .Y(n_737) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
NAND2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
endmodule