module real_aes_7549_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_691;
wire n_481;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g421 ( .A(n_0), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_1), .A2(n_127), .B(n_132), .C(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g239 ( .A(n_2), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_3), .A2(n_122), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_4), .B(n_199), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g200 ( .A1(n_5), .A2(n_122), .B(n_201), .Y(n_200) );
AND2x6_ASAP7_75t_L g127 ( .A(n_6), .B(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g120 ( .A1(n_7), .A2(n_121), .B(n_129), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_8), .B(n_40), .Y(n_422) );
INVx1_ASAP7_75t_L g540 ( .A(n_9), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_10), .B(n_171), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_11), .B(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g206 ( .A(n_12), .Y(n_206) );
INVx1_ASAP7_75t_L g119 ( .A(n_13), .Y(n_119) );
INVx1_ASAP7_75t_L g139 ( .A(n_14), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_15), .A2(n_140), .B(n_154), .C(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_16), .B(n_199), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_17), .B(n_156), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_18), .B(n_122), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_19), .B(n_464), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_20), .A2(n_187), .B(n_213), .C(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_21), .B(n_199), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_22), .B(n_171), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_23), .A2(n_136), .B(n_138), .C(n_140), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_24), .B(n_171), .Y(n_437) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_25), .Y(n_468) );
INVx1_ASAP7_75t_L g436 ( .A(n_26), .Y(n_436) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_27), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_28), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_29), .B(n_171), .Y(n_240) );
INVx1_ASAP7_75t_L g461 ( .A(n_30), .Y(n_461) );
INVx1_ASAP7_75t_L g218 ( .A(n_31), .Y(n_218) );
INVx2_ASAP7_75t_L g125 ( .A(n_32), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_33), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_34), .A2(n_187), .B(n_207), .C(n_449), .Y(n_448) );
INVxp67_ASAP7_75t_L g462 ( .A(n_35), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_36), .A2(n_127), .B(n_132), .C(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_37), .A2(n_132), .B(n_435), .C(n_440), .Y(n_434) );
CKINVDCx14_ASAP7_75t_R g447 ( .A(n_38), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_39), .A2(n_66), .B1(n_104), .B2(n_105), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_39), .Y(n_104) );
INVx1_ASAP7_75t_L g216 ( .A(n_41), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_42), .A2(n_158), .B(n_204), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_43), .B(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g708 ( .A1(n_44), .A2(n_83), .B1(n_709), .B2(n_710), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_44), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_45), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_46), .Y(n_458) );
INVx1_ASAP7_75t_L g506 ( .A(n_47), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_48), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_49), .B(n_122), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_50), .A2(n_132), .B1(n_213), .B2(n_215), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_51), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_52), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_53), .A2(n_204), .B(n_205), .C(n_207), .Y(n_203) );
CKINVDCx14_ASAP7_75t_R g537 ( .A(n_54), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_55), .Y(n_175) );
INVx1_ASAP7_75t_L g202 ( .A(n_56), .Y(n_202) );
AOI222xp33_ASAP7_75t_SL g102 ( .A1(n_57), .A2(n_103), .B1(n_106), .B2(n_690), .C1(n_691), .C2(n_692), .Y(n_102) );
INVx1_ASAP7_75t_L g128 ( .A(n_58), .Y(n_128) );
INVx1_ASAP7_75t_L g118 ( .A(n_59), .Y(n_118) );
INVx1_ASAP7_75t_SL g450 ( .A(n_60), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_61), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_62), .B(n_199), .Y(n_510) );
INVx1_ASAP7_75t_L g471 ( .A(n_63), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_SL g226 ( .A1(n_64), .A2(n_156), .B(n_207), .C(n_227), .Y(n_226) );
INVxp67_ASAP7_75t_L g228 ( .A(n_65), .Y(n_228) );
INVx1_ASAP7_75t_L g105 ( .A(n_66), .Y(n_105) );
INVx1_ASAP7_75t_L g700 ( .A(n_67), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_68), .A2(n_122), .B(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_69), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_70), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_71), .A2(n_122), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g166 ( .A(n_72), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_73), .A2(n_121), .B(n_457), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g433 ( .A(n_74), .Y(n_433) );
INVx1_ASAP7_75t_L g498 ( .A(n_75), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_76), .A2(n_127), .B(n_132), .C(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_77), .A2(n_122), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g501 ( .A(n_78), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_79), .B(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g116 ( .A(n_80), .Y(n_116) );
INVx1_ASAP7_75t_L g490 ( .A(n_81), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_82), .B(n_156), .Y(n_155) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_83), .A2(n_101), .B1(n_696), .B2(n_705), .C1(n_715), .C2(n_721), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_83), .Y(n_709) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_84), .A2(n_127), .B(n_132), .C(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g419 ( .A(n_85), .Y(n_419) );
OR2x2_ASAP7_75t_L g689 ( .A(n_85), .B(n_420), .Y(n_689) );
OR2x2_ASAP7_75t_L g704 ( .A(n_85), .B(n_695), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_86), .A2(n_132), .B(n_470), .C(n_474), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_87), .B(n_115), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_88), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_89), .A2(n_127), .B(n_132), .C(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_90), .Y(n_192) );
INVx1_ASAP7_75t_L g225 ( .A(n_91), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g130 ( .A(n_92), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_93), .B(n_153), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_94), .B(n_144), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_95), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_96), .A2(n_122), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g509 ( .A(n_97), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_98), .B(n_700), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_99), .Y(n_714) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g690 ( .A(n_103), .Y(n_690) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_416), .B1(n_423), .B2(n_687), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
OAI22xp5_ASAP7_75t_SL g691 ( .A1(n_108), .A2(n_418), .B1(n_424), .B2(n_689), .Y(n_691) );
OR4x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_312), .C(n_371), .D(n_398), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_254), .C(n_279), .Y(n_109) );
O2A1O1Ixp33_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_177), .B(n_197), .C(n_230), .Y(n_110) );
AOI211xp5_ASAP7_75t_SL g402 ( .A1(n_111), .A2(n_403), .B(n_405), .C(n_408), .Y(n_402) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_146), .Y(n_111) );
INVx1_ASAP7_75t_L g277 ( .A(n_112), .Y(n_277) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g252 ( .A(n_113), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g284 ( .A(n_113), .Y(n_284) );
AND2x2_ASAP7_75t_L g339 ( .A(n_113), .B(n_308), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_113), .B(n_195), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_113), .B(n_196), .Y(n_397) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g258 ( .A(n_114), .Y(n_258) );
AND2x2_ASAP7_75t_L g301 ( .A(n_114), .B(n_164), .Y(n_301) );
AND2x2_ASAP7_75t_L g319 ( .A(n_114), .B(n_196), .Y(n_319) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_143), .Y(n_114) );
INVx1_ASAP7_75t_L g176 ( .A(n_115), .Y(n_176) );
INVx2_ASAP7_75t_L g181 ( .A(n_115), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g432 ( .A1(n_115), .A2(n_167), .B(n_433), .C(n_434), .Y(n_432) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_115), .A2(n_535), .B(n_541), .Y(n_534) );
AND2x2_ASAP7_75t_SL g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AND2x2_ASAP7_75t_L g145 ( .A(n_116), .B(n_117), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_127), .Y(n_122) );
NAND2x1p5_ASAP7_75t_L g167 ( .A(n_123), .B(n_127), .Y(n_167) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g439 ( .A(n_124), .Y(n_439) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g133 ( .A(n_125), .Y(n_133) );
INVx1_ASAP7_75t_L g214 ( .A(n_125), .Y(n_214) );
INVx1_ASAP7_75t_L g134 ( .A(n_126), .Y(n_134) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_126), .Y(n_137) );
INVx3_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
INVx1_ASAP7_75t_L g156 ( .A(n_126), .Y(n_156) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_126), .Y(n_171) );
INVx4_ASAP7_75t_SL g142 ( .A(n_127), .Y(n_142) );
BUFx3_ASAP7_75t_L g440 ( .A(n_127), .Y(n_440) );
O2A1O1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_135), .C(n_142), .Y(n_129) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_131), .A2(n_142), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_131), .A2(n_142), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_131), .A2(n_142), .B(n_447), .C(n_448), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_SL g457 ( .A1(n_131), .A2(n_142), .B(n_458), .C(n_459), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g497 ( .A1(n_131), .A2(n_142), .B(n_498), .C(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_131), .A2(n_142), .B(n_506), .C(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_131), .A2(n_142), .B(n_537), .C(n_538), .Y(n_536) );
INVx5_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx3_ASAP7_75t_L g141 ( .A(n_133), .Y(n_141) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_133), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_136), .B(n_139), .Y(n_138) );
OAI22xp33_ASAP7_75t_L g460 ( .A1(n_136), .A2(n_153), .B1(n_461), .B2(n_462), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_136), .B(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_136), .B(n_509), .Y(n_508) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OAI22xp5_ASAP7_75t_SL g215 ( .A1(n_137), .A2(n_216), .B1(n_217), .B2(n_218), .Y(n_215) );
INVx2_ASAP7_75t_L g217 ( .A(n_137), .Y(n_217) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
OAI22xp33_ASAP7_75t_L g211 ( .A1(n_142), .A2(n_167), .B1(n_212), .B2(n_219), .Y(n_211) );
INVx1_ASAP7_75t_L g474 ( .A(n_142), .Y(n_474) );
INVx4_ASAP7_75t_L g163 ( .A(n_144), .Y(n_163) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_144), .A2(n_223), .B(n_229), .Y(n_222) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_144), .Y(n_444) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g160 ( .A(n_145), .Y(n_160) );
INVx4_ASAP7_75t_L g251 ( .A(n_146), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_146), .A2(n_307), .B(n_309), .Y(n_306) );
AND2x2_ASAP7_75t_L g387 ( .A(n_146), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_164), .Y(n_146) );
INVx1_ASAP7_75t_L g194 ( .A(n_147), .Y(n_194) );
AND2x2_ASAP7_75t_L g256 ( .A(n_147), .B(n_196), .Y(n_256) );
OR2x2_ASAP7_75t_L g285 ( .A(n_147), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g299 ( .A(n_147), .Y(n_299) );
INVx3_ASAP7_75t_L g308 ( .A(n_147), .Y(n_308) );
AND2x2_ASAP7_75t_L g318 ( .A(n_147), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g351 ( .A(n_147), .B(n_257), .Y(n_351) );
AND2x2_ASAP7_75t_L g375 ( .A(n_147), .B(n_331), .Y(n_375) );
OR2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_161), .Y(n_147) );
AOI21xp5_ASAP7_75t_SL g148 ( .A1(n_149), .A2(n_150), .B(n_159), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_155), .B(n_157), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_153), .A2(n_239), .B(n_240), .C(n_241), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g435 ( .A1(n_153), .A2(n_436), .B(n_437), .C(n_438), .Y(n_435) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_154), .B(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_154), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_154), .B(n_540), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_157), .A2(n_170), .B(n_172), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_157), .A2(n_471), .B(n_472), .C(n_473), .Y(n_470) );
O2A1O1Ixp5_ASAP7_75t_L g489 ( .A1(n_157), .A2(n_472), .B(n_490), .C(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g173 ( .A(n_159), .Y(n_173) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_160), .A2(n_211), .B(n_220), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_160), .B(n_221), .Y(n_220) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_160), .A2(n_235), .B(n_242), .Y(n_234) );
NOR2xp33_ASAP7_75t_SL g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx3_ASAP7_75t_L g199 ( .A(n_163), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_163), .B(n_442), .Y(n_441) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_163), .A2(n_467), .B(n_475), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_163), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g196 ( .A(n_164), .Y(n_196) );
AND2x2_ASAP7_75t_L g411 ( .A(n_164), .B(n_253), .Y(n_411) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_173), .B(n_174), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_168), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_167), .A2(n_236), .B(n_237), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_167), .A2(n_468), .B(n_469), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_167), .A2(n_487), .B(n_488), .Y(n_486) );
INVx4_ASAP7_75t_L g187 ( .A(n_171), .Y(n_187) );
INVx2_ASAP7_75t_L g204 ( .A(n_171), .Y(n_204) );
INVx1_ASAP7_75t_L g455 ( .A(n_173), .Y(n_455) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_173), .A2(n_480), .B(n_481), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_176), .B(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_176), .B(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_176), .A2(n_486), .B(n_492), .Y(n_485) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_179), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g331 ( .A(n_179), .B(n_319), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_179), .B(n_308), .Y(n_393) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g253 ( .A(n_180), .Y(n_253) );
AND2x2_ASAP7_75t_L g257 ( .A(n_180), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g298 ( .A(n_180), .B(n_299), .Y(n_298) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_191), .Y(n_180) );
INVx1_ASAP7_75t_L g464 ( .A(n_181), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_181), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_190), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_187), .B(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g207 ( .A(n_189), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_193), .B(n_294), .Y(n_316) );
INVx1_ASAP7_75t_L g355 ( .A(n_193), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_193), .B(n_282), .Y(n_399) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AND2x2_ASAP7_75t_L g262 ( .A(n_194), .B(n_257), .Y(n_262) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_196), .B(n_253), .Y(n_286) );
INVx1_ASAP7_75t_L g365 ( .A(n_196), .Y(n_365) );
AOI322xp5_ASAP7_75t_L g389 ( .A1(n_197), .A2(n_304), .A3(n_364), .B1(n_390), .B2(n_392), .C1(n_394), .C2(n_396), .Y(n_389) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_198), .B(n_209), .Y(n_197) );
AND2x2_ASAP7_75t_L g244 ( .A(n_198), .B(n_222), .Y(n_244) );
INVx1_ASAP7_75t_SL g247 ( .A(n_198), .Y(n_247) );
AND2x2_ASAP7_75t_L g249 ( .A(n_198), .B(n_210), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_198), .B(n_266), .Y(n_272) );
INVx2_ASAP7_75t_L g291 ( .A(n_198), .Y(n_291) );
AND2x2_ASAP7_75t_L g304 ( .A(n_198), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g342 ( .A(n_198), .B(n_266), .Y(n_342) );
BUFx2_ASAP7_75t_L g359 ( .A(n_198), .Y(n_359) );
AND2x2_ASAP7_75t_L g373 ( .A(n_198), .B(n_233), .Y(n_373) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_208), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_209), .B(n_261), .Y(n_288) );
AND2x2_ASAP7_75t_L g415 ( .A(n_209), .B(n_291), .Y(n_415) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_222), .Y(n_209) );
OR2x2_ASAP7_75t_L g260 ( .A(n_210), .B(n_261), .Y(n_260) );
INVx3_ASAP7_75t_L g266 ( .A(n_210), .Y(n_266) );
AND2x2_ASAP7_75t_L g311 ( .A(n_210), .B(n_234), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_210), .B(n_359), .Y(n_358) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_210), .Y(n_395) );
INVx2_ASAP7_75t_L g241 ( .A(n_213), .Y(n_241) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g472 ( .A(n_217), .Y(n_472) );
AND2x2_ASAP7_75t_L g246 ( .A(n_222), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g268 ( .A(n_222), .Y(n_268) );
BUFx2_ASAP7_75t_L g274 ( .A(n_222), .Y(n_274) );
AND2x2_ASAP7_75t_L g293 ( .A(n_222), .B(n_266), .Y(n_293) );
INVx3_ASAP7_75t_L g305 ( .A(n_222), .Y(n_305) );
OR2x2_ASAP7_75t_L g315 ( .A(n_222), .B(n_266), .Y(n_315) );
AOI31xp33_ASAP7_75t_SL g230 ( .A1(n_231), .A2(n_245), .A3(n_248), .B(n_250), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_244), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_232), .B(n_267), .Y(n_278) );
OR2x2_ASAP7_75t_L g302 ( .A(n_232), .B(n_272), .Y(n_302) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_233), .B(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g323 ( .A(n_233), .B(n_315), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_233), .B(n_305), .Y(n_333) );
AND2x2_ASAP7_75t_L g340 ( .A(n_233), .B(n_341), .Y(n_340) );
NAND2x1_ASAP7_75t_L g368 ( .A(n_233), .B(n_304), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_233), .B(n_359), .Y(n_369) );
AND2x2_ASAP7_75t_L g381 ( .A(n_233), .B(n_266), .Y(n_381) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx3_ASAP7_75t_L g261 ( .A(n_234), .Y(n_261) );
INVx1_ASAP7_75t_L g327 ( .A(n_244), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_244), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_246), .B(n_322), .Y(n_356) );
AND2x4_ASAP7_75t_L g267 ( .A(n_247), .B(n_268), .Y(n_267) );
CKINVDCx16_ASAP7_75t_R g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g346 ( .A(n_252), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_252), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g294 ( .A(n_253), .B(n_284), .Y(n_294) );
AND2x2_ASAP7_75t_L g388 ( .A(n_253), .B(n_258), .Y(n_388) );
INVx1_ASAP7_75t_L g413 ( .A(n_253), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_259), .B1(n_262), .B2(n_263), .C(n_269), .Y(n_254) );
CKINVDCx14_ASAP7_75t_R g275 ( .A(n_255), .Y(n_275) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_256), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_259), .B(n_310), .Y(n_329) );
INVx3_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g378 ( .A(n_260), .B(n_274), .Y(n_378) );
AND2x2_ASAP7_75t_L g292 ( .A(n_261), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g322 ( .A(n_261), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_261), .B(n_305), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g392 ( .A(n_261), .B(n_362), .C(n_393), .Y(n_392) );
AOI211xp5_ASAP7_75t_SL g325 ( .A1(n_262), .A2(n_326), .B(n_328), .C(n_336), .Y(n_325) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OAI22xp33_ASAP7_75t_L g314 ( .A1(n_264), .A2(n_315), .B1(n_316), .B2(n_317), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_265), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_265), .B(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g407 ( .A(n_267), .B(n_381), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_275), .B1(n_276), .B2(n_278), .Y(n_269) );
NOR2xp33_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_273), .B(n_322), .Y(n_353) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_276), .A2(n_368), .B1(n_399), .B2(n_406), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_287), .B1(n_289), .B2(n_294), .C(n_295), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI221xp5_ASAP7_75t_L g295 ( .A1(n_285), .A2(n_296), .B1(n_302), .B2(n_303), .C(n_306), .Y(n_295) );
INVx1_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_SL g310 ( .A(n_291), .Y(n_310) );
OR2x2_ASAP7_75t_L g383 ( .A(n_291), .B(n_315), .Y(n_383) );
AND2x2_ASAP7_75t_L g385 ( .A(n_291), .B(n_293), .Y(n_385) );
INVx1_ASAP7_75t_L g324 ( .A(n_294), .Y(n_324) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
AOI21xp33_ASAP7_75t_SL g354 ( .A1(n_297), .A2(n_355), .B(n_356), .Y(n_354) );
OR2x2_ASAP7_75t_L g361 ( .A(n_297), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g335 ( .A(n_298), .B(n_319), .Y(n_335) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp33_ASAP7_75t_SL g352 ( .A(n_303), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_304), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_305), .B(n_341), .Y(n_404) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_308), .A2(n_321), .B(n_323), .C(n_324), .Y(n_320) );
NAND2x1_ASAP7_75t_SL g345 ( .A(n_308), .B(n_346), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_309), .A2(n_358), .B1(n_360), .B2(n_363), .Y(n_357) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_311), .B(n_401), .Y(n_400) );
NAND5xp2_ASAP7_75t_L g312 ( .A(n_313), .B(n_325), .C(n_343), .D(n_357), .E(n_366), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_320), .Y(n_313) );
INVx1_ASAP7_75t_L g370 ( .A(n_316), .Y(n_370) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_318), .A2(n_337), .B1(n_377), .B2(n_379), .C(n_382), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_319), .B(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_322), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_322), .B(n_388), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B1(n_332), .B2(n_334), .Y(n_328) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_340), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AND2x2_ASAP7_75t_L g410 ( .A(n_339), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B1(n_351), .B2(n_352), .C(n_354), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g394 ( .A(n_349), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g401 ( .A(n_359), .Y(n_401) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_369), .B(n_370), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI211xp5_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_374), .B(n_376), .C(n_389), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_374), .A2(n_399), .B(n_400), .C(n_402), .Y(n_398) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_378), .B(n_380), .Y(n_379) );
AOI21xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_386), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .B(n_414), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
NOR2x2_ASAP7_75t_L g694 ( .A(n_419), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_420), .Y(n_695) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
XOR2xp5_ASAP7_75t_L g707 ( .A(n_424), .B(n_708), .Y(n_707) );
OR3x1_ASAP7_75t_L g424 ( .A(n_425), .B(n_598), .C(n_645), .Y(n_424) );
NAND3xp33_ASAP7_75t_SL g425 ( .A(n_426), .B(n_544), .C(n_569), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_484), .B1(n_511), .B2(n_514), .C(n_522), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_452), .B(n_477), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_429), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_429), .B(n_527), .Y(n_642) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_443), .Y(n_429) );
AND2x2_ASAP7_75t_L g513 ( .A(n_430), .B(n_483), .Y(n_513) );
AND2x2_ASAP7_75t_L g562 ( .A(n_430), .B(n_482), .Y(n_562) );
AND2x2_ASAP7_75t_L g583 ( .A(n_430), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g588 ( .A(n_430), .B(n_555), .Y(n_588) );
OR2x2_ASAP7_75t_L g596 ( .A(n_430), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g668 ( .A(n_430), .B(n_465), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_430), .B(n_617), .Y(n_682) );
INVx3_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g528 ( .A(n_431), .B(n_443), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_431), .B(n_465), .Y(n_529) );
AND2x4_ASAP7_75t_L g550 ( .A(n_431), .B(n_483), .Y(n_550) );
AND2x2_ASAP7_75t_L g580 ( .A(n_431), .B(n_454), .Y(n_580) );
AND2x2_ASAP7_75t_L g589 ( .A(n_431), .B(n_579), .Y(n_589) );
AND2x2_ASAP7_75t_L g605 ( .A(n_431), .B(n_466), .Y(n_605) );
OR2x2_ASAP7_75t_L g614 ( .A(n_431), .B(n_597), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_431), .B(n_555), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_431), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g634 ( .A(n_431), .B(n_479), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_431), .B(n_524), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_431), .B(n_584), .Y(n_673) );
OR2x6_ASAP7_75t_L g431 ( .A(n_432), .B(n_441), .Y(n_431) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_439), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g483 ( .A(n_443), .Y(n_483) );
AND2x2_ASAP7_75t_L g579 ( .A(n_443), .B(n_465), .Y(n_579) );
AND2x2_ASAP7_75t_L g584 ( .A(n_443), .B(n_466), .Y(n_584) );
INVx1_ASAP7_75t_L g640 ( .A(n_443), .Y(n_640) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B(n_451), .Y(n_443) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_444), .A2(n_496), .B(n_502), .Y(n_495) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_444), .A2(n_504), .B(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g549 ( .A(n_453), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_465), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_454), .B(n_513), .Y(n_512) );
BUFx3_ASAP7_75t_L g527 ( .A(n_454), .Y(n_527) );
OR2x2_ASAP7_75t_L g597 ( .A(n_454), .B(n_465), .Y(n_597) );
OR2x2_ASAP7_75t_L g658 ( .A(n_454), .B(n_565), .Y(n_658) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_463), .Y(n_454) );
INVx1_ASAP7_75t_L g480 ( .A(n_456), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_463), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_465), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g617 ( .A(n_465), .B(n_479), .Y(n_617) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g556 ( .A(n_466), .Y(n_556) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_478), .A2(n_662), .B1(n_666), .B2(n_669), .C(n_670), .Y(n_661) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_482), .Y(n_478) );
INVx1_ASAP7_75t_SL g525 ( .A(n_479), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_479), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g656 ( .A(n_479), .B(n_513), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_482), .B(n_527), .Y(n_648) );
AND2x2_ASAP7_75t_L g555 ( .A(n_483), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_SL g559 ( .A(n_484), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_484), .B(n_565), .Y(n_595) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
AND2x2_ASAP7_75t_L g521 ( .A(n_485), .B(n_495), .Y(n_521) );
INVx4_ASAP7_75t_L g533 ( .A(n_485), .Y(n_533) );
BUFx3_ASAP7_75t_L g575 ( .A(n_485), .Y(n_575) );
AND3x2_ASAP7_75t_L g590 ( .A(n_485), .B(n_591), .C(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g672 ( .A(n_494), .B(n_586), .Y(n_672) );
AND2x2_ASAP7_75t_L g680 ( .A(n_494), .B(n_565), .Y(n_680) );
INVx1_ASAP7_75t_SL g685 ( .A(n_494), .Y(n_685) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_503), .Y(n_494) );
INVx1_ASAP7_75t_SL g543 ( .A(n_495), .Y(n_543) );
AND2x2_ASAP7_75t_L g566 ( .A(n_495), .B(n_533), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_495), .B(n_517), .Y(n_568) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_495), .Y(n_608) );
OR2x2_ASAP7_75t_L g613 ( .A(n_495), .B(n_533), .Y(n_613) );
INVx2_ASAP7_75t_L g519 ( .A(n_503), .Y(n_519) );
AND2x2_ASAP7_75t_L g553 ( .A(n_503), .B(n_534), .Y(n_553) );
OR2x2_ASAP7_75t_L g573 ( .A(n_503), .B(n_534), .Y(n_573) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_503), .Y(n_593) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_512), .A2(n_552), .B(n_644), .Y(n_643) );
AOI322xp5_ASAP7_75t_L g679 ( .A1(n_514), .A2(n_524), .A3(n_550), .B1(n_680), .B2(n_681), .C1(n_683), .C2(n_686), .Y(n_679) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_520), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_516), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_517), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g542 ( .A(n_518), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g610 ( .A(n_519), .B(n_533), .Y(n_610) );
AND2x2_ASAP7_75t_L g677 ( .A(n_519), .B(n_534), .Y(n_677) );
INVx1_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g618 ( .A(n_521), .B(n_572), .Y(n_618) );
AOI31xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_526), .A3(n_529), .B(n_530), .Y(n_522) );
AND2x2_ASAP7_75t_L g577 ( .A(n_524), .B(n_555), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_524), .B(n_547), .Y(n_659) );
AND2x2_ASAP7_75t_L g678 ( .A(n_524), .B(n_583), .Y(n_678) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_527), .B(n_555), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_527), .B(n_584), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_527), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_527), .B(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_528), .B(n_584), .Y(n_616) );
INVx1_ASAP7_75t_L g660 ( .A(n_528), .Y(n_660) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_542), .Y(n_531) );
INVxp67_ASAP7_75t_L g612 ( .A(n_532), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_533), .B(n_543), .Y(n_548) );
INVx1_ASAP7_75t_L g654 ( .A(n_533), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_533), .B(n_631), .Y(n_665) );
BUFx3_ASAP7_75t_L g565 ( .A(n_534), .Y(n_565) );
AND2x2_ASAP7_75t_L g591 ( .A(n_534), .B(n_543), .Y(n_591) );
INVx2_ASAP7_75t_L g631 ( .A(n_534), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_542), .B(n_664), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_549), .B(n_551), .C(n_560), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_546), .A2(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_547), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_547), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g627 ( .A(n_548), .B(n_573), .Y(n_627) );
INVx3_ASAP7_75t_L g558 ( .A(n_550), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_554), .B1(n_557), .B2(n_559), .Y(n_551) );
OAI21xp5_ASAP7_75t_SL g576 ( .A1(n_553), .A2(n_577), .B(n_578), .Y(n_576) );
AND2x2_ASAP7_75t_L g602 ( .A(n_553), .B(n_566), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_553), .B(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g557 ( .A(n_556), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g626 ( .A(n_556), .Y(n_626) );
OAI21xp5_ASAP7_75t_SL g570 ( .A1(n_557), .A2(n_571), .B(n_576), .Y(n_570) );
OAI22xp33_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_563), .B1(n_567), .B2(n_568), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_562), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g586 ( .A(n_565), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_565), .B(n_608), .Y(n_607) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_581), .C(n_594), .Y(n_569) );
OAI22xp5_ASAP7_75t_SL g636 ( .A1(n_571), .A2(n_637), .B1(n_641), .B2(n_642), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g641 ( .A(n_573), .B(n_574), .Y(n_641) );
AND2x2_ASAP7_75t_L g649 ( .A(n_574), .B(n_630), .Y(n_649) );
CKINVDCx16_ASAP7_75t_R g574 ( .A(n_575), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_SL g657 ( .A1(n_575), .A2(n_658), .B(n_659), .C(n_660), .Y(n_657) );
OR2x2_ASAP7_75t_L g684 ( .A(n_575), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B(n_587), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_583), .A2(n_620), .B(n_621), .C(n_624), .Y(n_619) );
OAI21xp33_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_589), .B(n_590), .Y(n_587) );
AND2x2_ASAP7_75t_L g652 ( .A(n_591), .B(n_610), .Y(n_652) );
INVxp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g630 ( .A(n_593), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g635 ( .A(n_595), .Y(n_635) );
NAND3xp33_ASAP7_75t_SL g598 ( .A(n_599), .B(n_619), .C(n_632), .Y(n_598) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B(n_603), .C(n_611), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g669 ( .A(n_606), .Y(n_669) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g629 ( .A(n_608), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_608), .B(n_677), .Y(n_676) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_614), .C(n_615), .Y(n_611) );
INVx2_ASAP7_75t_SL g623 ( .A(n_613), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_614), .A2(n_625), .B1(n_627), .B2(n_628), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_617), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_636), .C(n_643), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVxp33_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g686 ( .A(n_640), .Y(n_686) );
NAND4xp25_ASAP7_75t_L g645 ( .A(n_646), .B(n_661), .C(n_674), .D(n_679), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B(n_650), .C(n_657), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B(n_655), .Y(n_650) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_651), .A2(n_671), .B(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_658), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_678), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
NAND2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_702), .Y(n_697) );
NOR2xp33_ASAP7_75t_SL g698 ( .A(n_699), .B(n_701), .Y(n_698) );
INVx1_ASAP7_75t_SL g720 ( .A(n_699), .Y(n_720) );
INVx1_ASAP7_75t_L g719 ( .A(n_701), .Y(n_719) );
OA21x2_ASAP7_75t_L g722 ( .A1(n_701), .A2(n_720), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_704), .Y(n_711) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_704), .Y(n_713) );
BUFx2_ASAP7_75t_L g723 ( .A(n_704), .Y(n_723) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_711), .B(n_712), .Y(n_706) );
NOR2xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_714), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_716), .Y(n_715) );
CKINVDCx6p67_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
endmodule