module fake_jpeg_31559_n_58 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

INVx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx24_ASAP7_75t_SL g37 ( 
.A(n_33),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_26),
.C(n_24),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_41),
.C(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_39),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_20),
.B(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_46),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_24),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_36),
.C(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_9),
.C(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_45),
.Y(n_55)
);

NOR5xp2_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.C(n_53),
.D(n_51),
.E(n_54),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_43),
.B1(n_49),
.B2(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_56),
.Y(n_58)
);


endmodule