module real_aes_7595_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g459 ( .A1(n_0), .A2(n_160), .B(n_460), .C(n_463), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_1), .B(n_454), .Y(n_465) );
INVx1_ASAP7_75t_L g423 ( .A(n_2), .Y(n_423) );
INVx1_ASAP7_75t_L g209 ( .A(n_3), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_4), .B(n_148), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_5), .A2(n_438), .B(n_508), .Y(n_507) );
AOI222xp33_ASAP7_75t_L g99 ( .A1(n_6), .A2(n_100), .B1(n_727), .B2(n_736), .C1(n_749), .C2(n_755), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_6), .A2(n_9), .B1(n_418), .B2(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_6), .Y(n_745) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_7), .A2(n_165), .B(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_8), .A2(n_37), .B1(n_121), .B2(n_133), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_9), .A2(n_105), .B1(n_106), .B2(n_418), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_9), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_10), .B(n_165), .Y(n_198) );
AND2x6_ASAP7_75t_L g136 ( .A(n_11), .B(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_12), .A2(n_136), .B(n_441), .C(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_13), .B(n_38), .Y(n_424) );
INVx1_ASAP7_75t_L g117 ( .A(n_14), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_15), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g203 ( .A(n_16), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_17), .B(n_148), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_18), .B(n_163), .Y(n_181) );
AO32x2_ASAP7_75t_L g157 ( .A1(n_19), .A2(n_158), .A3(n_162), .B1(n_164), .B2(n_165), .Y(n_157) );
AOI222xp33_ASAP7_75t_SL g101 ( .A1(n_20), .A2(n_91), .B1(n_102), .B2(n_720), .C1(n_721), .C2(n_723), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_20), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_21), .B(n_121), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_22), .B(n_163), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_23), .A2(n_53), .B1(n_121), .B2(n_133), .Y(n_161) );
AOI22xp33_ASAP7_75t_SL g174 ( .A1(n_24), .A2(n_78), .B1(n_121), .B2(n_125), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_25), .B(n_121), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_26), .A2(n_164), .B(n_441), .C(n_443), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_27), .A2(n_164), .B(n_441), .C(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_28), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_29), .B(n_113), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_30), .A2(n_438), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_31), .B(n_113), .Y(n_155) );
INVx2_ASAP7_75t_L g123 ( .A(n_32), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_33), .A2(n_472), .B(n_473), .C(n_477), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_34), .B(n_121), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_35), .B(n_113), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_36), .B(n_128), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_39), .B(n_437), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_40), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_41), .B(n_148), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_42), .B(n_438), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_43), .A2(n_472), .B(n_477), .C(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_44), .Y(n_748) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_45), .B(n_121), .Y(n_191) );
INVx1_ASAP7_75t_L g461 ( .A(n_46), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_47), .A2(n_86), .B1(n_133), .B2(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g500 ( .A(n_48), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_49), .B(n_121), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_50), .B(n_121), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_51), .B(n_438), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_52), .B(n_196), .Y(n_195) );
AOI22xp33_ASAP7_75t_SL g185 ( .A1(n_54), .A2(n_58), .B1(n_121), .B2(n_125), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_55), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_56), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_57), .B(n_121), .Y(n_222) );
INVx1_ASAP7_75t_L g137 ( .A(n_59), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_60), .B(n_438), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_61), .B(n_454), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_62), .A2(n_196), .B(n_206), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_63), .B(n_121), .Y(n_210) );
INVx1_ASAP7_75t_L g116 ( .A(n_64), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_65), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_66), .B(n_148), .Y(n_475) );
AO32x2_ASAP7_75t_L g170 ( .A1(n_67), .A2(n_164), .A3(n_165), .B1(n_171), .B2(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_68), .B(n_149), .Y(n_531) );
INVx1_ASAP7_75t_L g221 ( .A(n_69), .Y(n_221) );
INVx1_ASAP7_75t_L g146 ( .A(n_70), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_71), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_72), .B(n_445), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_73), .A2(n_441), .B(n_477), .C(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_74), .B(n_125), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_75), .Y(n_509) );
INVx1_ASAP7_75t_L g731 ( .A(n_76), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_77), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_79), .B(n_133), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_80), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_81), .B(n_125), .Y(n_152) );
INVx2_ASAP7_75t_L g114 ( .A(n_82), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_83), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_84), .B(n_135), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_85), .B(n_125), .Y(n_192) );
OR2x2_ASAP7_75t_L g421 ( .A(n_87), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g719 ( .A(n_87), .Y(n_719) );
OR2x2_ASAP7_75t_L g735 ( .A(n_87), .B(n_726), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_88), .A2(n_98), .B1(n_125), .B2(n_126), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_89), .B(n_438), .Y(n_470) );
INVx1_ASAP7_75t_L g474 ( .A(n_90), .Y(n_474) );
INVxp67_ASAP7_75t_L g512 ( .A(n_92), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_93), .B(n_125), .Y(n_219) );
INVx1_ASAP7_75t_L g487 ( .A(n_94), .Y(n_487) );
INVx1_ASAP7_75t_L g527 ( .A(n_95), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_96), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g502 ( .A(n_97), .B(n_113), .Y(n_502) );
INVxp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22x1_ASAP7_75t_SL g102 ( .A1(n_103), .A2(n_419), .B1(n_425), .B2(n_716), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g721 ( .A1(n_104), .A2(n_426), .B1(n_716), .B2(n_722), .Y(n_721) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_105), .A2(n_106), .B1(n_743), .B2(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_340), .Y(n_106) );
NAND5xp2_ASAP7_75t_L g107 ( .A(n_108), .B(n_259), .C(n_274), .D(n_300), .E(n_322), .Y(n_107) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_239), .Y(n_108) );
OAI221xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_176), .B1(n_212), .B2(n_228), .C(n_229), .Y(n_109) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_166), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_111), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_SL g416 ( .A(n_111), .Y(n_416) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_139), .Y(n_111) );
INVx1_ASAP7_75t_L g256 ( .A(n_112), .Y(n_256) );
AND2x2_ASAP7_75t_L g258 ( .A(n_112), .B(n_157), .Y(n_258) );
AND2x2_ASAP7_75t_L g268 ( .A(n_112), .B(n_156), .Y(n_268) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_112), .Y(n_286) );
INVx1_ASAP7_75t_L g296 ( .A(n_112), .Y(n_296) );
OR2x2_ASAP7_75t_L g334 ( .A(n_112), .B(n_233), .Y(n_334) );
INVx2_ASAP7_75t_L g384 ( .A(n_112), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_112), .B(n_232), .Y(n_401) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B(n_138), .Y(n_112) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_113), .A2(n_143), .B(n_155), .Y(n_142) );
INVx2_ASAP7_75t_L g175 ( .A(n_113), .Y(n_175) );
INVx1_ASAP7_75t_L g451 ( .A(n_113), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_113), .A2(n_470), .B(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_113), .A2(n_497), .B(n_498), .Y(n_496) );
AND2x2_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x2_ASAP7_75t_L g163 ( .A(n_114), .B(n_115), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_130), .B(n_136), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B(n_127), .Y(n_119) );
INVx3_ASAP7_75t_L g145 ( .A(n_121), .Y(n_145) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_121), .Y(n_489) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g133 ( .A(n_122), .Y(n_133) );
BUFx3_ASAP7_75t_L g173 ( .A(n_122), .Y(n_173) );
AND2x6_ASAP7_75t_L g441 ( .A(n_122), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g126 ( .A(n_123), .Y(n_126) );
INVx1_ASAP7_75t_L g197 ( .A(n_123), .Y(n_197) );
INVx2_ASAP7_75t_L g204 ( .A(n_125), .Y(n_204) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_129), .Y(n_135) );
INVx3_ASAP7_75t_L g149 ( .A(n_129), .Y(n_149) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_129), .Y(n_154) );
AND2x2_ASAP7_75t_L g439 ( .A(n_129), .B(n_197), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_129), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B(n_134), .Y(n_130) );
O2A1O1Ixp5_ASAP7_75t_L g220 ( .A1(n_134), .A2(n_208), .B(n_221), .C(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g158 ( .A1(n_135), .A2(n_159), .B1(n_160), .B2(n_161), .Y(n_158) );
OAI22xp5_ASAP7_75t_SL g171 ( .A1(n_135), .A2(n_149), .B1(n_172), .B2(n_174), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_135), .A2(n_160), .B1(n_184), .B2(n_185), .Y(n_183) );
INVx4_ASAP7_75t_L g462 ( .A(n_135), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_136), .A2(n_144), .B(n_150), .Y(n_143) );
BUFx3_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_136), .A2(n_190), .B(n_193), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_136), .A2(n_202), .B(n_207), .Y(n_201) );
AND2x4_ASAP7_75t_L g438 ( .A(n_136), .B(n_439), .Y(n_438) );
INVx4_ASAP7_75t_SL g464 ( .A(n_136), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_136), .B(n_439), .Y(n_528) );
NOR2xp67_ASAP7_75t_L g139 ( .A(n_140), .B(n_156), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_141), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_141), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_SL g316 ( .A(n_141), .B(n_256), .Y(n_316) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
INVx2_ASAP7_75t_L g233 ( .A(n_142), .Y(n_233) );
OR2x2_ASAP7_75t_L g295 ( .A(n_142), .B(n_296), .Y(n_295) );
O2A1O1Ixp5_ASAP7_75t_SL g144 ( .A1(n_145), .A2(n_146), .B(n_147), .C(n_148), .Y(n_144) );
INVx2_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_148), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_148), .A2(n_218), .B(n_219), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_148), .B(n_512), .Y(n_511) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g206 ( .A(n_153), .Y(n_206) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g445 ( .A(n_154), .Y(n_445) );
AND2x2_ASAP7_75t_L g234 ( .A(n_156), .B(n_170), .Y(n_234) );
AND2x2_ASAP7_75t_L g251 ( .A(n_156), .B(n_231), .Y(n_251) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g169 ( .A(n_157), .B(n_170), .Y(n_169) );
BUFx2_ASAP7_75t_L g254 ( .A(n_157), .Y(n_254) );
AND2x2_ASAP7_75t_L g383 ( .A(n_157), .B(n_384), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_160), .A2(n_194), .B(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_160), .A2(n_208), .B(n_209), .C(n_210), .Y(n_207) );
INVx2_ASAP7_75t_L g200 ( .A(n_162), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_162), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_163), .Y(n_165) );
NAND3xp33_ASAP7_75t_L g182 ( .A(n_164), .B(n_183), .C(n_186), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_164), .A2(n_217), .B(n_220), .Y(n_216) );
INVx4_ASAP7_75t_L g186 ( .A(n_165), .Y(n_186) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_165), .A2(n_189), .B(n_198), .Y(n_188) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_165), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_165), .A2(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g228 ( .A(n_166), .Y(n_228) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_169), .Y(n_166) );
AND2x2_ASAP7_75t_L g346 ( .A(n_167), .B(n_234), .Y(n_346) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g347 ( .A(n_168), .B(n_258), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_169), .A2(n_315), .B(n_317), .C(n_319), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_169), .B(n_315), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_169), .A2(n_245), .B1(n_388), .B2(n_389), .C(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g231 ( .A(n_170), .Y(n_231) );
INVx1_ASAP7_75t_L g267 ( .A(n_170), .Y(n_267) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_170), .Y(n_276) );
INVx2_ASAP7_75t_L g463 ( .A(n_173), .Y(n_463) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_173), .Y(n_476) );
INVx1_ASAP7_75t_L g448 ( .A(n_175), .Y(n_448) );
INVx1_ASAP7_75t_SL g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_187), .Y(n_177) );
AND2x2_ASAP7_75t_L g293 ( .A(n_178), .B(n_238), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_178), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_179), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g385 ( .A(n_179), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g417 ( .A(n_179), .Y(n_417) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx3_ASAP7_75t_L g247 ( .A(n_180), .Y(n_247) );
AND2x2_ASAP7_75t_L g273 ( .A(n_180), .B(n_227), .Y(n_273) );
NOR2x1_ASAP7_75t_L g282 ( .A(n_180), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g289 ( .A(n_180), .B(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g225 ( .A(n_181), .Y(n_225) );
AO21x1_ASAP7_75t_L g224 ( .A1(n_183), .A2(n_186), .B(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g454 ( .A(n_186), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_186), .B(n_479), .Y(n_478) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_186), .A2(n_484), .B(n_491), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_186), .B(n_492), .Y(n_491) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_186), .A2(n_526), .B(n_533), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_187), .B(n_329), .Y(n_364) );
INVx1_ASAP7_75t_SL g368 ( .A(n_187), .Y(n_368) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_199), .Y(n_187) );
INVx3_ASAP7_75t_L g227 ( .A(n_188), .Y(n_227) );
AND2x2_ASAP7_75t_L g238 ( .A(n_188), .B(n_215), .Y(n_238) );
AND2x2_ASAP7_75t_L g260 ( .A(n_188), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g305 ( .A(n_188), .B(n_299), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_188), .B(n_237), .Y(n_386) );
INVx2_ASAP7_75t_L g208 ( .A(n_196), .Y(n_208) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g226 ( .A(n_199), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g237 ( .A(n_199), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_199), .B(n_215), .Y(n_262) );
AND2x2_ASAP7_75t_L g298 ( .A(n_199), .B(n_299), .Y(n_298) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_211), .Y(n_199) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_200), .A2(n_216), .B(n_223), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .C(n_206), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_204), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_204), .A2(n_531), .B(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_206), .A2(n_487), .B(n_488), .C(n_489), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_208), .A2(n_444), .B(n_446), .Y(n_443) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_226), .Y(n_213) );
INVx1_ASAP7_75t_L g278 ( .A(n_214), .Y(n_278) );
AND2x2_ASAP7_75t_L g320 ( .A(n_214), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_214), .B(n_241), .Y(n_326) );
AOI21xp5_ASAP7_75t_SL g400 ( .A1(n_214), .A2(n_232), .B(n_255), .Y(n_400) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_224), .Y(n_214) );
OR2x2_ASAP7_75t_L g243 ( .A(n_215), .B(n_224), .Y(n_243) );
AND2x2_ASAP7_75t_L g290 ( .A(n_215), .B(n_227), .Y(n_290) );
INVx2_ASAP7_75t_L g299 ( .A(n_215), .Y(n_299) );
INVx1_ASAP7_75t_L g405 ( .A(n_215), .Y(n_405) );
AND2x2_ASAP7_75t_L g329 ( .A(n_224), .B(n_299), .Y(n_329) );
INVx1_ASAP7_75t_L g354 ( .A(n_224), .Y(n_354) );
AND2x2_ASAP7_75t_L g263 ( .A(n_226), .B(n_247), .Y(n_263) );
AND2x2_ASAP7_75t_L g275 ( .A(n_226), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_SL g393 ( .A(n_226), .Y(n_393) );
INVx2_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
AND2x2_ASAP7_75t_L g321 ( .A(n_227), .B(n_237), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_227), .B(n_405), .Y(n_404) );
OAI21xp33_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_234), .B(n_235), .Y(n_229) );
AND2x2_ASAP7_75t_L g336 ( .A(n_230), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g390 ( .A(n_230), .Y(n_390) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g310 ( .A(n_231), .Y(n_310) );
BUFx2_ASAP7_75t_L g409 ( .A(n_231), .Y(n_409) );
BUFx2_ASAP7_75t_L g280 ( .A(n_232), .Y(n_280) );
AND2x2_ASAP7_75t_L g382 ( .A(n_232), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g365 ( .A(n_233), .Y(n_365) );
AND2x4_ASAP7_75t_L g292 ( .A(n_234), .B(n_255), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_234), .B(n_316), .Y(n_328) );
AOI32xp33_ASAP7_75t_L g252 ( .A1(n_235), .A2(n_253), .A3(n_255), .B1(n_257), .B2(n_258), .Y(n_252) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
INVx3_ASAP7_75t_L g241 ( .A(n_236), .Y(n_241) );
OR2x2_ASAP7_75t_L g377 ( .A(n_236), .B(n_333), .Y(n_377) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g246 ( .A(n_237), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g353 ( .A(n_237), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g245 ( .A(n_238), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g257 ( .A(n_238), .B(n_247), .Y(n_257) );
INVx1_ASAP7_75t_L g378 ( .A(n_238), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_238), .B(n_353), .Y(n_411) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_244), .B(n_248), .C(n_252), .Y(n_239) );
OAI322xp33_ASAP7_75t_L g348 ( .A1(n_240), .A2(n_285), .A3(n_349), .B1(n_351), .B2(n_355), .C1(n_356), .C2(n_360), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVxp67_ASAP7_75t_L g313 ( .A(n_241), .Y(n_313) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g367 ( .A(n_243), .B(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_243), .B(n_283), .Y(n_414) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g306 ( .A(n_246), .Y(n_306) );
OR2x2_ASAP7_75t_L g392 ( .A(n_247), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_250), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g301 ( .A(n_251), .B(n_280), .Y(n_301) );
AND2x2_ASAP7_75t_L g372 ( .A(n_251), .B(n_285), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_251), .B(n_359), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g259 ( .A1(n_253), .A2(n_260), .B1(n_263), .B2(n_264), .C(n_269), .Y(n_259) );
OR2x2_ASAP7_75t_L g270 ( .A(n_253), .B(n_266), .Y(n_270) );
AND2x2_ASAP7_75t_L g358 ( .A(n_253), .B(n_359), .Y(n_358) );
AOI32xp33_ASAP7_75t_L g397 ( .A1(n_253), .A2(n_283), .A3(n_398), .B1(n_399), .B2(n_402), .Y(n_397) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_254), .B(n_290), .C(n_313), .Y(n_331) );
AND2x2_ASAP7_75t_L g357 ( .A(n_254), .B(n_350), .Y(n_357) );
INVxp67_ASAP7_75t_L g337 ( .A(n_255), .Y(n_337) );
BUFx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_258), .B(n_310), .Y(n_366) );
INVx2_ASAP7_75t_L g376 ( .A(n_258), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_258), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g345 ( .A(n_261), .Y(n_345) );
OR2x2_ASAP7_75t_L g271 ( .A(n_262), .B(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_264), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_267), .Y(n_350) );
AND2x2_ASAP7_75t_L g309 ( .A(n_268), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g355 ( .A(n_268), .Y(n_355) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_268), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AOI21xp33_ASAP7_75t_SL g294 ( .A1(n_270), .A2(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g388 ( .A(n_273), .B(n_298), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_277), .B(n_287), .C(n_294), .Y(n_274) );
AND2x2_ASAP7_75t_L g318 ( .A(n_276), .B(n_286), .Y(n_318) );
INVx2_ASAP7_75t_L g333 ( .A(n_276), .Y(n_333) );
OR2x2_ASAP7_75t_L g371 ( .A(n_276), .B(n_334), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_276), .B(n_414), .Y(n_413) );
AOI211xp5_ASAP7_75t_SL g277 ( .A1(n_278), .A2(n_279), .B(n_281), .C(n_284), .Y(n_277) );
INVxp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_280), .B(n_318), .Y(n_317) );
OAI211xp5_ASAP7_75t_L g399 ( .A1(n_281), .A2(n_376), .B(n_400), .C(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2x1p5_ASAP7_75t_L g297 ( .A(n_282), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g339 ( .A(n_283), .B(n_329), .Y(n_339) );
INVx1_ASAP7_75t_L g344 ( .A(n_283), .Y(n_344) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVxp33_ASAP7_75t_L g395 ( .A(n_289), .Y(n_395) );
AND2x2_ASAP7_75t_L g374 ( .A(n_290), .B(n_353), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_295), .A2(n_357), .B(n_358), .Y(n_356) );
OAI322xp33_ASAP7_75t_L g375 ( .A1(n_297), .A2(n_376), .A3(n_377), .B1(n_378), .B2(n_379), .C1(n_381), .C2(n_385), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B1(n_307), .B2(n_311), .C(n_314), .Y(n_300) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g352 ( .A(n_305), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g396 ( .A(n_309), .Y(n_396) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_312), .B(n_332), .Y(n_398) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g361 ( .A(n_321), .B(n_329), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_325), .B1(n_327), .B2(n_329), .C(n_330), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_325), .A2(n_342), .B1(n_346), .B2(n_347), .C(n_348), .Y(n_341) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_329), .B(n_344), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B1(n_335), .B2(n_338), .Y(n_330) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx2_ASAP7_75t_SL g359 ( .A(n_334), .Y(n_359) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND5xp2_ASAP7_75t_L g340 ( .A(n_341), .B(n_362), .C(n_387), .D(n_397), .E(n_407), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_343), .B(n_345), .Y(n_342) );
NOR4xp25_ASAP7_75t_L g415 ( .A(n_344), .B(n_350), .C(n_416), .D(n_417), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_347), .A2(n_408), .B1(n_410), .B2(n_412), .C(n_415), .Y(n_407) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g406 ( .A(n_353), .Y(n_406) );
OAI322xp33_ASAP7_75t_L g363 ( .A1(n_357), .A2(n_364), .A3(n_365), .B1(n_366), .B2(n_367), .C1(n_369), .C2(n_373), .Y(n_363) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_375), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g408 ( .A(n_383), .B(n_409), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B1(n_395), .B2(n_396), .Y(n_391) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g722 ( .A(n_420), .Y(n_722) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g718 ( .A(n_422), .B(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g726 ( .A(n_422), .Y(n_726) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_SL g426 ( .A(n_427), .B(n_671), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_606), .Y(n_427) );
NAND4xp25_ASAP7_75t_SL g428 ( .A(n_429), .B(n_551), .C(n_575), .D(n_598), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_493), .B1(n_523), .B2(n_535), .C(n_538), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_466), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_432), .A2(n_452), .B1(n_494), .B2(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_432), .B(n_467), .Y(n_609) );
AND2x2_ASAP7_75t_L g628 ( .A(n_432), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_432), .B(n_612), .Y(n_698) );
AND2x4_ASAP7_75t_L g432 ( .A(n_433), .B(n_452), .Y(n_432) );
AND2x2_ASAP7_75t_L g566 ( .A(n_433), .B(n_467), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_433), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g589 ( .A(n_433), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g594 ( .A(n_433), .B(n_453), .Y(n_594) );
INVx2_ASAP7_75t_L g626 ( .A(n_433), .Y(n_626) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_433), .Y(n_670) );
AND2x2_ASAP7_75t_L g687 ( .A(n_433), .B(n_564), .Y(n_687) );
INVx5_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g605 ( .A(n_434), .B(n_564), .Y(n_605) );
AND2x4_ASAP7_75t_L g619 ( .A(n_434), .B(n_452), .Y(n_619) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_434), .Y(n_623) );
AND2x2_ASAP7_75t_L g643 ( .A(n_434), .B(n_558), .Y(n_643) );
AND2x2_ASAP7_75t_L g693 ( .A(n_434), .B(n_468), .Y(n_693) );
AND2x2_ASAP7_75t_L g703 ( .A(n_434), .B(n_453), .Y(n_703) );
OR2x6_ASAP7_75t_L g434 ( .A(n_435), .B(n_449), .Y(n_434) );
AOI21xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_440), .B(n_448), .Y(n_435) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx5_ASAP7_75t_L g458 ( .A(n_441), .Y(n_458) );
INVx2_ASAP7_75t_L g447 ( .A(n_445), .Y(n_447) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_447), .A2(n_474), .B(n_475), .C(n_476), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_447), .A2(n_476), .B(n_500), .C(n_501), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AND2x2_ASAP7_75t_L g559 ( .A(n_452), .B(n_467), .Y(n_559) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_452), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_452), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g649 ( .A(n_452), .Y(n_649) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g537 ( .A(n_453), .B(n_482), .Y(n_537) );
AND2x2_ASAP7_75t_L g564 ( .A(n_453), .B(n_483), .Y(n_564) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B(n_465), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_458), .B(n_459), .C(n_464), .Y(n_456) );
INVx2_ASAP7_75t_L g472 ( .A(n_458), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_458), .A2(n_464), .B(n_509), .C(n_510), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g477 ( .A(n_464), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_466), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_480), .Y(n_466) );
OR2x2_ASAP7_75t_L g590 ( .A(n_467), .B(n_481), .Y(n_590) );
AND2x2_ASAP7_75t_L g627 ( .A(n_467), .B(n_537), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_467), .B(n_558), .Y(n_638) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_467), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_467), .B(n_594), .Y(n_711) );
INVx5_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g536 ( .A(n_468), .Y(n_536) );
AND2x2_ASAP7_75t_L g545 ( .A(n_468), .B(n_481), .Y(n_545) );
AND2x2_ASAP7_75t_L g661 ( .A(n_468), .B(n_556), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_468), .B(n_594), .Y(n_683) );
OR2x6_ASAP7_75t_L g468 ( .A(n_469), .B(n_478), .Y(n_468) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_481), .Y(n_629) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_482), .Y(n_581) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g558 ( .A(n_483), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_490), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_494), .B(n_571), .Y(n_690) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_495), .B(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g542 ( .A(n_495), .B(n_543), .Y(n_542) );
INVx5_ASAP7_75t_SL g550 ( .A(n_495), .Y(n_550) );
OR2x2_ASAP7_75t_L g573 ( .A(n_495), .B(n_543), .Y(n_573) );
OR2x2_ASAP7_75t_L g583 ( .A(n_495), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g646 ( .A(n_495), .B(n_505), .Y(n_646) );
AND2x2_ASAP7_75t_SL g684 ( .A(n_495), .B(n_504), .Y(n_684) );
NOR4xp25_ASAP7_75t_L g705 ( .A(n_495), .B(n_626), .C(n_706), .D(n_707), .Y(n_705) );
AND2x2_ASAP7_75t_L g715 ( .A(n_495), .B(n_547), .Y(n_715) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g540 ( .A(n_504), .B(n_536), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_504), .B(n_542), .Y(n_709) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
OR2x2_ASAP7_75t_L g549 ( .A(n_505), .B(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g556 ( .A(n_505), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_505), .B(n_525), .Y(n_568) );
INVxp67_ASAP7_75t_L g571 ( .A(n_505), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_505), .B(n_543), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_505), .B(n_515), .Y(n_637) );
AND2x2_ASAP7_75t_L g652 ( .A(n_505), .B(n_547), .Y(n_652) );
OR2x2_ASAP7_75t_L g681 ( .A(n_505), .B(n_515), .Y(n_681) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_513), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_514), .B(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_514), .B(n_550), .Y(n_689) );
OR2x2_ASAP7_75t_L g710 ( .A(n_514), .B(n_587), .Y(n_710) );
INVx1_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g524 ( .A(n_515), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g547 ( .A(n_515), .B(n_543), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_515), .B(n_525), .Y(n_562) );
AND2x2_ASAP7_75t_L g632 ( .A(n_515), .B(n_556), .Y(n_632) );
AND2x2_ASAP7_75t_L g666 ( .A(n_515), .B(n_550), .Y(n_666) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_516), .B(n_550), .Y(n_569) );
AND2x2_ASAP7_75t_L g597 ( .A(n_516), .B(n_525), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_523), .B(n_605), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_524), .A2(n_612), .B1(n_648), .B2(n_665), .C(n_667), .Y(n_664) );
INVx5_ASAP7_75t_SL g543 ( .A(n_525), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_529), .Y(n_526) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
OAI33xp33_ASAP7_75t_L g563 ( .A1(n_536), .A2(n_564), .A3(n_565), .B1(n_567), .B2(n_570), .B3(n_574), .Y(n_563) );
OR2x2_ASAP7_75t_L g579 ( .A(n_536), .B(n_580), .Y(n_579) );
AOI322xp5_ASAP7_75t_L g688 ( .A1(n_536), .A2(n_605), .A3(n_612), .B1(n_689), .B2(n_690), .C1(n_691), .C2(n_694), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_536), .B(n_564), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_SL g712 ( .A1(n_536), .A2(n_564), .B(n_713), .C(n_715), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_537), .A2(n_552), .B1(n_557), .B2(n_560), .C(n_563), .Y(n_551) );
INVx1_ASAP7_75t_L g644 ( .A(n_537), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_537), .B(n_693), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_541), .B1(n_544), .B2(n_546), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g621 ( .A(n_542), .B(n_556), .Y(n_621) );
AND2x2_ASAP7_75t_L g679 ( .A(n_542), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g587 ( .A(n_543), .B(n_550), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_543), .B(n_556), .Y(n_615) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_545), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_545), .B(n_623), .Y(n_677) );
OAI321xp33_ASAP7_75t_L g696 ( .A1(n_545), .A2(n_618), .A3(n_697), .B1(n_698), .B2(n_699), .C(n_700), .Y(n_696) );
INVx1_ASAP7_75t_L g663 ( .A(n_546), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_547), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g602 ( .A(n_547), .B(n_550), .Y(n_602) );
AOI321xp33_ASAP7_75t_L g660 ( .A1(n_547), .A2(n_564), .A3(n_661), .B1(n_662), .B2(n_663), .C(n_664), .Y(n_660) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g577 ( .A(n_549), .B(n_562), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_550), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_550), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_550), .B(n_636), .Y(n_673) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g596 ( .A(n_554), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g561 ( .A(n_555), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g669 ( .A(n_556), .Y(n_669) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_559), .B(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g592 ( .A(n_564), .Y(n_592) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_566), .B(n_601), .Y(n_650) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OR2x2_ASAP7_75t_L g614 ( .A(n_569), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g659 ( .A(n_569), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_570), .A2(n_617), .B1(n_620), .B2(n_622), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g714 ( .A(n_573), .B(n_637), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_578), .B1(n_582), .B2(n_588), .C(n_591), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx2_ASAP7_75t_L g612 ( .A(n_581), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_SL g658 ( .A(n_584), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_586), .B(n_636), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_586), .A2(n_654), .B(n_656), .Y(n_653) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g699 ( .A(n_587), .B(n_681), .Y(n_699) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_SL g601 ( .A(n_590), .Y(n_601) );
AOI21xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g645 ( .A(n_597), .B(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_L g707 ( .A(n_597), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B(n_603), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_601), .B(n_619), .Y(n_655) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g676 ( .A(n_605), .Y(n_676) );
NAND5xp2_ASAP7_75t_L g606 ( .A(n_607), .B(n_624), .C(n_633), .D(n_653), .E(n_660), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B(n_613), .C(n_616), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g648 ( .A(n_612), .Y(n_648) );
CKINVDCx16_ASAP7_75t_R g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_620), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g662 ( .A(n_622), .Y(n_662) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_628), .B(n_630), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_625), .A2(n_679), .B1(n_682), .B2(n_684), .C(n_685), .Y(n_678) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AOI321xp33_ASAP7_75t_L g633 ( .A1(n_626), .A2(n_634), .A3(n_638), .B1(n_639), .B2(n_645), .C(n_647), .Y(n_633) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g704 ( .A(n_638), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_640), .B(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g656 ( .A(n_641), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NOR2xp67_ASAP7_75t_SL g668 ( .A(n_642), .B(n_649), .Y(n_668) );
AOI321xp33_ASAP7_75t_SL g700 ( .A1(n_645), .A2(n_701), .A3(n_702), .B1(n_703), .B2(n_704), .C(n_705), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B(n_650), .C(n_651), .Y(n_647) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_658), .B(n_666), .Y(n_695) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .C(n_670), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_696), .C(n_708), .Y(n_671) );
OAI211xp5_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_674), .B(n_678), .C(n_688), .Y(n_672) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_676), .B(n_677), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_677), .A2(n_709), .B1(n_710), .B2(n_711), .C(n_712), .Y(n_708) );
INVx1_ASAP7_75t_L g697 ( .A(n_679), .Y(n_697) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g701 ( .A(n_699), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
CKINVDCx14_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2x2_ASAP7_75t_L g725 ( .A(n_719), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
NAND2xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_733), .Y(n_728) );
NOR2xp33_ASAP7_75t_SL g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_SL g754 ( .A(n_730), .Y(n_754) );
INVx1_ASAP7_75t_L g753 ( .A(n_732), .Y(n_753) );
OA21x2_ASAP7_75t_L g756 ( .A1(n_732), .A2(n_754), .B(n_757), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_733), .A2(n_738), .B(n_746), .Y(n_737) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_735), .Y(n_747) );
BUFx2_ASAP7_75t_L g757 ( .A(n_735), .Y(n_757) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_SL g746 ( .A(n_747), .B(n_748), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
endmodule