module fake_aes_703_n_1251 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1251);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1251;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_634;
wire n_307;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_659;
wire n_432;
wire n_386;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_416;
wire n_536;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_755;
wire n_848;
wire n_1031;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g299 ( .A(n_269), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_126), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_35), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_192), .Y(n_302) );
CKINVDCx16_ASAP7_75t_R g303 ( .A(n_27), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_218), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_196), .Y(n_305) );
INVxp67_ASAP7_75t_L g306 ( .A(n_146), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_108), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_235), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_160), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_45), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_294), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_262), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_195), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_239), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_191), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_81), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_240), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_156), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_183), .Y(n_319) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_247), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_171), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_41), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_24), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
INVxp33_ASAP7_75t_SL g325 ( .A(n_104), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_54), .Y(n_326) );
INVxp33_ASAP7_75t_SL g327 ( .A(n_284), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_292), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_238), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_107), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_95), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_275), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_139), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_245), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_155), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_71), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_12), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_193), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_251), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_213), .Y(n_340) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_121), .Y(n_341) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_276), .Y(n_342) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_273), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_28), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_64), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_59), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_228), .Y(n_347) );
INVxp33_ASAP7_75t_L g348 ( .A(n_236), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_79), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_56), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_128), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_154), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_62), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g354 ( .A(n_177), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_200), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_34), .Y(n_356) );
CKINVDCx16_ASAP7_75t_R g357 ( .A(n_80), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_129), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_76), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_43), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_254), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_176), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_145), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_76), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_25), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_22), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_115), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_255), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_165), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_113), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_31), .Y(n_371) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_151), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_162), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_96), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_221), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_207), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_119), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_48), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_246), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_45), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_173), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_204), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_282), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_29), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_24), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_263), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_105), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_136), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_283), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_184), .Y(n_390) );
INVxp33_ASAP7_75t_L g391 ( .A(n_74), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_44), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_43), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_56), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_167), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_270), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_106), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_288), .Y(n_398) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_169), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_252), .Y(n_400) );
INVxp33_ASAP7_75t_SL g401 ( .A(n_64), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_194), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_172), .Y(n_403) );
INVxp33_ASAP7_75t_SL g404 ( .A(n_51), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_229), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_23), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_178), .Y(n_407) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_133), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_134), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_81), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_101), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_92), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_35), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_38), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_130), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_2), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_234), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_30), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_111), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_112), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_293), .Y(n_421) );
INVxp33_ASAP7_75t_SL g422 ( .A(n_250), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_265), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_65), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_222), .Y(n_425) );
INVxp33_ASAP7_75t_SL g426 ( .A(n_51), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_264), .Y(n_427) );
INVxp33_ASAP7_75t_SL g428 ( .A(n_122), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_206), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_37), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_86), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_59), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_268), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_42), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_4), .Y(n_435) );
INVxp33_ASAP7_75t_L g436 ( .A(n_187), .Y(n_436) );
INVxp33_ASAP7_75t_L g437 ( .A(n_253), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_55), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_7), .Y(n_439) );
BUFx10_ASAP7_75t_L g440 ( .A(n_164), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_158), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_257), .Y(n_442) );
INVxp33_ASAP7_75t_SL g443 ( .A(n_274), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_98), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_55), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_186), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_135), .Y(n_447) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_19), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_25), .Y(n_449) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_299), .A2(n_0), .B(n_1), .Y(n_450) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_299), .A2(n_0), .B(n_1), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_309), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_350), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_341), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_350), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_350), .B(n_2), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_342), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_354), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_302), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_347), .B(n_3), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_347), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_332), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_417), .B(n_3), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_302), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_417), .B(n_429), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_332), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_429), .B(n_4), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_303), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_333), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_310), .B(n_5), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_442), .B(n_5), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_313), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_309), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_310), .B(n_6), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_333), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_334), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_336), .B(n_6), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_334), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_309), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_309), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_335), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_313), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_335), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_391), .B(n_7), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_473), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_456), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_462), .B(n_305), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_473), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_456), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_456), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_473), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_473), .Y(n_492) );
AND2x4_ASAP7_75t_SL g493 ( .A(n_470), .B(n_339), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_456), .B(n_326), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_465), .B(n_348), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_473), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_450), .B(n_444), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_456), .Y(n_498) );
INVx3_ASAP7_75t_L g499 ( .A(n_450), .Y(n_499) );
OAI22xp5_ASAP7_75t_SL g500 ( .A1(n_468), .A2(n_344), .B1(n_418), .B2(n_393), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_450), .Y(n_501) );
INVx4_ASAP7_75t_L g502 ( .A(n_450), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_470), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_453), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_450), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_462), .B(n_446), .C(n_444), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_455), .Y(n_509) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_473), .Y(n_510) );
BUFx3_ASAP7_75t_L g511 ( .A(n_455), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_466), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_465), .B(n_440), .Y(n_513) );
BUFx10_ASAP7_75t_L g514 ( .A(n_461), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_450), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_473), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_470), .B(n_326), .Y(n_517) );
OAI221xp5_ASAP7_75t_L g518 ( .A1(n_477), .A2(n_448), .B1(n_345), .B2(n_336), .C(n_384), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_452), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_466), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_469), .B(n_305), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_451), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_474), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g524 ( .A(n_451), .B(n_446), .Y(n_524) );
CKINVDCx11_ASAP7_75t_R g525 ( .A(n_468), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_490), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_490), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_490), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_495), .B(n_461), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_490), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_499), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_504), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_511), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_495), .B(n_474), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_486), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_493), .Y(n_536) );
INVx4_ASAP7_75t_L g537 ( .A(n_494), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_503), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_511), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_504), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_525), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_506), .Y(n_542) );
OR2x6_ASAP7_75t_L g543 ( .A(n_517), .B(n_474), .Y(n_543) );
NOR3xp33_ASAP7_75t_SL g544 ( .A(n_518), .B(n_464), .C(n_459), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_486), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_525), .Y(n_546) );
OR2x4_ASAP7_75t_L g547 ( .A(n_489), .B(n_471), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_503), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_523), .B(n_460), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_489), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_523), .B(n_460), .Y(n_551) );
INVx8_ASAP7_75t_L g552 ( .A(n_517), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_499), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_517), .Y(n_554) );
AND3x2_ASAP7_75t_SL g555 ( .A(n_514), .B(n_378), .C(n_365), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_513), .B(n_463), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_513), .B(n_463), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_517), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_493), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_506), .Y(n_560) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_515), .A2(n_467), .B(n_477), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_499), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_499), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_499), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_513), .B(n_467), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_494), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_514), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_517), .B(n_469), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_498), .Y(n_569) );
BUFx8_ASAP7_75t_L g570 ( .A(n_494), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_512), .B(n_457), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_494), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_509), .Y(n_573) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_511), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_512), .B(n_475), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_509), .Y(n_576) );
NOR2x1p5_ASAP7_75t_L g577 ( .A(n_500), .B(n_457), .Y(n_577) );
INVx5_ASAP7_75t_L g578 ( .A(n_494), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_498), .B(n_471), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_501), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_511), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_514), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_512), .B(n_475), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_502), .Y(n_584) );
NAND2x1p5_ASAP7_75t_L g585 ( .A(n_502), .B(n_451), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_520), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_520), .B(n_454), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_520), .Y(n_588) );
OR2x6_ASAP7_75t_L g589 ( .A(n_497), .B(n_451), .Y(n_589) );
NOR3xp33_ASAP7_75t_SL g590 ( .A(n_518), .B(n_472), .C(n_482), .Y(n_590) );
INVx2_ASAP7_75t_SL g591 ( .A(n_514), .Y(n_591) );
NOR3xp33_ASAP7_75t_SL g592 ( .A(n_500), .B(n_482), .C(n_357), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_487), .B(n_476), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_487), .B(n_476), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_514), .B(n_458), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_493), .B(n_478), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_565), .B(n_493), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_537), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_565), .B(n_484), .Y(n_599) );
OAI21x1_ASAP7_75t_L g600 ( .A1(n_584), .A2(n_505), .B(n_501), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_556), .B(n_521), .Y(n_601) );
BUFx3_ASAP7_75t_L g602 ( .A(n_570), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_596), .A2(n_377), .B1(n_339), .B2(n_401), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_566), .Y(n_604) );
CKINVDCx8_ASAP7_75t_R g605 ( .A(n_541), .Y(n_605) );
INVx3_ASAP7_75t_L g606 ( .A(n_537), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_570), .Y(n_607) );
AOI222xp33_ASAP7_75t_L g608 ( .A1(n_549), .A2(n_432), .B1(n_344), .B2(n_438), .C1(n_418), .C2(n_393), .Y(n_608) );
BUFx3_ASAP7_75t_L g609 ( .A(n_570), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_557), .B(n_521), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_566), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_529), .B(n_401), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_588), .B(n_502), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_533), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_543), .B(n_502), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_543), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_549), .A2(n_377), .B1(n_426), .B2(n_404), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_531), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_538), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_566), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_551), .B(n_484), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_554), .Y(n_622) );
NOR2xp67_ASAP7_75t_L g623 ( .A(n_541), .B(n_507), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_586), .A2(n_522), .B(n_515), .Y(n_624) );
BUFx3_ASAP7_75t_L g625 ( .A(n_533), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_551), .B(n_478), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_543), .A2(n_426), .B1(n_404), .B2(n_502), .Y(n_627) );
NAND2x1_ASAP7_75t_L g628 ( .A(n_537), .B(n_501), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_531), .Y(n_629) );
AND2x4_ASAP7_75t_SL g630 ( .A(n_536), .B(n_432), .Y(n_630) );
INVx3_ASAP7_75t_L g631 ( .A(n_528), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_561), .A2(n_522), .B1(n_507), .B2(n_481), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_586), .A2(n_505), .B(n_501), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_553), .A2(n_505), .B(n_501), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_538), .B(n_438), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_533), .Y(n_636) );
CKINVDCx8_ASAP7_75t_R g637 ( .A(n_546), .Y(n_637) );
AO31x2_ASAP7_75t_L g638 ( .A1(n_535), .A2(n_481), .A3(n_483), .B(n_447), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_553), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_562), .A2(n_564), .B(n_563), .Y(n_640) );
CKINVDCx11_ASAP7_75t_R g641 ( .A(n_536), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_534), .B(n_325), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_588), .B(n_505), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_554), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_562), .A2(n_505), .B(n_497), .Y(n_645) );
NOR2xp67_ASAP7_75t_SL g646 ( .A(n_567), .B(n_323), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_543), .A2(n_323), .B1(n_380), .B2(n_337), .Y(n_647) );
INVx5_ASAP7_75t_L g648 ( .A(n_528), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_546), .Y(n_649) );
INVx4_ASAP7_75t_L g650 ( .A(n_552), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_558), .B(n_301), .Y(n_651) );
INVx3_ASAP7_75t_L g652 ( .A(n_528), .Y(n_652) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_567), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_558), .Y(n_654) );
AOI21xp33_ASAP7_75t_L g655 ( .A1(n_559), .A2(n_437), .B(n_436), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_552), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_563), .A2(n_524), .B(n_497), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_579), .B(n_483), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_548), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_579), .B(n_497), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_552), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_552), .Y(n_662) );
OR2x6_ASAP7_75t_L g663 ( .A(n_577), .B(n_524), .Y(n_663) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_592), .Y(n_664) );
OR2x6_ASAP7_75t_L g665 ( .A(n_572), .B(n_524), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_590), .B(n_337), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_564), .A2(n_524), .B(n_519), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_578), .Y(n_668) );
BUFx4_ASAP7_75t_SL g669 ( .A(n_589), .Y(n_669) );
O2A1O1Ixp5_ASAP7_75t_L g670 ( .A1(n_584), .A2(n_330), .B(n_340), .C(n_324), .Y(n_670) );
BUFx4f_ASAP7_75t_SL g671 ( .A(n_547), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_579), .B(n_380), .Y(n_672) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_568), .A2(n_445), .B1(n_364), .B2(n_394), .C1(n_345), .C2(n_360), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_593), .B(n_445), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_580), .A2(n_519), .B(n_488), .Y(n_675) );
INVx3_ASAP7_75t_L g676 ( .A(n_528), .Y(n_676) );
BUFx3_ASAP7_75t_L g677 ( .A(n_533), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_580), .A2(n_519), .B(n_488), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g679 ( .A1(n_572), .A2(n_327), .B(n_325), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_547), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_544), .B(n_451), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_594), .B(n_451), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_591), .B(n_316), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_561), .B(n_327), .Y(n_684) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_533), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_575), .A2(n_519), .B(n_488), .Y(n_686) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_555), .B(n_447), .Y(n_687) );
BUFx3_ASAP7_75t_L g688 ( .A(n_539), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_561), .A2(n_428), .B1(n_443), .B2(n_422), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_547), .B(n_422), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_584), .Y(n_691) );
CKINVDCx5p33_ASAP7_75t_R g692 ( .A(n_649), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_597), .B(n_571), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_691), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_660), .A2(n_582), .B1(n_591), .B2(n_583), .Y(n_695) );
BUFx3_ASAP7_75t_L g696 ( .A(n_602), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_619), .A2(n_587), .B1(n_595), .B2(n_535), .Y(n_697) );
BUFx3_ASAP7_75t_L g698 ( .A(n_602), .Y(n_698) );
BUFx12f_ASAP7_75t_L g699 ( .A(n_649), .Y(n_699) );
BUFx3_ASAP7_75t_L g700 ( .A(n_609), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_630), .A2(n_555), .B1(n_443), .B2(n_428), .Y(n_701) );
AO21x2_ASAP7_75t_L g702 ( .A1(n_681), .A2(n_645), .B(n_684), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_659), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_687), .A2(n_550), .B1(n_569), .B2(n_545), .Y(n_704) );
INVxp67_ASAP7_75t_L g705 ( .A(n_601), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_635), .B(n_578), .Y(n_706) );
OAI21x1_ASAP7_75t_L g707 ( .A1(n_600), .A2(n_585), .B(n_540), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_672), .B(n_578), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_621), .B(n_578), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_599), .B(n_578), .Y(n_710) );
OA21x2_ASAP7_75t_L g711 ( .A1(n_670), .A2(n_550), .B(n_545), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_617), .B(n_532), .Y(n_712) );
INVx5_ASAP7_75t_SL g713 ( .A(n_687), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_642), .A2(n_569), .B1(n_560), .B2(n_542), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_642), .A2(n_576), .B1(n_573), .B2(n_526), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_624), .A2(n_633), .B(n_667), .Y(n_716) );
NAND2xp33_ASAP7_75t_R g717 ( .A(n_669), .B(n_589), .Y(n_717) );
INVx3_ASAP7_75t_L g718 ( .A(n_650), .Y(n_718) );
CKINVDCx6p67_ASAP7_75t_R g719 ( .A(n_641), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_680), .A2(n_526), .B1(n_527), .B2(n_528), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_603), .A2(n_527), .B1(n_530), .B2(n_581), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_612), .A2(n_530), .B1(n_581), .B2(n_589), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_691), .Y(n_723) );
NAND2xp33_ASAP7_75t_R g724 ( .A(n_669), .B(n_589), .Y(n_724) );
OAI21x1_ASAP7_75t_L g725 ( .A1(n_657), .A2(n_585), .B(n_330), .Y(n_725) );
INVxp67_ASAP7_75t_L g726 ( .A(n_610), .Y(n_726) );
BUFx3_ASAP7_75t_L g727 ( .A(n_609), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_612), .A2(n_349), .B1(n_356), .B2(n_346), .C(n_322), .Y(n_728) );
OA21x2_ASAP7_75t_L g729 ( .A1(n_670), .A2(n_640), .B(n_634), .Y(n_729) );
OA21x2_ASAP7_75t_L g730 ( .A1(n_632), .A2(n_340), .B(n_324), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_613), .A2(n_574), .B(n_539), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_650), .Y(n_732) );
NAND3xp33_ASAP7_75t_SL g733 ( .A(n_608), .B(n_338), .C(n_315), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_626), .B(n_530), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_618), .Y(n_735) );
OR2x6_ASAP7_75t_L g736 ( .A(n_607), .B(n_539), .Y(n_736) );
AND2x4_ASAP7_75t_L g737 ( .A(n_656), .B(n_539), .Y(n_737) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_641), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_651), .A2(n_353), .B1(n_366), .B2(n_359), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_614), .B(n_574), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_674), .B(n_574), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_605), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_653), .A2(n_440), .B1(n_338), .B2(n_370), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_627), .A2(n_574), .B1(n_315), .B2(n_379), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_604), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_611), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_618), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_629), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_620), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_671), .A2(n_353), .B1(n_385), .B2(n_371), .Y(n_750) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_614), .Y(n_751) );
INVx8_ASAP7_75t_L g752 ( .A(n_648), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_671), .A2(n_353), .B1(n_406), .B2(n_392), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_616), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_616), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_613), .A2(n_320), .B(n_319), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_666), .A2(n_353), .B1(n_414), .B2(n_413), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_615), .A2(n_353), .B1(n_424), .B2(n_416), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_638), .Y(n_759) );
OR2x6_ASAP7_75t_L g760 ( .A(n_663), .B(n_365), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_658), .A2(n_370), .B1(n_387), .B2(n_379), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g762 ( .A(n_637), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g763 ( .A1(n_690), .A2(n_435), .B1(n_439), .B2(n_434), .C(n_431), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_661), .B(n_449), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_682), .A2(n_410), .B(n_430), .C(n_378), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_615), .A2(n_430), .B1(n_410), .B2(n_304), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_643), .A2(n_343), .B(n_321), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_663), .A2(n_307), .B1(n_308), .B2(n_300), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_638), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_673), .B(n_387), .Y(n_770) );
NAND3xp33_ASAP7_75t_SL g771 ( .A(n_664), .B(n_405), .C(n_396), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_629), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_639), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g774 ( .A1(n_679), .A2(n_306), .B1(n_420), .B2(n_421), .C(n_403), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_647), .B(n_396), .Y(n_775) );
O2A1O1Ixp33_ASAP7_75t_SL g776 ( .A1(n_643), .A2(n_311), .B(n_314), .C(n_312), .Y(n_776) );
INVxp33_ASAP7_75t_SL g777 ( .A(n_646), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_638), .Y(n_778) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_614), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_675), .A2(n_399), .B(n_372), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_689), .B(n_405), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_598), .Y(n_782) );
OR2x2_ASAP7_75t_L g783 ( .A(n_689), .B(n_412), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_663), .A2(n_412), .B1(n_423), .B2(n_408), .Y(n_784) );
AND2x4_ASAP7_75t_L g785 ( .A(n_598), .B(n_317), .Y(n_785) );
A2O1A1Ixp33_ASAP7_75t_L g786 ( .A1(n_632), .A2(n_395), .B(n_390), .C(n_318), .Y(n_786) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_664), .A2(n_409), .B1(n_328), .B2(n_329), .C(n_373), .Y(n_787) );
CKINVDCx8_ASAP7_75t_R g788 ( .A(n_668), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_606), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_638), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_683), .A2(n_352), .B1(n_358), .B2(n_355), .Y(n_791) );
AOI211xp5_ASAP7_75t_L g792 ( .A1(n_733), .A2(n_623), .B(n_655), .C(n_662), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_703), .B(n_713), .Y(n_793) );
OA21x2_ASAP7_75t_L g794 ( .A1(n_759), .A2(n_686), .B(n_678), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_705), .A2(n_683), .B1(n_622), .B2(n_644), .C(n_654), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_725), .A2(n_652), .B(n_631), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_726), .Y(n_797) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_713), .A2(n_665), .B1(n_648), .B2(n_362), .Y(n_798) );
OAI21x1_ASAP7_75t_L g799 ( .A1(n_707), .A2(n_652), .B(n_631), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_770), .A2(n_665), .B1(n_628), .B2(n_423), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_712), .B(n_648), .Y(n_801) );
AOI222xp33_ASAP7_75t_L g802 ( .A1(n_728), .A2(n_398), .B1(n_376), .B2(n_361), .C1(n_381), .C2(n_382), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_717), .Y(n_803) );
OAI22xp33_ASAP7_75t_L g804 ( .A1(n_717), .A2(n_724), .B1(n_760), .B2(n_783), .Y(n_804) );
NAND3xp33_ASAP7_75t_L g805 ( .A(n_765), .B(n_648), .C(n_368), .Y(n_805) );
AOI221xp5_ASAP7_75t_L g806 ( .A1(n_763), .A2(n_419), .B1(n_411), .B2(n_425), .C(n_427), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_764), .Y(n_807) );
OA21x2_ASAP7_75t_L g808 ( .A1(n_769), .A2(n_479), .B(n_452), .Y(n_808) );
OAI21xp5_ASAP7_75t_SL g809 ( .A1(n_701), .A2(n_369), .B(n_367), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_764), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_713), .A2(n_665), .B1(n_362), .B2(n_363), .Y(n_811) );
OA21x2_ASAP7_75t_L g812 ( .A1(n_778), .A2(n_479), .B(n_452), .Y(n_812) );
OAI21x1_ASAP7_75t_L g813 ( .A1(n_716), .A2(n_676), .B(n_479), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_745), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_746), .Y(n_815) );
AOI211xp5_ASAP7_75t_L g816 ( .A1(n_787), .A2(n_375), .B(n_383), .C(n_374), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_735), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_747), .Y(n_818) );
OA21x2_ASAP7_75t_L g819 ( .A1(n_790), .A2(n_786), .B(n_765), .Y(n_819) );
OAI211xp5_ASAP7_75t_L g820 ( .A1(n_704), .A2(n_388), .B(n_389), .C(n_386), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_749), .Y(n_821) );
BUFx3_ASAP7_75t_L g822 ( .A(n_752), .Y(n_822) );
AND2x4_ASAP7_75t_L g823 ( .A(n_718), .B(n_625), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_781), .A2(n_688), .B1(n_677), .B2(n_636), .Y(n_824) );
NOR3xp33_ASAP7_75t_SL g825 ( .A(n_692), .B(n_400), .C(n_397), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_714), .B(n_677), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_748), .Y(n_827) );
AOI222xp33_ASAP7_75t_L g828 ( .A1(n_704), .A2(n_415), .B1(n_441), .B2(n_407), .C1(n_402), .C2(n_433), .Y(n_828) );
BUFx2_ASAP7_75t_L g829 ( .A(n_696), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_785), .Y(n_830) );
OAI22xp33_ASAP7_75t_L g831 ( .A1(n_724), .A2(n_636), .B1(n_685), .B2(n_614), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_760), .A2(n_363), .B1(n_351), .B2(n_688), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_775), .B(n_8), .Y(n_833) );
OAI21xp33_ASAP7_75t_L g834 ( .A1(n_791), .A2(n_351), .B(n_390), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g835 ( .A1(n_729), .A2(n_685), .B(n_636), .Y(n_835) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_752), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_760), .B(n_8), .Y(n_837) );
AOI221x1_ASAP7_75t_L g838 ( .A1(n_786), .A2(n_452), .B1(n_479), .B2(n_480), .C(n_309), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_693), .A2(n_685), .B1(n_395), .B2(n_331), .Y(n_839) );
AND2x4_ASAP7_75t_L g840 ( .A(n_718), .B(n_685), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_772), .Y(n_841) );
INVx3_ASAP7_75t_L g842 ( .A(n_752), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_693), .B(n_9), .Y(n_843) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_729), .A2(n_488), .B(n_485), .Y(n_844) );
AOI22xp33_ASAP7_75t_SL g845 ( .A1(n_738), .A2(n_331), .B1(n_11), .B2(n_9), .Y(n_845) );
AOI222xp33_ASAP7_75t_L g846 ( .A1(n_706), .A2(n_331), .B1(n_480), .B2(n_12), .C1(n_13), .C2(n_14), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_754), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_710), .B(n_10), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_732), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_696), .B(n_10), .Y(n_850) );
AOI221xp5_ASAP7_75t_L g851 ( .A1(n_757), .A2(n_331), .B1(n_480), .B2(n_508), .C(n_516), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_755), .Y(n_852) );
AOI222xp33_ASAP7_75t_L g853 ( .A1(n_709), .A2(n_11), .B1(n_13), .B2(n_14), .C1(n_15), .C2(n_16), .Y(n_853) );
AOI21xp5_ASAP7_75t_L g854 ( .A1(n_729), .A2(n_508), .B(n_485), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_694), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g856 ( .A1(n_715), .A2(n_516), .B1(n_508), .B2(n_485), .C(n_496), .Y(n_856) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_715), .A2(n_741), .B(n_722), .Y(n_857) );
AOI21xp5_ASAP7_75t_SL g858 ( .A1(n_695), .A2(n_730), .B(n_751), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g859 ( .A1(n_721), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_859) );
AOI22xp33_ASAP7_75t_SL g860 ( .A1(n_738), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_708), .A2(n_516), .B1(n_485), .B2(n_496), .Y(n_861) );
AND2x6_ASAP7_75t_SL g862 ( .A(n_719), .B(n_18), .Y(n_862) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_736), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_791), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_777), .A2(n_20), .B1(n_21), .B2(n_23), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_698), .B(n_26), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_768), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_698), .B(n_29), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_723), .Y(n_869) );
OAI211xp5_ASAP7_75t_SL g870 ( .A1(n_750), .A2(n_30), .B(n_31), .C(n_32), .Y(n_870) );
INVx4_ASAP7_75t_L g871 ( .A(n_742), .Y(n_871) );
AND2x4_ASAP7_75t_L g872 ( .A(n_732), .B(n_32), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_761), .A2(n_510), .B1(n_496), .B2(n_492), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_773), .Y(n_874) );
BUFx4f_ASAP7_75t_SL g875 ( .A(n_699), .Y(n_875) );
AO21x2_ASAP7_75t_L g876 ( .A1(n_702), .A2(n_492), .B(n_491), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_753), .A2(n_510), .B1(n_496), .B2(n_492), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_766), .A2(n_33), .B1(n_34), .B2(n_36), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_766), .B(n_36), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_700), .B(n_37), .Y(n_880) );
NAND2x1_ASAP7_75t_L g881 ( .A(n_736), .B(n_491), .Y(n_881) );
AOI221xp5_ASAP7_75t_L g882 ( .A1(n_739), .A2(n_510), .B1(n_496), .B2(n_492), .C(n_491), .Y(n_882) );
OAI22xp33_ASAP7_75t_L g883 ( .A1(n_744), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_727), .A2(n_510), .B1(n_496), .B2(n_492), .Y(n_884) );
AOI21xp33_ASAP7_75t_SL g885 ( .A1(n_762), .A2(n_39), .B(n_40), .Y(n_885) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_739), .A2(n_510), .B1(n_496), .B2(n_492), .C(n_491), .Y(n_886) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_758), .B(n_492), .C(n_491), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_727), .Y(n_888) );
OAI22xp33_ASAP7_75t_L g889 ( .A1(n_697), .A2(n_41), .B1(n_42), .B2(n_44), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_784), .B(n_46), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_807), .A2(n_702), .B1(n_758), .B2(n_736), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_810), .A2(n_730), .B1(n_734), .B2(n_711), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_797), .B(n_771), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_814), .Y(n_894) );
NAND4xp25_ASAP7_75t_SL g895 ( .A(n_860), .B(n_743), .C(n_774), .D(n_788), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_837), .B(n_46), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_815), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_833), .B(n_47), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_806), .B(n_802), .Y(n_899) );
INVx5_ASAP7_75t_L g900 ( .A(n_836), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_822), .B(n_47), .Y(n_901) );
AOI221x1_ASAP7_75t_SL g902 ( .A1(n_865), .A2(n_48), .B1(n_49), .B2(n_50), .C(n_52), .Y(n_902) );
AOI222xp33_ASAP7_75t_L g903 ( .A1(n_806), .A2(n_737), .B1(n_782), .B2(n_789), .C1(n_720), .C2(n_740), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_821), .Y(n_904) );
INVx3_ASAP7_75t_L g905 ( .A(n_836), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_794), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g907 ( .A(n_809), .B(n_782), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_804), .A2(n_737), .B1(n_720), .B2(n_776), .Y(n_908) );
INVx2_ASAP7_75t_L g909 ( .A(n_794), .Y(n_909) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_863), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_836), .Y(n_911) );
AO21x2_ASAP7_75t_L g912 ( .A1(n_835), .A2(n_776), .B(n_740), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_863), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_870), .A2(n_711), .B1(n_767), .B2(n_780), .Y(n_914) );
AOI221xp5_ASAP7_75t_L g915 ( .A1(n_859), .A2(n_756), .B1(n_731), .B2(n_751), .C(n_779), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g916 ( .A(n_800), .B(n_49), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_847), .Y(n_917) );
AOI211xp5_ASAP7_75t_SL g918 ( .A1(n_803), .A2(n_50), .B(n_52), .C(n_53), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_825), .B(n_53), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_811), .A2(n_779), .B1(n_751), .B2(n_58), .Y(n_920) );
OA21x2_ASAP7_75t_L g921 ( .A1(n_835), .A2(n_779), .B(n_751), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_859), .A2(n_779), .B1(n_510), .B2(n_496), .C(n_492), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_852), .Y(n_923) );
AOI21xp5_ASAP7_75t_L g924 ( .A1(n_858), .A2(n_510), .B(n_491), .Y(n_924) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_831), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_867), .A2(n_510), .B1(n_491), .B2(n_58), .C(n_60), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_803), .A2(n_54), .B1(n_57), .B2(n_60), .Y(n_927) );
AND2x4_ASAP7_75t_L g928 ( .A(n_801), .B(n_90), .Y(n_928) );
AOI31xp33_ASAP7_75t_L g929 ( .A1(n_860), .A2(n_57), .A3(n_61), .B(n_62), .Y(n_929) );
INVxp67_ASAP7_75t_L g930 ( .A(n_850), .Y(n_930) );
OA21x2_ASAP7_75t_L g931 ( .A1(n_813), .A2(n_491), .B(n_93), .Y(n_931) );
OR2x2_ASAP7_75t_L g932 ( .A(n_829), .B(n_61), .Y(n_932) );
AOI22xp33_ASAP7_75t_SL g933 ( .A1(n_872), .A2(n_63), .B1(n_65), .B2(n_66), .Y(n_933) );
INVx3_ASAP7_75t_L g934 ( .A(n_842), .Y(n_934) );
AOI22xp33_ASAP7_75t_SL g935 ( .A1(n_872), .A2(n_63), .B1(n_66), .B2(n_67), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_825), .B(n_67), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_795), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_937) );
BUFx2_ASAP7_75t_L g938 ( .A(n_842), .Y(n_938) );
INVx2_ASAP7_75t_SL g939 ( .A(n_823), .Y(n_939) );
AO21x2_ASAP7_75t_L g940 ( .A1(n_876), .A2(n_69), .B(n_70), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_866), .B(n_71), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g942 ( .A1(n_864), .A2(n_72), .B1(n_73), .B2(n_74), .C(n_75), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_874), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_870), .A2(n_72), .B1(n_73), .B2(n_75), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g945 ( .A1(n_889), .A2(n_77), .B1(n_78), .B2(n_79), .C(n_80), .Y(n_945) );
NOR2x1_ASAP7_75t_L g946 ( .A(n_793), .B(n_77), .Y(n_946) );
AO21x1_ASAP7_75t_SL g947 ( .A1(n_824), .A2(n_78), .B(n_82), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_855), .Y(n_948) );
OAI33xp33_ASAP7_75t_L g949 ( .A1(n_878), .A2(n_82), .A3(n_83), .B1(n_84), .B2(n_85), .B3(n_86), .Y(n_949) );
OAI221xp5_ASAP7_75t_L g950 ( .A1(n_845), .A2(n_83), .B1(n_84), .B2(n_85), .C(n_87), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_876), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_811), .A2(n_87), .B1(n_88), .B2(n_89), .Y(n_952) );
BUFx3_ASAP7_75t_L g953 ( .A(n_881), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_832), .A2(n_88), .B1(n_89), .B2(n_91), .Y(n_954) );
OAI22xp33_ASAP7_75t_L g955 ( .A1(n_879), .A2(n_94), .B1(n_97), .B2(n_99), .Y(n_955) );
OR2x2_ASAP7_75t_L g956 ( .A(n_868), .B(n_100), .Y(n_956) );
AND2x4_ASAP7_75t_L g957 ( .A(n_840), .B(n_102), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_880), .B(n_103), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_828), .B(n_109), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_869), .Y(n_960) );
OR2x6_ASAP7_75t_L g961 ( .A(n_823), .B(n_110), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_845), .B(n_114), .Y(n_962) );
INVx1_ASAP7_75t_SL g963 ( .A(n_875), .Y(n_963) );
INVxp67_ASAP7_75t_SL g964 ( .A(n_831), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_853), .A2(n_116), .B1(n_117), .B2(n_118), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_819), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_832), .A2(n_120), .B1(n_123), .B2(n_124), .Y(n_967) );
AND4x1_ASAP7_75t_L g968 ( .A(n_846), .B(n_125), .C(n_127), .D(n_131), .Y(n_968) );
AND2x4_ASAP7_75t_L g969 ( .A(n_840), .B(n_132), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_830), .B(n_298), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_808), .Y(n_971) );
BUFx2_ASAP7_75t_L g972 ( .A(n_849), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_808), .Y(n_973) );
NOR2xp67_ASAP7_75t_L g974 ( .A(n_871), .B(n_137), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_816), .B(n_138), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_817), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_843), .B(n_297), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_795), .A2(n_140), .B1(n_141), .B2(n_142), .Y(n_978) );
AOI221xp5_ASAP7_75t_SL g979 ( .A1(n_885), .A2(n_296), .B1(n_144), .B2(n_147), .C(n_148), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_818), .Y(n_980) );
NOR2x1_ASAP7_75t_L g981 ( .A(n_871), .B(n_143), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_812), .Y(n_982) );
OR2x2_ASAP7_75t_L g983 ( .A(n_888), .B(n_149), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_819), .A2(n_150), .B1(n_152), .B2(n_153), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_827), .Y(n_985) );
NAND2xp5_ASAP7_75t_SL g986 ( .A(n_798), .B(n_157), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_883), .A2(n_159), .B1(n_161), .B2(n_163), .Y(n_987) );
OAI21xp33_ASAP7_75t_SL g988 ( .A1(n_799), .A2(n_166), .B(n_168), .Y(n_988) );
AOI21xp5_ASAP7_75t_L g989 ( .A1(n_844), .A2(n_170), .B(n_174), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g990 ( .A1(n_902), .A2(n_890), .B1(n_834), .B2(n_820), .C(n_792), .Y(n_990) );
INVx1_ASAP7_75t_SL g991 ( .A(n_911), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_917), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_923), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_894), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_897), .B(n_841), .Y(n_995) );
INVxp67_ASAP7_75t_L g996 ( .A(n_901), .Y(n_996) );
OAI33xp33_ASAP7_75t_L g997 ( .A1(n_952), .A2(n_848), .A3(n_805), .B1(n_862), .B2(n_826), .B3(n_887), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_904), .B(n_857), .Y(n_998) );
AOI21xp5_ASAP7_75t_SL g999 ( .A1(n_986), .A2(n_820), .B(n_886), .Y(n_999) );
NOR3xp33_ASAP7_75t_L g1000 ( .A(n_895), .B(n_798), .C(n_849), .Y(n_1000) );
NAND3xp33_ASAP7_75t_L g1001 ( .A(n_918), .B(n_851), .C(n_839), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_966), .B(n_812), .Y(n_1002) );
OR2x2_ASAP7_75t_L g1003 ( .A(n_910), .B(n_844), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_899), .A2(n_886), .B1(n_882), .B2(n_877), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_966), .B(n_796), .Y(n_1005) );
OAI31xp33_ASAP7_75t_SL g1006 ( .A1(n_962), .A2(n_882), .A3(n_856), .B(n_838), .Y(n_1006) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_929), .A2(n_854), .B1(n_861), .B2(n_873), .C(n_884), .Y(n_1007) );
INVx3_ASAP7_75t_L g1008 ( .A(n_953), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_943), .B(n_854), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_893), .B(n_175), .Y(n_1010) );
XOR2x2_ASAP7_75t_L g1011 ( .A(n_963), .B(n_179), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_906), .Y(n_1012) );
INVx1_ASAP7_75t_SL g1013 ( .A(n_900), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_906), .Y(n_1014) );
INVx1_ASAP7_75t_SL g1015 ( .A(n_900), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_948), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_913), .B(n_180), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_909), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_960), .B(n_181), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_976), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_980), .Y(n_1021) );
AOI33xp33_ASAP7_75t_L g1022 ( .A1(n_933), .A2(n_182), .A3(n_185), .B1(n_188), .B2(n_189), .B3(n_190), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_985), .B(n_197), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_896), .B(n_198), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_909), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_951), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_951), .Y(n_1027) );
INVx4_ASAP7_75t_L g1028 ( .A(n_961), .Y(n_1028) );
OAI33xp33_ASAP7_75t_L g1029 ( .A1(n_932), .A2(n_199), .A3(n_201), .B1(n_202), .B2(n_203), .B3(n_205), .Y(n_1029) );
AOI211xp5_ASAP7_75t_SL g1030 ( .A1(n_950), .A2(n_920), .B(n_954), .C(n_916), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_913), .B(n_208), .Y(n_1031) );
NAND3xp33_ASAP7_75t_SL g1032 ( .A(n_935), .B(n_209), .C(n_210), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_930), .B(n_295), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_938), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_971), .B(n_211), .Y(n_1035) );
INVxp67_ASAP7_75t_SL g1036 ( .A(n_971), .Y(n_1036) );
INVx2_ASAP7_75t_L g1037 ( .A(n_973), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_973), .B(n_212), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_982), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_982), .Y(n_1040) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_961), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_941), .B(n_214), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_940), .B(n_215), .Y(n_1043) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_972), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_898), .B(n_216), .Y(n_1045) );
AOI31xp33_ASAP7_75t_L g1046 ( .A1(n_927), .A2(n_217), .A3(n_219), .B(n_220), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_940), .B(n_223), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_946), .Y(n_1048) );
AOI33xp33_ASAP7_75t_L g1049 ( .A1(n_919), .A2(n_224), .A3(n_225), .B1(n_226), .B2(n_227), .B3(n_230), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_965), .A2(n_944), .B1(n_937), .B2(n_978), .Y(n_1050) );
INVxp67_ASAP7_75t_L g1051 ( .A(n_905), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_983), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_892), .B(n_231), .Y(n_1053) );
NOR2x1_ASAP7_75t_L g1054 ( .A(n_981), .B(n_232), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_936), .B(n_907), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_965), .A2(n_233), .B1(n_237), .B2(n_241), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_921), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_907), .B(n_291), .Y(n_1058) );
AOI33xp33_ASAP7_75t_L g1059 ( .A1(n_944), .A2(n_242), .A3(n_243), .B1(n_244), .B2(n_248), .B3(n_249), .Y(n_1059) );
INVx4_ASAP7_75t_L g1060 ( .A(n_900), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_934), .Y(n_1061) );
AOI22xp33_ASAP7_75t_SL g1062 ( .A1(n_925), .A2(n_256), .B1(n_258), .B2(n_259), .Y(n_1062) );
INVx3_ASAP7_75t_L g1063 ( .A(n_953), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_934), .Y(n_1064) );
NAND3xp33_ASAP7_75t_L g1065 ( .A(n_968), .B(n_260), .C(n_261), .Y(n_1065) );
AND2x4_ASAP7_75t_L g1066 ( .A(n_925), .B(n_266), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_928), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_912), .Y(n_1068) );
AND2x4_ASAP7_75t_L g1069 ( .A(n_964), .B(n_267), .Y(n_1069) );
NAND3xp33_ASAP7_75t_L g1070 ( .A(n_945), .B(n_271), .C(n_272), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_892), .B(n_277), .Y(n_1071) );
OR2x2_ASAP7_75t_SL g1072 ( .A(n_956), .B(n_278), .Y(n_1072) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_939), .B(n_279), .Y(n_1073) );
AOI221xp5_ASAP7_75t_L g1074 ( .A1(n_949), .A2(n_942), .B1(n_926), .B2(n_975), .C(n_959), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_921), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_928), .Y(n_1076) );
INVx2_ASAP7_75t_L g1077 ( .A(n_912), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_928), .Y(n_1078) );
INVx2_ASAP7_75t_L g1079 ( .A(n_931), .Y(n_1079) );
OR2x2_ASAP7_75t_L g1080 ( .A(n_939), .B(n_280), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1009), .B(n_964), .Y(n_1081) );
AOI21xp33_ASAP7_75t_L g1082 ( .A1(n_1041), .A2(n_903), .B(n_979), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_992), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_993), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_998), .B(n_891), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_994), .Y(n_1086) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_1044), .B(n_891), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_998), .B(n_900), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1012), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_991), .B(n_958), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1009), .B(n_984), .Y(n_1091) );
HB1xp67_ASAP7_75t_L g1092 ( .A(n_1036), .Y(n_1092) );
NOR2xp67_ASAP7_75t_L g1093 ( .A(n_1028), .B(n_986), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_995), .B(n_908), .Y(n_1094) );
INVx5_ASAP7_75t_L g1095 ( .A(n_1060), .Y(n_1095) );
INVx2_ASAP7_75t_L g1096 ( .A(n_1012), .Y(n_1096) );
OR2x6_ASAP7_75t_L g1097 ( .A(n_1028), .B(n_957), .Y(n_1097) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_1025), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1016), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1055), .B(n_947), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_996), .B(n_969), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1020), .Y(n_1102) );
OR2x2_ASAP7_75t_L g1103 ( .A(n_1021), .B(n_957), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_1025), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1052), .B(n_957), .Y(n_1105) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_1000), .A2(n_974), .B1(n_978), .B2(n_977), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1034), .B(n_969), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1028), .B(n_970), .Y(n_1108) );
NAND2x1_ASAP7_75t_L g1109 ( .A(n_1008), .B(n_931), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1014), .Y(n_1110) );
NAND2x1_ASAP7_75t_L g1111 ( .A(n_1008), .B(n_931), .Y(n_1111) );
INVx1_ASAP7_75t_SL g1112 ( .A(n_1013), .Y(n_1112) );
INVx2_ASAP7_75t_L g1113 ( .A(n_1014), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1002), .B(n_914), .Y(n_1114) );
NOR2xp33_ASAP7_75t_L g1115 ( .A(n_997), .B(n_955), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1061), .Y(n_1116) );
NOR2xp33_ASAP7_75t_R g1117 ( .A(n_1060), .B(n_987), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1005), .B(n_914), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1067), .B(n_915), .Y(n_1119) );
NAND5xp2_ASAP7_75t_L g1120 ( .A(n_1030), .B(n_987), .C(n_922), .D(n_989), .E(n_924), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_1003), .B(n_967), .Y(n_1121) );
AND2x2_ASAP7_75t_SL g1122 ( .A(n_1066), .B(n_955), .Y(n_1122) );
INVxp67_ASAP7_75t_SL g1123 ( .A(n_1026), .Y(n_1123) );
NAND2x1p5_ASAP7_75t_L g1124 ( .A(n_1060), .B(n_988), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1064), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1005), .B(n_285), .Y(n_1126) );
NAND2xp5_ASAP7_75t_SL g1127 ( .A(n_1066), .B(n_286), .Y(n_1127) );
NOR2x1_ASAP7_75t_R g1128 ( .A(n_1011), .B(n_287), .Y(n_1128) );
INVx5_ASAP7_75t_L g1129 ( .A(n_1066), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_1011), .Y(n_1130) );
INVx1_ASAP7_75t_SL g1131 ( .A(n_1015), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1031), .B(n_289), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1017), .Y(n_1133) );
INVxp67_ASAP7_75t_L g1134 ( .A(n_1048), .Y(n_1134) );
NOR2x1_ASAP7_75t_L g1135 ( .A(n_1054), .B(n_290), .Y(n_1135) );
INVx2_ASAP7_75t_L g1136 ( .A(n_1018), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1018), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1076), .B(n_1078), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1051), .B(n_990), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1037), .Y(n_1140) );
NAND2xp33_ASAP7_75t_L g1141 ( .A(n_1065), .B(n_1080), .Y(n_1141) );
OR2x6_ASAP7_75t_L g1142 ( .A(n_1069), .B(n_1063), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1031), .B(n_1063), .Y(n_1143) );
INVxp67_ASAP7_75t_L g1144 ( .A(n_1008), .Y(n_1144) );
BUFx2_ASAP7_75t_L g1145 ( .A(n_1063), .Y(n_1145) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1039), .B(n_1040), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_1122), .A2(n_1050), .B1(n_1074), .B2(n_1029), .Y(n_1147) );
OAI221xp5_ASAP7_75t_L g1148 ( .A1(n_1139), .A2(n_1134), .B1(n_1082), .B2(n_1115), .C(n_1130), .Y(n_1148) );
OAI222xp33_ASAP7_75t_L g1149 ( .A1(n_1097), .A2(n_1069), .B1(n_1080), .B2(n_1073), .C1(n_1043), .C2(n_1047), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1083), .Y(n_1150) );
AOI21xp33_ASAP7_75t_L g1151 ( .A1(n_1115), .A2(n_1010), .B(n_1033), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1084), .Y(n_1152) );
NAND4xp25_ASAP7_75t_L g1153 ( .A(n_1120), .B(n_1024), .C(n_1058), .D(n_1045), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1086), .Y(n_1154) );
NAND2xp5_ASAP7_75t_SL g1155 ( .A(n_1122), .B(n_1069), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1099), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1143), .B(n_1040), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1102), .Y(n_1158) );
AOI21xp33_ASAP7_75t_L g1159 ( .A1(n_1134), .A2(n_1046), .B(n_1042), .Y(n_1159) );
A2O1A1Ixp33_ASAP7_75t_L g1160 ( .A1(n_1129), .A2(n_1049), .B(n_1059), .C(n_1022), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1116), .Y(n_1161) );
NAND4xp75_ASAP7_75t_L g1162 ( .A(n_1093), .B(n_1047), .C(n_1043), .D(n_1053), .Y(n_1162) );
NOR2x1p5_ASAP7_75t_L g1163 ( .A(n_1130), .B(n_1032), .Y(n_1163) );
AOI22x1_ASAP7_75t_L g1164 ( .A1(n_1112), .A2(n_1073), .B1(n_1072), .B2(n_1053), .Y(n_1164) );
AOI322xp5_ASAP7_75t_L g1165 ( .A1(n_1100), .A2(n_1019), .A3(n_1071), .B1(n_1004), .B2(n_1007), .C1(n_1023), .C2(n_1056), .Y(n_1165) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_1097), .A2(n_1001), .B1(n_1019), .B2(n_1070), .Y(n_1166) );
OAI21xp5_ASAP7_75t_L g1167 ( .A1(n_1127), .A2(n_999), .B(n_1049), .Y(n_1167) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1089), .Y(n_1168) );
INVx1_ASAP7_75t_SL g1169 ( .A(n_1131), .Y(n_1169) );
AND2x4_ASAP7_75t_L g1170 ( .A(n_1142), .B(n_1057), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1089), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1125), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1085), .B(n_1027), .Y(n_1173) );
OR2x2_ASAP7_75t_L g1174 ( .A(n_1092), .B(n_1057), .Y(n_1174) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_1097), .A2(n_1072), .B1(n_1142), .B2(n_1129), .Y(n_1175) );
OAI21xp5_ASAP7_75t_L g1176 ( .A1(n_1127), .A2(n_999), .B(n_1022), .Y(n_1176) );
OAI221xp5_ASAP7_75t_L g1177 ( .A1(n_1106), .A2(n_1062), .B1(n_1006), .B2(n_1068), .C(n_1075), .Y(n_1177) );
AOI22xp5_ASAP7_75t_L g1178 ( .A1(n_1101), .A2(n_1023), .B1(n_1035), .B2(n_1038), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1098), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1098), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1104), .Y(n_1181) );
O2A1O1Ixp33_ASAP7_75t_SL g1182 ( .A1(n_1128), .A2(n_1075), .B(n_1059), .C(n_1079), .Y(n_1182) );
AOI22xp33_ASAP7_75t_SL g1183 ( .A1(n_1129), .A2(n_1035), .B1(n_1038), .B2(n_1079), .Y(n_1183) );
AOI21xp33_ASAP7_75t_L g1184 ( .A1(n_1087), .A2(n_1077), .B(n_1144), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1088), .Y(n_1185) );
OAI22xp33_ASAP7_75t_L g1186 ( .A1(n_1142), .A2(n_1077), .B1(n_1129), .B2(n_1095), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1150), .Y(n_1187) );
INVx2_ASAP7_75t_SL g1188 ( .A(n_1174), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1185), .B(n_1118), .Y(n_1189) );
NAND3xp33_ASAP7_75t_L g1190 ( .A(n_1148), .B(n_1144), .C(n_1141), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1152), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1154), .Y(n_1192) );
XNOR2x2_ASAP7_75t_L g1193 ( .A(n_1155), .B(n_1090), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1157), .B(n_1114), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1156), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1173), .B(n_1146), .Y(n_1196) );
CKINVDCx5p33_ASAP7_75t_R g1197 ( .A(n_1169), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1158), .Y(n_1198) );
OAI21xp33_ASAP7_75t_L g1199 ( .A1(n_1147), .A2(n_1117), .B(n_1114), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1170), .B(n_1081), .Y(n_1200) );
NOR2xp33_ASAP7_75t_L g1201 ( .A(n_1151), .B(n_1105), .Y(n_1201) );
AOI21xp33_ASAP7_75t_SL g1202 ( .A1(n_1155), .A2(n_1124), .B(n_1103), .Y(n_1202) );
AOI21xp33_ASAP7_75t_L g1203 ( .A1(n_1147), .A2(n_1108), .B(n_1119), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1161), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1179), .B(n_1133), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1172), .Y(n_1206) );
NAND4xp75_ASAP7_75t_L g1207 ( .A(n_1167), .B(n_1135), .C(n_1132), .D(n_1126), .Y(n_1207) );
NOR2x1_ASAP7_75t_L g1208 ( .A(n_1175), .B(n_1145), .Y(n_1208) );
AOI21xp5_ASAP7_75t_L g1209 ( .A1(n_1182), .A2(n_1095), .B(n_1124), .Y(n_1209) );
INVx3_ASAP7_75t_L g1210 ( .A(n_1170), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1180), .Y(n_1211) );
NOR2x1_ASAP7_75t_L g1212 ( .A(n_1176), .B(n_1126), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1181), .Y(n_1213) );
XNOR2x2_ASAP7_75t_L g1214 ( .A(n_1193), .B(n_1162), .Y(n_1214) );
AOI221xp5_ASAP7_75t_L g1215 ( .A1(n_1203), .A2(n_1184), .B1(n_1159), .B2(n_1182), .C(n_1177), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_1199), .A2(n_1163), .B1(n_1153), .B2(n_1166), .Y(n_1216) );
AOI21xp5_ASAP7_75t_L g1217 ( .A1(n_1209), .A2(n_1160), .B(n_1149), .Y(n_1217) );
NAND2xp5_ASAP7_75t_SL g1218 ( .A(n_1208), .B(n_1197), .Y(n_1218) );
CKINVDCx16_ASAP7_75t_R g1219 ( .A(n_1212), .Y(n_1219) );
NAND2x1_ASAP7_75t_L g1220 ( .A(n_1210), .B(n_1188), .Y(n_1220) );
AOI31xp33_ASAP7_75t_L g1221 ( .A1(n_1197), .A2(n_1160), .A3(n_1186), .B(n_1183), .Y(n_1221) );
NAND2xp5_ASAP7_75t_SL g1222 ( .A(n_1202), .B(n_1164), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g1223 ( .A1(n_1201), .A2(n_1094), .B1(n_1107), .B2(n_1178), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1196), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1196), .Y(n_1225) );
INVx2_ASAP7_75t_SL g1226 ( .A(n_1188), .Y(n_1226) );
AO22x2_ASAP7_75t_L g1227 ( .A1(n_1187), .A2(n_1171), .B1(n_1168), .B2(n_1138), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1227), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1227), .Y(n_1229) );
AND2x4_ASAP7_75t_L g1230 ( .A(n_1218), .B(n_1210), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_1215), .A2(n_1201), .B1(n_1190), .B2(n_1206), .Y(n_1231) );
HB1xp67_ASAP7_75t_L g1232 ( .A(n_1220), .Y(n_1232) );
AOI21xp5_ASAP7_75t_L g1233 ( .A1(n_1222), .A2(n_1149), .B(n_1186), .Y(n_1233) );
O2A1O1Ixp33_ASAP7_75t_L g1234 ( .A1(n_1221), .A2(n_1198), .B(n_1191), .C(n_1192), .Y(n_1234) );
NOR2xp33_ASAP7_75t_R g1235 ( .A(n_1219), .B(n_1095), .Y(n_1235) );
OAI322xp33_ASAP7_75t_L g1236 ( .A1(n_1214), .A2(n_1189), .A3(n_1204), .B1(n_1195), .B2(n_1205), .C1(n_1213), .C2(n_1211), .Y(n_1236) );
NOR2x1_ASAP7_75t_L g1237 ( .A(n_1217), .B(n_1207), .Y(n_1237) );
NAND4xp25_ASAP7_75t_L g1238 ( .A(n_1216), .B(n_1165), .C(n_1121), .D(n_1183), .Y(n_1238) );
NAND3xp33_ASAP7_75t_SL g1239 ( .A(n_1216), .B(n_1117), .C(n_1109), .Y(n_1239) );
OAI21xp33_ASAP7_75t_SL g1240 ( .A1(n_1226), .A2(n_1194), .B(n_1200), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1224), .Y(n_1241) );
AOI221xp5_ASAP7_75t_L g1242 ( .A1(n_1225), .A2(n_1091), .B1(n_1168), .B2(n_1171), .C(n_1140), .Y(n_1242) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_1223), .A2(n_1123), .B1(n_1111), .B2(n_1137), .Y(n_1243) );
NOR2xp33_ASAP7_75t_L g1244 ( .A(n_1236), .B(n_1231), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1231), .B(n_1233), .Y(n_1245) );
OAI221xp5_ASAP7_75t_L g1246 ( .A1(n_1237), .A2(n_1234), .B1(n_1238), .B2(n_1240), .C(n_1232), .Y(n_1246) );
AO22x2_ASAP7_75t_L g1247 ( .A1(n_1245), .A2(n_1229), .B1(n_1228), .B2(n_1239), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1247), .Y(n_1248) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_1248), .A2(n_1244), .B1(n_1246), .B2(n_1230), .C(n_1243), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g1250 ( .A1(n_1249), .A2(n_1235), .B1(n_1241), .B2(n_1242), .Y(n_1250) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_1250), .A2(n_1096), .B1(n_1110), .B2(n_1113), .C(n_1136), .Y(n_1251) );
endmodule