module fake_aes_3140_n_463 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_463);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_463;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_73;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_67;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g66 ( .A(n_34), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_52), .Y(n_67) );
INVx1_ASAP7_75t_SL g68 ( .A(n_51), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_50), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_23), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_15), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_38), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_45), .Y(n_73) );
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_40), .Y(n_74) );
INVxp33_ASAP7_75t_L g75 ( .A(n_11), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_64), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_5), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_20), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_21), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_42), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_6), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_57), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_32), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_10), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_65), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_49), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
INVx2_ASAP7_75t_SL g88 ( .A(n_18), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_3), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_1), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_41), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_58), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_62), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_21), .Y(n_94) );
INVxp67_ASAP7_75t_L g95 ( .A(n_25), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_53), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_37), .Y(n_98) );
INVx1_ASAP7_75t_SL g99 ( .A(n_4), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_39), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_77), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_74), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_66), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_68), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_88), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_98), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_88), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_98), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_99), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_70), .B(n_0), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_83), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_95), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_90), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_85), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_86), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_71), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_67), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_100), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_87), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_71), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_120), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_120), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_105), .B(n_100), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_112), .B(n_69), .Y(n_126) );
OAI22xp33_ASAP7_75t_SL g127 ( .A1(n_111), .A2(n_81), .B1(n_96), .B2(n_78), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_122), .A2(n_75), .B1(n_96), .B2(n_81), .Y(n_128) );
OR2x2_ASAP7_75t_SL g129 ( .A(n_110), .B(n_78), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_116), .B(n_79), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_103), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_106), .B(n_69), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_122), .A2(n_114), .B1(n_115), .B2(n_117), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_120), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_120), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_120), .Y(n_136) );
NAND2x1p5_ASAP7_75t_L g137 ( .A(n_105), .B(n_72), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_116), .B(n_79), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_120), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_119), .B(n_72), .Y(n_140) );
OR2x6_ASAP7_75t_L g141 ( .A(n_111), .B(n_89), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_119), .B(n_89), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_107), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_101), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_107), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_138), .B(n_113), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_141), .B(n_108), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_141), .Y(n_148) );
NOR2xp33_ASAP7_75t_R g149 ( .A(n_131), .B(n_110), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_141), .Y(n_150) );
OAI21xp5_ASAP7_75t_L g151 ( .A1(n_137), .A2(n_121), .B(n_93), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_141), .B(n_84), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_138), .B(n_104), .Y(n_154) );
OR2x2_ASAP7_75t_L g155 ( .A(n_131), .B(n_102), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_138), .B(n_94), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_138), .B(n_130), .Y(n_157) );
OR2x2_ASAP7_75t_L g158 ( .A(n_133), .B(n_102), .Y(n_158) );
NOR3xp33_ASAP7_75t_SL g159 ( .A(n_128), .B(n_92), .C(n_97), .Y(n_159) );
NAND3xp33_ASAP7_75t_L g160 ( .A(n_132), .B(n_91), .C(n_76), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_137), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_137), .Y(n_162) );
NOR3xp33_ASAP7_75t_L g163 ( .A(n_128), .B(n_91), .C(n_76), .Y(n_163) );
OAI21xp33_ASAP7_75t_L g164 ( .A1(n_130), .A2(n_107), .B(n_109), .Y(n_164) );
AND3x1_ASAP7_75t_SL g165 ( .A(n_129), .B(n_118), .C(n_97), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_132), .B(n_109), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_145), .Y(n_167) );
INVx2_ASAP7_75t_SL g168 ( .A(n_142), .Y(n_168) );
AND3x1_ASAP7_75t_SL g169 ( .A(n_129), .B(n_73), .C(n_80), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_145), .Y(n_171) );
INVxp67_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
OR2x6_ASAP7_75t_SL g173 ( .A(n_140), .B(n_93), .Y(n_173) );
BUFx4f_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_126), .B(n_109), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_167), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_161), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_157), .B(n_140), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_147), .B(n_127), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_157), .A2(n_127), .B1(n_143), .B2(n_125), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_149), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_151), .A2(n_143), .B(n_125), .C(n_145), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_157), .B(n_143), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_168), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_174), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_167), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_166), .A2(n_136), .B(n_123), .Y(n_189) );
INVx6_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_167), .Y(n_191) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_171), .A2(n_139), .B(n_135), .Y(n_192) );
BUFx10_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_152), .A2(n_145), .B1(n_73), .B2(n_80), .Y(n_194) );
OAI221xp5_ASAP7_75t_L g195 ( .A1(n_163), .A2(n_82), .B1(n_145), .B2(n_136), .C(n_123), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_152), .A2(n_145), .B1(n_82), .B2(n_135), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_146), .B(n_0), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_148), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_174), .A2(n_139), .B(n_135), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_147), .B(n_139), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_174), .B(n_134), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_150), .B(n_1), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_173), .B(n_2), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_156), .B(n_2), .Y(n_205) );
INVxp67_ASAP7_75t_SL g206 ( .A(n_205), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_204), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g208 ( .A(n_193), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_178), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_178), .B(n_155), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_189), .A2(n_154), .B(n_171), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_191), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_179), .B(n_173), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_190), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_193), .B(n_149), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_205), .A2(n_172), .B1(n_159), .B2(n_156), .Y(n_216) );
OAI22xp33_ASAP7_75t_L g217 ( .A1(n_182), .A2(n_158), .B1(n_155), .B2(n_170), .Y(n_217) );
OR2x6_ASAP7_75t_L g218 ( .A(n_178), .B(n_156), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_179), .B(n_175), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_181), .B(n_175), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_205), .Y(n_221) );
AOI221xp5_ASAP7_75t_L g222 ( .A1(n_181), .A2(n_158), .B1(n_175), .B2(n_160), .C(n_164), .Y(n_222) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_183), .A2(n_169), .B(n_165), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_204), .Y(n_224) );
AOI221xp5_ASAP7_75t_L g225 ( .A1(n_180), .A2(n_167), .B1(n_134), .B2(n_124), .C(n_6), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_184), .B(n_3), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g227 ( .A(n_205), .B(n_134), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_205), .A2(n_124), .B1(n_134), .B2(n_7), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_203), .A2(n_134), .B1(n_124), .B2(n_7), .Y(n_229) );
OAI211xp5_ASAP7_75t_L g230 ( .A1(n_216), .A2(n_203), .B(n_197), .C(n_194), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_213), .A2(n_203), .B1(n_202), .B2(n_190), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_206), .A2(n_202), .B1(n_185), .B2(n_187), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_211), .A2(n_189), .B(n_199), .Y(n_233) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_220), .A2(n_199), .B(n_192), .Y(n_234) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_228), .A2(n_192), .B(n_176), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_213), .B(n_177), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_221), .B(n_177), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_207), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_212), .Y(n_239) );
AOI221xp5_ASAP7_75t_L g240 ( .A1(n_217), .A2(n_187), .B1(n_185), .B2(n_195), .C(n_184), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_208), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g242 ( .A1(n_221), .A2(n_202), .B1(n_193), .B2(n_190), .Y(n_242) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_222), .A2(n_195), .B1(n_184), .B2(n_202), .C(n_194), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_216), .A2(n_202), .B1(n_190), .B2(n_200), .Y(n_245) );
OAI21xp5_ASAP7_75t_SL g246 ( .A1(n_227), .A2(n_186), .B(n_196), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_212), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_210), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_227), .A2(n_190), .B1(n_200), .B2(n_196), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_239), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_238), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_239), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_241), .Y(n_253) );
OAI211xp5_ASAP7_75t_SL g254 ( .A1(n_240), .A2(n_210), .B(n_229), .C(n_226), .Y(n_254) );
OAI33xp33_ASAP7_75t_L g255 ( .A1(n_238), .A2(n_228), .A3(n_224), .B1(n_215), .B2(n_219), .B3(n_201), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_239), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_236), .B(n_227), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_236), .B(n_224), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_239), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_232), .A2(n_218), .B1(n_208), .B2(n_209), .Y(n_260) );
INVxp67_ASAP7_75t_L g261 ( .A(n_248), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_244), .B(n_223), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
OAI31xp33_ASAP7_75t_L g264 ( .A1(n_230), .A2(n_186), .A3(n_214), .B(n_198), .Y(n_264) );
OAI31xp33_ASAP7_75t_L g265 ( .A1(n_230), .A2(n_186), .A3(n_214), .B(n_198), .Y(n_265) );
OAI221xp5_ASAP7_75t_L g266 ( .A1(n_240), .A2(n_218), .B1(n_225), .B2(n_200), .C(n_214), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_244), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_234), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_234), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_268), .B(n_234), .Y(n_270) );
NOR2x1_ASAP7_75t_SL g271 ( .A(n_260), .B(n_246), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_251), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_251), .B(n_236), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_267), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_250), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_267), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g277 ( .A1(n_261), .A2(n_231), .B1(n_245), .B2(n_243), .C(n_246), .Y(n_277) );
NAND2x1p5_ASAP7_75t_L g278 ( .A(n_256), .B(n_239), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_250), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_262), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_268), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_268), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_262), .Y(n_283) );
INVx4_ASAP7_75t_L g284 ( .A(n_250), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_269), .B(n_234), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_269), .B(n_233), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_260), .B(n_264), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_269), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_252), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_263), .B(n_233), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_266), .A2(n_243), .B1(n_223), .B2(n_241), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_259), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_258), .B(n_237), .Y(n_294) );
AOI322xp5_ASAP7_75t_L g295 ( .A1(n_258), .A2(n_241), .A3(n_232), .B1(n_242), .B2(n_237), .C1(n_10), .C2(n_11), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_252), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_258), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_256), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_286), .B(n_257), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_297), .B(n_261), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_286), .B(n_257), .Y(n_301) );
NAND4xp25_ASAP7_75t_SL g302 ( .A(n_295), .B(n_266), .C(n_265), .D(n_264), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g303 ( .A(n_295), .B(n_265), .C(n_253), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_289), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_280), .B(n_257), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_289), .Y(n_306) );
AND2x2_ASAP7_75t_SL g307 ( .A(n_284), .B(n_237), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_272), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_286), .B(n_259), .Y(n_309) );
CKINVDCx16_ASAP7_75t_R g310 ( .A(n_294), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_270), .B(n_259), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_294), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_297), .B(n_253), .Y(n_313) );
NOR4xp25_ASAP7_75t_SL g314 ( .A(n_288), .B(n_254), .C(n_255), .D(n_223), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g315 ( .A(n_294), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_280), .B(n_259), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_283), .B(n_263), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_270), .B(n_263), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_270), .B(n_263), .Y(n_320) );
NOR2xp33_ASAP7_75t_SL g321 ( .A(n_284), .B(n_241), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_273), .B(n_242), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_274), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_290), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_285), .B(n_263), .Y(n_325) );
AOI31xp33_ASAP7_75t_L g326 ( .A1(n_292), .A2(n_255), .A3(n_249), .B(n_254), .Y(n_326) );
AO21x2_ASAP7_75t_L g327 ( .A1(n_291), .A2(n_235), .B(n_249), .Y(n_327) );
NOR4xp25_ASAP7_75t_SL g328 ( .A(n_277), .B(n_4), .C(n_5), .D(n_8), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_285), .B(n_256), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_273), .B(n_256), .Y(n_330) );
OR2x6_ASAP7_75t_L g331 ( .A(n_284), .B(n_275), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_290), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_274), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_283), .B(n_235), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_296), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_276), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_287), .B(n_235), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_276), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_287), .B(n_9), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_281), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_324), .Y(n_341) );
NOR4xp25_ASAP7_75t_L g342 ( .A(n_302), .B(n_277), .C(n_292), .D(n_296), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_332), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_310), .B(n_281), .Y(n_344) );
AOI32xp33_ASAP7_75t_L g345 ( .A1(n_312), .A2(n_284), .A3(n_285), .B1(n_279), .B2(n_275), .Y(n_345) );
OAI33xp33_ASAP7_75t_L g346 ( .A1(n_300), .A2(n_281), .A3(n_282), .B1(n_271), .B2(n_293), .B3(n_15), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_315), .B(n_271), .Y(n_347) );
AOI211xp5_ASAP7_75t_L g348 ( .A1(n_303), .A2(n_291), .B(n_279), .C(n_275), .Y(n_348) );
OAI322xp33_ASAP7_75t_L g349 ( .A1(n_339), .A2(n_282), .A3(n_293), .B1(n_298), .B2(n_278), .C1(n_16), .C2(n_17), .Y(n_349) );
OAI311xp33_ASAP7_75t_L g350 ( .A1(n_339), .A2(n_298), .A3(n_12), .B1(n_13), .C1(n_14), .Y(n_350) );
NAND2x1_ASAP7_75t_L g351 ( .A(n_331), .B(n_282), .Y(n_351) );
NAND2xp33_ASAP7_75t_L g352 ( .A(n_319), .B(n_298), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_307), .A2(n_298), .B1(n_291), .B2(n_293), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_335), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_299), .B(n_291), .Y(n_355) );
O2A1O1Ixp33_ASAP7_75t_L g356 ( .A1(n_326), .A2(n_218), .B(n_200), .C(n_291), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_307), .A2(n_218), .B1(n_200), .B2(n_278), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_340), .Y(n_358) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_314), .B(n_124), .C(n_134), .Y(n_359) );
OAI31xp33_ASAP7_75t_L g360 ( .A1(n_321), .A2(n_278), .A3(n_198), .B(n_13), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_299), .B(n_278), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_322), .A2(n_218), .B1(n_200), .B2(n_193), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_313), .B(n_9), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_331), .A2(n_193), .B1(n_198), .B2(n_247), .Y(n_364) );
NAND3xp33_ASAP7_75t_SL g365 ( .A(n_328), .B(n_12), .C(n_14), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_333), .A2(n_124), .B1(n_17), .B2(n_18), .C(n_19), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_336), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_338), .Y(n_368) );
AO21x1_ASAP7_75t_L g369 ( .A1(n_338), .A2(n_16), .B(n_19), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_301), .B(n_20), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_301), .B(n_22), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_308), .B(n_22), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_331), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_331), .A2(n_247), .B1(n_239), .B2(n_212), .Y(n_374) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_334), .A2(n_24), .B(n_124), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_319), .A2(n_247), .B1(n_212), .B2(n_188), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_319), .A2(n_247), .B(n_212), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_323), .B(n_305), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_305), .B(n_24), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_304), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_311), .B(n_247), .Y(n_381) );
CKINVDCx14_ASAP7_75t_R g382 ( .A(n_329), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_330), .A2(n_247), .B1(n_188), .B2(n_176), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_340), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_344), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_341), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_343), .B(n_304), .Y(n_387) );
NOR3xp33_ASAP7_75t_SL g388 ( .A(n_346), .B(n_306), .C(n_327), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_354), .B(n_306), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_382), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_358), .Y(n_391) );
XNOR2x2_ASAP7_75t_L g392 ( .A(n_370), .B(n_317), .Y(n_392) );
NOR4xp25_ASAP7_75t_SL g393 ( .A(n_375), .B(n_327), .C(n_334), .D(n_337), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_378), .B(n_309), .Y(n_394) );
AND3x2_ASAP7_75t_L g395 ( .A(n_348), .B(n_318), .C(n_320), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_373), .B(n_318), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_358), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_346), .B(n_337), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_367), .Y(n_399) );
NAND3xp33_ASAP7_75t_L g400 ( .A(n_342), .B(n_316), .C(n_325), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_371), .B(n_316), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_368), .B(n_247), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_355), .B(n_26), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_361), .B(n_27), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_380), .B(n_28), .Y(n_405) );
NAND2x1_ASAP7_75t_L g406 ( .A(n_347), .B(n_188), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_SL g407 ( .A1(n_363), .A2(n_176), .B(n_30), .C(n_31), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_384), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_351), .Y(n_409) );
NOR3xp33_ASAP7_75t_SL g410 ( .A(n_350), .B(n_29), .C(n_33), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_381), .B(n_35), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_372), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_379), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_352), .Y(n_414) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_356), .B(n_191), .C(n_36), .Y(n_415) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_349), .B(n_191), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_369), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_398), .B(n_345), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_390), .A2(n_353), .B1(n_364), .B2(n_374), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_417), .B(n_365), .C(n_366), .Y(n_420) );
O2A1O1Ixp5_ASAP7_75t_L g421 ( .A1(n_398), .A2(n_376), .B(n_377), .C(n_359), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_400), .A2(n_365), .B1(n_357), .B2(n_360), .C(n_362), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_390), .A2(n_383), .B(n_192), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_387), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_385), .Y(n_425) );
OAI321xp33_ASAP7_75t_L g426 ( .A1(n_415), .A2(n_191), .A3(n_44), .B1(n_46), .B2(n_47), .C(n_48), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_389), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_392), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_412), .B(n_43), .Y(n_429) );
OA22x2_ASAP7_75t_L g430 ( .A1(n_395), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_430) );
XNOR2x1_ASAP7_75t_L g431 ( .A(n_392), .B(n_59), .Y(n_431) );
AOI22xp5_ASAP7_75t_SL g432 ( .A1(n_391), .A2(n_60), .B1(n_61), .B2(n_191), .Y(n_432) );
AOI322xp5_ASAP7_75t_L g433 ( .A1(n_388), .A2(n_413), .A3(n_397), .B1(n_401), .B2(n_386), .C1(n_394), .C2(n_414), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_406), .A2(n_407), .B(n_416), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_399), .Y(n_435) );
NOR2x1p5_ASAP7_75t_L g436 ( .A(n_409), .B(n_412), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_428), .A2(n_410), .B1(n_396), .B2(n_409), .C(n_403), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_431), .A2(n_396), .B1(n_393), .B2(n_404), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_425), .Y(n_439) );
INVx3_ASAP7_75t_SL g440 ( .A(n_432), .Y(n_440) );
OAI322xp33_ASAP7_75t_L g441 ( .A1(n_419), .A2(n_408), .A3(n_402), .B1(n_405), .B2(n_404), .C1(n_411), .C2(n_407), .Y(n_441) );
NAND2xp33_ASAP7_75t_SL g442 ( .A(n_436), .B(n_411), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_433), .B(n_427), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_430), .A2(n_422), .B1(n_434), .B2(n_424), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_420), .A2(n_421), .B1(n_435), .B2(n_423), .C(n_429), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_430), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_426), .B(n_421), .C(n_428), .Y(n_447) );
NAND3xp33_ASAP7_75t_SL g448 ( .A(n_433), .B(n_421), .C(n_434), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_419), .A2(n_418), .B1(n_431), .B2(n_428), .Y(n_449) );
NOR2xp67_ASAP7_75t_SL g450 ( .A(n_434), .B(n_390), .Y(n_450) );
NOR3xp33_ASAP7_75t_L g451 ( .A(n_421), .B(n_428), .C(n_420), .Y(n_451) );
NAND2x1p5_ASAP7_75t_SL g452 ( .A(n_450), .B(n_448), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_439), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_449), .A2(n_440), .B1(n_443), .B2(n_444), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_439), .B(n_451), .Y(n_455) );
AO22x2_ASAP7_75t_L g456 ( .A1(n_454), .A2(n_447), .B1(n_446), .B2(n_438), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_453), .Y(n_457) );
NOR4xp25_ASAP7_75t_SL g458 ( .A(n_452), .B(n_442), .C(n_445), .D(n_437), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_457), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_456), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_460), .B(n_455), .Y(n_461) );
OAI221xp5_ASAP7_75t_R g462 ( .A1(n_461), .A2(n_456), .B1(n_458), .B2(n_455), .C(n_459), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_462), .A2(n_442), .B(n_441), .Y(n_463) );
endmodule