module fake_jpeg_27687_n_167 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_30),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_45),
.Y(n_61)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_1),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_26),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_48),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_31),
.B1(n_26),
.B2(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_23),
.B1(n_27),
.B2(n_9),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_57),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_16),
.Y(n_71)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_46),
.C(n_2),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_21),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_68),
.Y(n_77)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_52),
.B1(n_58),
.B2(n_49),
.Y(n_90)
);

OAI32xp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_38),
.A3(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_80),
.B1(n_86),
.B2(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_12),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_19),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_74),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_28),
.B(n_22),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_39),
.B1(n_28),
.B2(n_14),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_1),
.B(n_3),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_29),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_64),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_27),
.B(n_7),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_89),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_6),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_12),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_74),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_50),
.B1(n_68),
.B2(n_55),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_99),
.B1(n_94),
.B2(n_92),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_50),
.B1(n_55),
.B2(n_13),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_73),
.C(n_87),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_105),
.C(n_106),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_88),
.B(n_70),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_96),
.B(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_72),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_122),
.B(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_116),
.C(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_113),
.B1(n_117),
.B2(n_111),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_105),
.C(n_96),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_126),
.C(n_135),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_106),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_130),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_102),
.B(n_77),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_144),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.C(n_112),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_127),
.B1(n_134),
.B2(n_136),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_151),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_131),
.C(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_152),
.Y(n_153)
);

AOI321xp33_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_133),
.A3(n_123),
.B1(n_128),
.B2(n_89),
.C(n_107),
.Y(n_148)
);

NOR4xp25_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_97),
.C(n_119),
.D(n_107),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_141),
.B(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_155),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

AOI31xp67_ASAP7_75t_SL g158 ( 
.A1(n_156),
.A2(n_119),
.A3(n_139),
.B(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_161),
.Y(n_163)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_159),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_157),
.B(n_114),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_160),
.C(n_149),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.C(n_76),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_144),
.C(n_138),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_76),
.Y(n_167)
);


endmodule