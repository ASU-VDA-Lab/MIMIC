module fake_jpeg_6276_n_231 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_2),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_26),
.Y(n_37)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_13),
.B1(n_20),
.B2(n_21),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_12),
.B1(n_22),
.B2(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_42),
.B1(n_23),
.B2(n_14),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_21),
.B1(n_25),
.B2(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_12),
.B1(n_22),
.B2(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_41),
.B1(n_28),
.B2(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_56),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_28),
.B1(n_41),
.B2(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_57),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_31),
.C(n_24),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_19),
.C(n_31),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_21),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_70),
.B(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_78),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_18),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_53),
.C(n_56),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_54),
.B1(n_28),
.B2(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_91),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_94),
.B1(n_51),
.B2(n_62),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_90),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_54),
.B1(n_60),
.B2(n_44),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_85),
.B1(n_77),
.B2(n_67),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_60),
.B1(n_38),
.B2(n_27),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_69),
.B(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_38),
.B1(n_39),
.B2(n_24),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_98),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_68),
.B1(n_64),
.B2(n_65),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_101),
.B1(n_102),
.B2(n_110),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_64),
.B1(n_67),
.B2(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_108),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_76),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_74),
.B1(n_70),
.B2(n_71),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_117),
.C(n_43),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_81),
.C(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_89),
.B(n_93),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_129),
.B(n_16),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_80),
.B1(n_82),
.B2(n_79),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_126),
.B1(n_19),
.B2(n_71),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_85),
.B1(n_81),
.B2(n_44),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_62),
.B1(n_13),
.B2(n_36),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_85),
.B1(n_49),
.B2(n_12),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_72),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_22),
.B(n_19),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_102),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_130),
.A2(n_72),
.B(n_18),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g131 ( 
.A(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_99),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_122),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_95),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_141),
.C(n_147),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_139),
.B(n_140),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_75),
.B1(n_36),
.B2(n_29),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_75),
.B(n_29),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_149),
.B1(n_152),
.B2(n_13),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_36),
.B1(n_40),
.B2(n_17),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_59),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_62),
.B1(n_13),
.B2(n_17),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_17),
.B1(n_62),
.B2(n_15),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_126),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_59),
.C(n_52),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_127),
.C(n_114),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_13),
.B1(n_17),
.B2(n_15),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVxp33_ASAP7_75t_SL g155 ( 
.A(n_144),
.Y(n_155)
);

AO221x1_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_143),
.B1(n_146),
.B2(n_149),
.C(n_3),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_167),
.C(n_152),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_132),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_163),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_120),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_118),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_116),
.B1(n_129),
.B2(n_52),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_116),
.Y(n_166)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_147),
.C(n_151),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_52),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_15),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_134),
.B1(n_136),
.B2(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_150),
.B(n_145),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_176),
.C(n_183),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_15),
.C(n_1),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_159),
.B(n_157),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_154),
.B1(n_168),
.B2(n_8),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_0),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_181),
.B(n_10),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_15),
.C(n_1),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_158),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_10),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_176),
.B(n_179),
.Y(n_203)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_172),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_15),
.C(n_7),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_194),
.C(n_196),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_182),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_2),
.C(n_3),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_201),
.B(n_196),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_204),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_182),
.B1(n_184),
.B2(n_178),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_206),
.C(n_190),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_180),
.B(n_183),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_194),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_203),
.B(n_205),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_170),
.Y(n_204)
);

AOI221xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_7),
.B1(n_10),
.B2(n_9),
.C(n_8),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_11),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_211),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_4),
.B(n_5),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_187),
.C(n_11),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_2),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_187),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_214),
.B(n_11),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_208),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_216),
.A2(n_221),
.B(n_5),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_5),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_4),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_4),
.Y(n_221)
);

AO21x2_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_224),
.B(n_5),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_223),
.A2(n_220),
.B(n_6),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_227),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_225),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_6),
.Y(n_231)
);


endmodule