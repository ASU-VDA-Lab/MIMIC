module fake_netlist_1_5655_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
AND2x2_ASAP7_75t_SL g10 ( .A(n_0), .B(n_5), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_10), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_12), .B(n_3), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_11), .B(n_4), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_10), .B1(n_13), .B2(n_14), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_17), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_13), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_15), .Y(n_26) );
NOR2x1_ASAP7_75t_SL g27 ( .A(n_26), .B(n_23), .Y(n_27) );
XNOR2xp5_ASAP7_75t_L g28 ( .A(n_25), .B(n_23), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OR5x1_ASAP7_75t_L g32 ( .A(n_30), .B(n_27), .C(n_6), .D(n_7), .E(n_8), .Y(n_32) );
AND3x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_9), .C(n_32), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
endmodule