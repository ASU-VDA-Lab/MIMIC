module fake_netlist_6_568_n_2299 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_356, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2299);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_356;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2299;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2291;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_2273;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_2069;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_2292;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_2016;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_2263;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_2298;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_652;
wire n_2154;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_2233;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2116;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_131),
.Y(n_569)
);

BUFx2_ASAP7_75t_SL g570 ( 
.A(n_400),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_68),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_119),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_24),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_255),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_377),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_159),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_522),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_6),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_21),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_59),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_322),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_186),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_216),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_349),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_145),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_311),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_195),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_271),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_220),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_22),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_250),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_385),
.Y(n_592)
);

CKINVDCx16_ASAP7_75t_R g593 ( 
.A(n_540),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_194),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_112),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_447),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_294),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_478),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_314),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_205),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_289),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_181),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_329),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_77),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_382),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_550),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_551),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_328),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g609 ( 
.A(n_320),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_346),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_452),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_75),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_312),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_184),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_78),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_538),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_496),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_473),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_418),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_38),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_45),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_271),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_37),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_318),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_439),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_520),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_159),
.Y(n_627)
);

BUFx10_ASAP7_75t_L g628 ( 
.A(n_167),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_388),
.Y(n_629)
);

CKINVDCx14_ASAP7_75t_R g630 ( 
.A(n_352),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_83),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_106),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_98),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_412),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_286),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_183),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_280),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_468),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_297),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_104),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_555),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_48),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_399),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_230),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_289),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_68),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_421),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_558),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_484),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_10),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_141),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_235),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_434),
.Y(n_653)
);

BUFx5_ASAP7_75t_L g654 ( 
.A(n_229),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_267),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_506),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_326),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_324),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_174),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_486),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_343),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_160),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_288),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_60),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_476),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_161),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_160),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_93),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_189),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_374),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_278),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_190),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_200),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_125),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_480),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_236),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_285),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_459),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_387),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_256),
.Y(n_680)
);

CKINVDCx16_ASAP7_75t_R g681 ( 
.A(n_269),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_509),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_72),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_157),
.Y(n_684)
);

CKINVDCx14_ASAP7_75t_R g685 ( 
.A(n_141),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_158),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_497),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_152),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_544),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_528),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_256),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_149),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_279),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_72),
.Y(n_694)
);

CKINVDCx14_ASAP7_75t_R g695 ( 
.A(n_110),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_375),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_241),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_446),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_337),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_292),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_32),
.Y(n_701)
);

CKINVDCx16_ASAP7_75t_R g702 ( 
.A(n_389),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_67),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_243),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_211),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_524),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_138),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_410),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_179),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_21),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_504),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_384),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_435),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_239),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_117),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_373),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_521),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_97),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_48),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_477),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_406),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_85),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_455),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_149),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_411),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_365),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_130),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_197),
.Y(n_728)
);

CKINVDCx16_ASAP7_75t_R g729 ( 
.A(n_121),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_227),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_293),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_233),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_284),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_268),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_443),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_111),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_533),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_316),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_567),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_325),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_440),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_50),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_56),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_286),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_241),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_531),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_144),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_264),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_394),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_417),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_305),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_395),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_327),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_183),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_519),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_129),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_330),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_157),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_431),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_396),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_39),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_565),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_371),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_517),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_86),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_4),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_39),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_76),
.Y(n_768)
);

CKINVDCx16_ASAP7_75t_R g769 ( 
.A(n_208),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_265),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_465),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_97),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_83),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_398),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_99),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_466),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_292),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_403),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_166),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_222),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_363),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_585),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_654),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_654),
.Y(n_784)
);

INVxp33_ASAP7_75t_SL g785 ( 
.A(n_730),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_654),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_654),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_585),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_654),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_654),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_685),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_654),
.Y(n_792)
);

CKINVDCx16_ASAP7_75t_R g793 ( 
.A(n_681),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_685),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_601),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_601),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_733),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_695),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_733),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_594),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_729),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_695),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_603),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_586),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_733),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_733),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_573),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_706),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_735),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_582),
.Y(n_810)
);

CKINVDCx14_ASAP7_75t_R g811 ( 
.A(n_630),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_571),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_769),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_589),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_569),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_602),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_612),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_593),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_579),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_572),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_574),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_571),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_594),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_613),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_643),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_620),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_623),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_635),
.Y(n_828)
);

INVxp33_ASAP7_75t_SL g829 ( 
.A(n_579),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_580),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_636),
.Y(n_831)
);

INVxp33_ASAP7_75t_L g832 ( 
.A(n_637),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_645),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_696),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_646),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_650),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_641),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_651),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_576),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_652),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_719),
.Y(n_841)
);

INVxp33_ASAP7_75t_SL g842 ( 
.A(n_580),
.Y(n_842)
);

INVxp33_ASAP7_75t_L g843 ( 
.A(n_662),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_578),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_664),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_671),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_673),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_583),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_719),
.Y(n_849)
);

INVxp33_ASAP7_75t_L g850 ( 
.A(n_677),
.Y(n_850)
);

INVxp33_ASAP7_75t_L g851 ( 
.A(n_680),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_683),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_583),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_686),
.Y(n_854)
);

INVxp33_ASAP7_75t_L g855 ( 
.A(n_688),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_691),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_587),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_625),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_692),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_693),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_701),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_703),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_709),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_595),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_586),
.Y(n_865)
);

INVxp33_ASAP7_75t_SL g866 ( 
.A(n_590),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_718),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_732),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_742),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_743),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_747),
.Y(n_871)
);

BUFx10_ASAP7_75t_L g872 ( 
.A(n_597),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_600),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_590),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_758),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_604),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_761),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_586),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_765),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_591),
.Y(n_880)
);

OAI21x1_ASAP7_75t_L g881 ( 
.A1(n_783),
.A2(n_771),
.B(n_619),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_806),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_825),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_825),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_806),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_825),
.Y(n_886)
);

OA21x2_ASAP7_75t_L g887 ( 
.A1(n_784),
.A2(n_619),
.B(n_592),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_825),
.Y(n_888)
);

OAI22x1_ASAP7_75t_SL g889 ( 
.A1(n_782),
.A2(n_591),
.B1(n_773),
.B2(n_772),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_783),
.B(n_641),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_797),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_792),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_825),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_792),
.B(n_771),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_786),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_799),
.B(n_771),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_837),
.B(n_630),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_787),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_805),
.B(n_581),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_815),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_834),
.B(n_609),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_789),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_790),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_795),
.B(n_702),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_812),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_812),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_822),
.B(n_592),
.Y(n_907)
);

AO22x1_ASAP7_75t_L g908 ( 
.A1(n_803),
.A2(n_773),
.B1(n_775),
.B2(n_772),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_822),
.A2(n_740),
.B(n_647),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_848),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_848),
.Y(n_911)
);

BUFx8_ASAP7_75t_L g912 ( 
.A(n_796),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_853),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_801),
.Y(n_914)
);

OA21x2_ASAP7_75t_L g915 ( 
.A1(n_853),
.A2(n_614),
.B(n_587),
.Y(n_915)
);

OA21x2_ASAP7_75t_L g916 ( 
.A1(n_857),
.A2(n_740),
.B(n_647),
.Y(n_916)
);

NOR2x1_ASAP7_75t_L g917 ( 
.A(n_857),
.B(n_570),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_807),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_811),
.B(n_779),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_810),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_791),
.B(n_607),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_791),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_SL g923 ( 
.A(n_794),
.B(n_625),
.Y(n_923)
);

INVx6_ASAP7_75t_L g924 ( 
.A(n_872),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_814),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_872),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_816),
.Y(n_927)
);

AND2x2_ASAP7_75t_SL g928 ( 
.A(n_818),
.B(n_643),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_817),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_824),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_826),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_827),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_828),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_831),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_833),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_815),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_835),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_836),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_838),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_840),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_845),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_846),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_884),
.Y(n_943)
);

BUFx10_ASAP7_75t_L g944 ( 
.A(n_921),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_900),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_904),
.B(n_793),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_R g947 ( 
.A(n_936),
.B(n_820),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_927),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_914),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_922),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_922),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_928),
.B(n_794),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_883),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_924),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_927),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_927),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_R g957 ( 
.A(n_923),
.B(n_820),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_890),
.Y(n_958)
);

AND3x2_ASAP7_75t_L g959 ( 
.A(n_923),
.B(n_653),
.C(n_614),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_R g960 ( 
.A(n_924),
.B(n_821),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_928),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_931),
.Y(n_962)
);

INVx5_ASAP7_75t_L g963 ( 
.A(n_884),
.Y(n_963)
);

INVx5_ASAP7_75t_L g964 ( 
.A(n_884),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_924),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_931),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_924),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_897),
.B(n_798),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_883),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_924),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_897),
.B(n_829),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_932),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_932),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_912),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_901),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_R g976 ( 
.A(n_926),
.B(n_821),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_934),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_928),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_926),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_926),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_912),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_926),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_926),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_926),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_890),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_926),
.B(n_839),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_883),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_904),
.B(n_829),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_912),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_919),
.B(n_839),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_934),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_912),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_889),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_R g994 ( 
.A(n_919),
.B(n_844),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_889),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_908),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_908),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_918),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_918),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_918),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_935),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_918),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_941),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_941),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_890),
.B(n_798),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_895),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_SL g1007 ( 
.A(n_899),
.Y(n_1007)
);

NOR2xp67_ASAP7_75t_L g1008 ( 
.A(n_938),
.B(n_873),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_883),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_918),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_895),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_R g1012 ( 
.A(n_938),
.B(n_844),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_918),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_933),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_R g1015 ( 
.A(n_938),
.B(n_864),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_R g1016 ( 
.A(n_915),
.B(n_785),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_895),
.Y(n_1017)
);

NOR2xp67_ASAP7_75t_L g1018 ( 
.A(n_938),
.B(n_873),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_933),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_884),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_R g1021 ( 
.A(n_915),
.B(n_785),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_933),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_933),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_933),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_884),
.Y(n_1025)
);

INVx5_ASAP7_75t_L g1026 ( 
.A(n_1020),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_988),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_988),
.B(n_842),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_967),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_958),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_985),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_971),
.B(n_842),
.Y(n_1032)
);

AND2x6_ASAP7_75t_L g1033 ( 
.A(n_971),
.B(n_596),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_962),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_954),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_975),
.B(n_813),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1006),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_966),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_945),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1011),
.B(n_902),
.Y(n_1040)
);

AND2x6_ASAP7_75t_L g1041 ( 
.A(n_948),
.B(n_606),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_968),
.B(n_866),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_944),
.B(n_866),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_944),
.B(n_864),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1017),
.B(n_902),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_960),
.B(n_802),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_972),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_1016),
.Y(n_1048)
);

BUFx8_ASAP7_75t_SL g1049 ( 
.A(n_949),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_965),
.Y(n_1050)
);

INVx6_ASAP7_75t_L g1051 ( 
.A(n_1020),
.Y(n_1051)
);

AND2x2_ASAP7_75t_SL g1052 ( 
.A(n_961),
.B(n_819),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_973),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_977),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_991),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_952),
.B(n_876),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_946),
.B(n_876),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_1001),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_998),
.B(n_902),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_955),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_956),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_978),
.B(n_802),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_970),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_953),
.Y(n_1064)
);

INVx4_ASAP7_75t_SL g1065 ( 
.A(n_1007),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_990),
.B(n_808),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_969),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_987),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_1020),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_1009),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1016),
.A2(n_738),
.B1(n_890),
.B2(n_917),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1012),
.B(n_872),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1020),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1008),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_994),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1015),
.B(n_809),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1025),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_1025),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1018),
.Y(n_1079)
);

BUFx10_ASAP7_75t_L g1080 ( 
.A(n_950),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1003),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1025),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_957),
.B(n_830),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1005),
.B(n_996),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_1004),
.Y(n_1085)
);

NAND3xp33_ASAP7_75t_L g1086 ( 
.A(n_1021),
.B(n_880),
.C(n_874),
.Y(n_1086)
);

AND2x6_ASAP7_75t_L g1087 ( 
.A(n_1025),
.B(n_608),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_951),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_999),
.B(n_903),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1000),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1007),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_1021),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_959),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1002),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1010),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_976),
.B(n_738),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_947),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_947),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_974),
.B(n_804),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_989),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_997),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_986),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1013),
.B(n_903),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_1014),
.Y(n_1104)
);

OAI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_992),
.A2(n_666),
.B1(n_676),
.B2(n_655),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_981),
.Y(n_1106)
);

NAND2xp33_ASAP7_75t_L g1107 ( 
.A(n_1019),
.B(n_577),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1022),
.B(n_847),
.Y(n_1108)
);

CKINVDCx16_ASAP7_75t_R g1109 ( 
.A(n_993),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1023),
.B(n_584),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_995),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_1024),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_979),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_943),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_943),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_943),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_943),
.B(n_852),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_963),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_963),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_963),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_980),
.B(n_865),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_982),
.B(n_903),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_963),
.Y(n_1123)
);

AND2x6_ASAP7_75t_L g1124 ( 
.A(n_983),
.B(n_611),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_984),
.B(n_878),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_964),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_964),
.Y(n_1127)
);

BUFx4f_ASAP7_75t_L g1128 ( 
.A(n_964),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_964),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_971),
.B(n_887),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_958),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_958),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_958),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_958),
.B(n_854),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_975),
.B(n_858),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_949),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_971),
.B(n_887),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_949),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_958),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_971),
.B(n_617),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_988),
.B(n_665),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_958),
.B(n_856),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_958),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_958),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_971),
.B(n_887),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_954),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_988),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_958),
.Y(n_1148)
);

INVxp33_ASAP7_75t_L g1149 ( 
.A(n_947),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_945),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_949),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_958),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_988),
.B(n_917),
.C(n_899),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_958),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_958),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_971),
.A2(n_915),
.B1(n_887),
.B2(n_916),
.Y(n_1156)
);

AND2x6_ASAP7_75t_L g1157 ( 
.A(n_971),
.B(n_618),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_958),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1141),
.B(n_933),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1141),
.B(n_894),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1027),
.B(n_894),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_1076),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_L g1163 ( 
.A(n_1033),
.B(n_598),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1027),
.B(n_894),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1059),
.A2(n_916),
.B(n_892),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1147),
.B(n_899),
.Y(n_1166)
);

NOR3xp33_ASAP7_75t_L g1167 ( 
.A(n_1028),
.B(n_762),
.C(n_725),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1034),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1147),
.B(n_899),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1028),
.B(n_1032),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_1058),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1092),
.A2(n_915),
.B1(n_744),
.B2(n_779),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1054),
.B(n_907),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1093),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1054),
.B(n_907),
.Y(n_1175)
);

AND2x6_ASAP7_75t_SL g1176 ( 
.A(n_1099),
.B(n_767),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1038),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1112),
.B(n_858),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1032),
.B(n_832),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1066),
.B(n_584),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1048),
.B(n_907),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1092),
.A2(n_915),
.B1(n_744),
.B2(n_704),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1048),
.B(n_843),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1083),
.B(n_782),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1047),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1136),
.B(n_850),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1042),
.A2(n_881),
.B(n_638),
.C(n_661),
.Y(n_1187)
);

OAI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1056),
.A2(n_668),
.B1(n_684),
.B2(n_642),
.C(n_588),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1090),
.B(n_690),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1033),
.A2(n_896),
.B1(n_682),
.B2(n_689),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1085),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1049),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1059),
.B(n_907),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1130),
.A2(n_629),
.B(n_713),
.C(n_712),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1055),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1053),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1089),
.B(n_898),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1089),
.B(n_898),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1094),
.B(n_690),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_1088),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1060),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1103),
.B(n_898),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1033),
.A2(n_704),
.B1(n_780),
.B2(n_770),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1136),
.B(n_788),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1086),
.B(n_851),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1061),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1138),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1030),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1149),
.B(n_1057),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1103),
.B(n_898),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1095),
.B(n_898),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1130),
.B(n_898),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1081),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1080),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_L g1215 ( 
.A(n_1029),
.B(n_859),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1137),
.B(n_716),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1104),
.B(n_776),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1134),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1137),
.B(n_726),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1151),
.B(n_788),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1145),
.A2(n_916),
.B(n_892),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1134),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_L g1223 ( 
.A(n_1033),
.B(n_599),
.Y(n_1223)
);

NOR2xp67_ASAP7_75t_L g1224 ( 
.A(n_1029),
.B(n_860),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1140),
.A2(n_896),
.B1(n_757),
.B2(n_760),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1080),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1140),
.A2(n_896),
.B1(n_774),
.B2(n_746),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1145),
.B(n_882),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1142),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1104),
.B(n_776),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1108),
.B(n_781),
.Y(n_1231)
);

NOR3xp33_ASAP7_75t_L g1232 ( 
.A(n_1062),
.B(n_781),
.C(n_861),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1140),
.A2(n_916),
.B1(n_881),
.B2(n_909),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1030),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1108),
.B(n_882),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1073),
.Y(n_1236)
);

NAND3xp33_ASAP7_75t_L g1237 ( 
.A(n_1036),
.B(n_823),
.C(n_800),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1142),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1151),
.B(n_855),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1140),
.A2(n_605),
.B1(n_616),
.B2(n_610),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1074),
.B(n_885),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1079),
.B(n_885),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1121),
.B(n_800),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1071),
.B(n_624),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1140),
.B(n_892),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1157),
.B(n_905),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1157),
.B(n_905),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1157),
.B(n_906),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1077),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1052),
.B(n_626),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1035),
.B(n_1050),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1097),
.B(n_823),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1097),
.B(n_841),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1157),
.B(n_1153),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1084),
.B(n_841),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1125),
.B(n_849),
.Y(n_1256)
);

AO22x1_ASAP7_75t_L g1257 ( 
.A1(n_1157),
.A2(n_775),
.B1(n_615),
.B2(n_622),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1031),
.B(n_906),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1101),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1131),
.B(n_910),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1037),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1101),
.A2(n_849),
.B1(n_621),
.B2(n_631),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1068),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1154),
.B(n_910),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1043),
.B(n_1044),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1096),
.B(n_627),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1063),
.B(n_634),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1132),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1155),
.B(n_913),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_SL g1270 ( 
.A(n_1111),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1156),
.B(n_920),
.Y(n_1271)
);

XNOR2x2_ASAP7_75t_L g1272 ( 
.A(n_1135),
.B(n_628),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1063),
.B(n_1075),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1039),
.B(n_920),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1070),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1133),
.B(n_632),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1146),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1139),
.B(n_920),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1070),
.Y(n_1279)
);

BUFx8_ASAP7_75t_L g1280 ( 
.A(n_1106),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1143),
.B(n_925),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1064),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1150),
.B(n_925),
.Y(n_1283)
);

OR2x6_ASAP7_75t_L g1284 ( 
.A(n_1099),
.B(n_862),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1144),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1158),
.A2(n_649),
.B1(n_656),
.B2(n_648),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1148),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1152),
.B(n_1122),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1067),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1072),
.B(n_633),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1098),
.B(n_639),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1122),
.B(n_925),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1113),
.B(n_657),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1040),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1102),
.B(n_929),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1040),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1102),
.B(n_929),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1046),
.B(n_863),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1110),
.B(n_929),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1045),
.B(n_1117),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1045),
.A2(n_937),
.B(n_939),
.C(n_930),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1117),
.B(n_930),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1107),
.B(n_930),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1069),
.B(n_658),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1082),
.B(n_937),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1078),
.B(n_937),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_1091),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1078),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1051),
.Y(n_1309)
);

NAND2xp33_ASAP7_75t_SL g1310 ( 
.A(n_1100),
.B(n_660),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1051),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1109),
.A2(n_736),
.B1(n_751),
.B2(n_667),
.Y(n_1312)
);

NOR2xp67_ASAP7_75t_SL g1313 ( 
.A(n_1026),
.B(n_643),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1041),
.A2(n_881),
.B1(n_909),
.B2(n_687),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1069),
.B(n_939),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1051),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1069),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1041),
.B(n_939),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1041),
.B(n_940),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1065),
.B(n_940),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_SL g1321 ( 
.A(n_1099),
.B(n_575),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1026),
.B(n_670),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1041),
.B(n_1124),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1115),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1041),
.B(n_940),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1116),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_SL g1327 ( 
.A(n_1105),
.B(n_575),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1126),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1026),
.B(n_675),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1026),
.B(n_678),
.Y(n_1330)
);

NOR2xp67_ASAP7_75t_L g1331 ( 
.A(n_1114),
.B(n_867),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1065),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1065),
.B(n_1105),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1118),
.B(n_640),
.Y(n_1334)
);

NOR2xp67_ASAP7_75t_L g1335 ( 
.A(n_1119),
.B(n_868),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1124),
.B(n_942),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1128),
.B(n_679),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1124),
.B(n_942),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1123),
.Y(n_1339)
);

AOI222xp33_ASAP7_75t_L g1340 ( 
.A1(n_1124),
.A2(n_628),
.B1(n_707),
.B2(n_705),
.C1(n_870),
.C2(n_869),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1127),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1124),
.B(n_1120),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1129),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1120),
.B(n_942),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1087),
.B(n_891),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1087),
.B(n_698),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1087),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1087),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1087),
.B(n_644),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1141),
.B(n_891),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1112),
.B(n_699),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1047),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1170),
.B(n_708),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1170),
.B(n_711),
.Y(n_1354)
);

CKINVDCx10_ASAP7_75t_R g1355 ( 
.A(n_1270),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1212),
.A2(n_909),
.B(n_888),
.Y(n_1356)
);

NOR3xp33_ASAP7_75t_L g1357 ( 
.A(n_1265),
.B(n_875),
.C(n_871),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1172),
.A2(n_888),
.B(n_884),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1172),
.A2(n_893),
.B(n_888),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1343),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_L g1361 ( 
.A1(n_1159),
.A2(n_877),
.B(n_879),
.C(n_886),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1162),
.A2(n_720),
.B1(n_721),
.B2(n_717),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1271),
.A2(n_886),
.B(n_778),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1182),
.A2(n_893),
.B(n_888),
.Y(n_1364)
);

NOR3xp33_ASAP7_75t_L g1365 ( 
.A(n_1179),
.B(n_663),
.C(n_659),
.Y(n_1365)
);

O2A1O1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1179),
.A2(n_886),
.B(n_575),
.C(n_705),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1165),
.A2(n_886),
.B(n_739),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1201),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1191),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1197),
.A2(n_893),
.B(n_888),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1167),
.A2(n_749),
.B1(n_750),
.B2(n_737),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1168),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1167),
.A2(n_753),
.B(n_755),
.C(n_752),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1209),
.B(n_1162),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1204),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1220),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1198),
.A2(n_1210),
.B(n_1202),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1209),
.B(n_669),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1255),
.B(n_672),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1266),
.A2(n_763),
.B(n_764),
.C(n_759),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1255),
.B(n_1183),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1165),
.A2(n_694),
.B(n_674),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1193),
.A2(n_893),
.B(n_911),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1300),
.A2(n_893),
.B(n_911),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1183),
.B(n_697),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1274),
.B(n_628),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1252),
.B(n_700),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1173),
.A2(n_911),
.B(n_687),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1175),
.A2(n_1221),
.B(n_1254),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1252),
.B(n_710),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1208),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1350),
.B(n_714),
.Y(n_1392)
);

AO21x1_ASAP7_75t_L g1393 ( 
.A1(n_1194),
.A2(n_687),
.B(n_643),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1177),
.Y(n_1394)
);

AND2x2_ASAP7_75t_SL g1395 ( 
.A(n_1327),
.B(n_723),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1288),
.B(n_715),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1343),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1195),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1283),
.B(n_722),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1259),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1206),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1294),
.B(n_724),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1258),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1221),
.A2(n_911),
.B(n_741),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1260),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1243),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1296),
.B(n_727),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1161),
.B(n_728),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1164),
.B(n_731),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1238),
.B(n_734),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1228),
.A2(n_911),
.B(n_741),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1270),
.B(n_705),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1216),
.A2(n_748),
.B(n_745),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1343),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1238),
.B(n_313),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1160),
.A2(n_911),
.B(n_741),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1282),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1332),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1188),
.A2(n_707),
.B(n_756),
.C(n_754),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1256),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1289),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1219),
.A2(n_768),
.B(n_766),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1166),
.B(n_1169),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1253),
.B(n_777),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1181),
.A2(n_741),
.B(n_723),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1292),
.B(n_723),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1264),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1269),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1174),
.Y(n_1429)
);

NOR2xp67_ASAP7_75t_L g1430 ( 
.A(n_1186),
.B(n_315),
.Y(n_1430)
);

AOI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1211),
.A2(n_723),
.B(n_319),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1184),
.B(n_1239),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1207),
.B(n_707),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1208),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1342),
.A2(n_321),
.B(n_317),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1245),
.A2(n_331),
.B(n_323),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1303),
.A2(n_333),
.B(n_332),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1295),
.B(n_0),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1277),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1297),
.B(n_0),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1174),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1232),
.B(n_334),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1232),
.B(n_335),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1205),
.B(n_1352),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1205),
.B(n_1),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1233),
.A2(n_338),
.B(n_336),
.Y(n_1446)
);

OAI21xp33_ASAP7_75t_L g1447 ( 
.A1(n_1253),
.A2(n_1),
.B(n_2),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1203),
.A2(n_340),
.B1(n_341),
.B2(n_339),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1233),
.A2(n_344),
.B(n_342),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1185),
.B(n_2),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1246),
.A2(n_347),
.B(n_345),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1187),
.A2(n_568),
.B(n_350),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1291),
.B(n_1180),
.Y(n_1453)
);

NOR3xp33_ASAP7_75t_L g1454 ( 
.A(n_1237),
.B(n_3),
.C(n_4),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1215),
.B(n_348),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1196),
.B(n_3),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1287),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1218),
.B(n_351),
.Y(n_1458)
);

AO21x1_ASAP7_75t_L g1459 ( 
.A1(n_1194),
.A2(n_5),
.B(n_6),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1247),
.A2(n_354),
.B(n_353),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1263),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1248),
.A2(n_356),
.B(n_355),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1275),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1290),
.A2(n_8),
.B(n_5),
.C(n_7),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1235),
.B(n_7),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1234),
.B(n_8),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1250),
.A2(n_1244),
.B(n_1333),
.C(n_1199),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1314),
.A2(n_358),
.B(n_357),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1314),
.A2(n_566),
.B(n_360),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1290),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1301),
.A2(n_361),
.B(n_359),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1302),
.A2(n_364),
.B(n_362),
.Y(n_1472)
);

NOR3xp33_ASAP7_75t_L g1473 ( 
.A(n_1178),
.B(n_9),
.C(n_11),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1163),
.A2(n_367),
.B(n_366),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1279),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1340),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1224),
.B(n_368),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1213),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1223),
.A2(n_370),
.B(n_369),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1261),
.B(n_12),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1299),
.B(n_13),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1278),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1222),
.B(n_372),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1301),
.A2(n_378),
.B(n_376),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1203),
.A2(n_1338),
.B(n_1336),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1229),
.B(n_14),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1236),
.Y(n_1487)
);

AND2x2_ASAP7_75t_SL g1488 ( 
.A(n_1321),
.B(n_15),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1323),
.A2(n_1344),
.B(n_1306),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1281),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1189),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_R g1492 ( 
.A(n_1310),
.B(n_379),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1320),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1298),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1276),
.B(n_16),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1276),
.B(n_1241),
.Y(n_1496)
);

NOR3xp33_ASAP7_75t_L g1497 ( 
.A(n_1312),
.B(n_17),
.C(n_18),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1242),
.B(n_18),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1334),
.B(n_19),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1334),
.B(n_19),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1200),
.B(n_1268),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1285),
.B(n_20),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1339),
.B(n_20),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1341),
.B(n_22),
.Y(n_1504)
);

NOR2xp67_ASAP7_75t_L g1505 ( 
.A(n_1214),
.B(n_380),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1315),
.A2(n_383),
.B(n_381),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1171),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1251),
.B(n_386),
.Y(n_1508)
);

INVxp67_ASAP7_75t_L g1509 ( 
.A(n_1231),
.Y(n_1509)
);

NOR2xp67_ASAP7_75t_L g1510 ( 
.A(n_1226),
.B(n_390),
.Y(n_1510)
);

AO21x1_ASAP7_75t_L g1511 ( 
.A1(n_1318),
.A2(n_23),
.B(n_24),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1257),
.B(n_23),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1319),
.A2(n_392),
.B(n_391),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1307),
.B(n_25),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1325),
.A2(n_397),
.B(n_393),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1251),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1262),
.B(n_25),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1305),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1304),
.A2(n_402),
.B(n_401),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1308),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1331),
.B(n_26),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1335),
.B(n_1349),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1347),
.A2(n_405),
.B(n_404),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1317),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1249),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1324),
.B(n_26),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1307),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1322),
.A2(n_408),
.B(n_407),
.Y(n_1528)
);

NOR3xp33_ASAP7_75t_L g1529 ( 
.A(n_1351),
.B(n_27),
.C(n_28),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1329),
.A2(n_413),
.B(n_409),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1190),
.A2(n_415),
.B(n_414),
.Y(n_1531)
);

O2A1O1Ixp5_ASAP7_75t_L g1532 ( 
.A1(n_1346),
.A2(n_419),
.B(n_420),
.C(n_416),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1286),
.B(n_422),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1330),
.A2(n_424),
.B(n_423),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1324),
.B(n_29),
.Y(n_1535)
);

AOI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1348),
.A2(n_426),
.B(n_425),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1326),
.B(n_30),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1337),
.A2(n_428),
.B(n_427),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1262),
.B(n_429),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1251),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1328),
.A2(n_432),
.B(n_430),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1309),
.A2(n_436),
.B(n_433),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1311),
.A2(n_438),
.B(n_437),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1284),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1316),
.B(n_30),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1192),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1249),
.A2(n_442),
.B(n_441),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1273),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1345),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1225),
.A2(n_445),
.B1(n_448),
.B2(n_444),
.Y(n_1550)
);

AO21x2_ASAP7_75t_L g1551 ( 
.A1(n_1425),
.A2(n_1227),
.B(n_1240),
.Y(n_1551)
);

NOR2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1546),
.B(n_1272),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1377),
.A2(n_1267),
.B(n_1230),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1372),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1461),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1406),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1381),
.B(n_1217),
.Y(n_1557)
);

BUFx4f_ASAP7_75t_SL g1558 ( 
.A(n_1360),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1394),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1369),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1522),
.A2(n_1293),
.B(n_1313),
.Y(n_1561)
);

BUFx12f_ASAP7_75t_L g1562 ( 
.A(n_1439),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1379),
.B(n_1284),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1389),
.A2(n_1284),
.B(n_450),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1375),
.B(n_1280),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1398),
.Y(n_1566)
);

NAND3xp33_ASAP7_75t_SL g1567 ( 
.A(n_1497),
.B(n_1176),
.C(n_1280),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_1429),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1360),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1453),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1496),
.A2(n_34),
.B1(n_31),
.B2(n_33),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1420),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1374),
.B(n_34),
.Y(n_1573)
);

AO21x1_ASAP7_75t_L g1574 ( 
.A1(n_1469),
.A2(n_35),
.B(n_36),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1423),
.A2(n_451),
.B(n_449),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1355),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1378),
.B(n_35),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1467),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1432),
.B(n_40),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1392),
.B(n_40),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1495),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1376),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1360),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1395),
.B(n_41),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1400),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1489),
.A2(n_454),
.B(n_453),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1414),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1478),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_L g1589 ( 
.A(n_1387),
.B(n_42),
.C(n_43),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1353),
.B(n_44),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1354),
.B(n_44),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1485),
.A2(n_457),
.B(n_456),
.Y(n_1592)
);

A2O1A1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1469),
.A2(n_1500),
.B(n_1499),
.C(n_1424),
.Y(n_1593)
);

O2A1O1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1445),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1386),
.B(n_1494),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_SL g1596 ( 
.A1(n_1539),
.A2(n_1443),
.B(n_1442),
.C(n_1533),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1414),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1444),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1485),
.A2(n_460),
.B(n_458),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1390),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1426),
.A2(n_462),
.B(n_461),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1493),
.B(n_51),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1356),
.A2(n_464),
.B(n_463),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1414),
.Y(n_1604)
);

NOR3xp33_ASAP7_75t_L g1605 ( 
.A(n_1476),
.B(n_52),
.C(n_53),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1403),
.B(n_52),
.Y(n_1606)
);

AOI21xp33_ASAP7_75t_L g1607 ( 
.A1(n_1413),
.A2(n_53),
.B(n_54),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1397),
.B(n_467),
.Y(n_1608)
);

BUFx8_ASAP7_75t_L g1609 ( 
.A(n_1540),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1452),
.A2(n_470),
.B(n_469),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1405),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_R g1612 ( 
.A(n_1493),
.B(n_471),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1493),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1452),
.A2(n_474),
.B(n_472),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1427),
.B(n_55),
.Y(n_1615)
);

AO32x2_ASAP7_75t_L g1616 ( 
.A1(n_1448),
.A2(n_59),
.A3(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_1616)
);

OAI22x1_ASAP7_75t_L g1617 ( 
.A1(n_1517),
.A2(n_1509),
.B1(n_1516),
.B2(n_1508),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1428),
.B(n_61),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1368),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1365),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1385),
.B(n_1396),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1397),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1401),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1430),
.A2(n_1488),
.B1(n_1399),
.B2(n_1410),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1417),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1482),
.B(n_62),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1490),
.B(n_63),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1391),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1421),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1402),
.B(n_64),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1441),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1407),
.B(n_65),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1441),
.B(n_65),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1408),
.B(n_66),
.Y(n_1634)
);

O2A1O1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1464),
.A2(n_69),
.B(n_66),
.C(n_67),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1409),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1636)
);

INVx4_ASAP7_75t_L g1637 ( 
.A(n_1418),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1457),
.A2(n_73),
.B1(n_70),
.B2(n_71),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1463),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1468),
.A2(n_479),
.B(n_475),
.Y(n_1640)
);

OAI22x1_ASAP7_75t_L g1641 ( 
.A1(n_1516),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1475),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1357),
.B(n_74),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1487),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1438),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1548),
.B(n_1507),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1548),
.B(n_1501),
.Y(n_1647)
);

OAI21xp33_ASAP7_75t_SL g1648 ( 
.A1(n_1471),
.A2(n_79),
.B(n_80),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1415),
.B(n_79),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1391),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1433),
.B(n_1465),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1474),
.A2(n_482),
.B(n_481),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1440),
.B(n_80),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1544),
.B(n_81),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1434),
.A2(n_84),
.B1(n_81),
.B2(n_82),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1479),
.A2(n_485),
.B(n_483),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1447),
.A2(n_1419),
.B1(n_1473),
.B2(n_1454),
.C(n_1529),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1362),
.B(n_82),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_SL g1659 ( 
.A(n_1527),
.B(n_84),
.C(n_85),
.Y(n_1659)
);

AOI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1404),
.A2(n_488),
.B(n_487),
.Y(n_1660)
);

NAND2x1_ASAP7_75t_SL g1661 ( 
.A(n_1508),
.B(n_86),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1422),
.B(n_87),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1492),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1367),
.A2(n_490),
.B(n_489),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1415),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1498),
.B(n_87),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1514),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1412),
.B(n_88),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1518),
.B(n_88),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1418),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1531),
.A2(n_1366),
.B(n_1484),
.C(n_1471),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1367),
.A2(n_1449),
.B(n_1446),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1525),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1524),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1458),
.B(n_564),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1549),
.B(n_89),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1458),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1524),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1531),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1502),
.B(n_92),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1524),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1481),
.B(n_93),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1486),
.B(n_94),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1412),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1418),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1363),
.A2(n_492),
.B(n_491),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1470),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1483),
.B(n_95),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1450),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1483),
.B(n_563),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1371),
.B(n_96),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1503),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1480),
.B(n_98),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1434),
.B(n_99),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1466),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1520),
.B(n_100),
.Y(n_1696)
);

INVx4_ASAP7_75t_L g1697 ( 
.A(n_1505),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1456),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1373),
.B(n_101),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1512),
.A2(n_1491),
.B(n_1521),
.C(n_1484),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1504),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1545),
.B(n_102),
.Y(n_1702)
);

A2O1A1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1382),
.A2(n_106),
.B(n_103),
.C(n_105),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1380),
.A2(n_108),
.B(n_105),
.C(n_107),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1382),
.B(n_107),
.Y(n_1705)
);

BUFx8_ASAP7_75t_SL g1706 ( 
.A(n_1526),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1510),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1707)
);

O2A1O1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1537),
.A2(n_112),
.B(n_109),
.C(n_111),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1535),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1361),
.A2(n_494),
.B(n_493),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1532),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1523),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1511),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1358),
.A2(n_498),
.B(n_495),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1455),
.B(n_113),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1359),
.A2(n_500),
.B(n_499),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1431),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1459),
.B(n_1477),
.Y(n_1718)
);

O2A1O1Ixp5_ASAP7_75t_L g1719 ( 
.A1(n_1393),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1538),
.B(n_116),
.Y(n_1720)
);

AOI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1370),
.A2(n_562),
.B(n_502),
.Y(n_1721)
);

AND2x6_ASAP7_75t_L g1722 ( 
.A(n_1536),
.B(n_501),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_SL g1723 ( 
.A(n_1519),
.B(n_117),
.C(n_118),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1364),
.A2(n_1383),
.B(n_1435),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1550),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1384),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1416),
.B(n_120),
.Y(n_1727)
);

INVx4_ASAP7_75t_L g1728 ( 
.A(n_1528),
.Y(n_1728)
);

BUFx4f_ASAP7_75t_L g1729 ( 
.A(n_1530),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1411),
.B(n_121),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1593),
.A2(n_1472),
.B(n_1437),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1672),
.A2(n_1436),
.B(n_1451),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1554),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1559),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1671),
.A2(n_1534),
.B(n_1460),
.C(n_1462),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1724),
.A2(n_1515),
.B(n_1513),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1566),
.Y(n_1737)
);

OAI21x1_ASAP7_75t_L g1738 ( 
.A1(n_1726),
.A2(n_1547),
.B(n_1506),
.Y(n_1738)
);

AOI31xp67_ASAP7_75t_L g1739 ( 
.A1(n_1718),
.A2(n_1388),
.A3(n_1541),
.B(n_1543),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1700),
.A2(n_1577),
.B(n_1621),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1610),
.A2(n_1542),
.B(n_505),
.Y(n_1741)
);

NOR2x1_ASAP7_75t_L g1742 ( 
.A(n_1697),
.B(n_503),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1557),
.B(n_122),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1563),
.B(n_122),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1555),
.Y(n_1745)
);

BUFx6f_ASAP7_75t_L g1746 ( 
.A(n_1587),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1614),
.A2(n_1553),
.B(n_1729),
.Y(n_1747)
);

AOI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1607),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.C(n_126),
.Y(n_1748)
);

A2O1A1Ixp33_ASAP7_75t_L g1749 ( 
.A1(n_1651),
.A2(n_1666),
.B(n_1657),
.C(n_1662),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1729),
.A2(n_561),
.B(n_508),
.Y(n_1750)
);

OAI21x1_ASAP7_75t_L g1751 ( 
.A1(n_1603),
.A2(n_510),
.B(n_507),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1692),
.B(n_123),
.Y(n_1752)
);

OAI21x1_ASAP7_75t_L g1753 ( 
.A1(n_1660),
.A2(n_512),
.B(n_511),
.Y(n_1753)
);

AO31x2_ASAP7_75t_L g1754 ( 
.A1(n_1574),
.A2(n_127),
.A3(n_124),
.B(n_126),
.Y(n_1754)
);

AND2x6_ASAP7_75t_L g1755 ( 
.A(n_1675),
.B(n_513),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1596),
.A2(n_560),
.B(n_515),
.Y(n_1756)
);

AO22x2_ASAP7_75t_L g1757 ( 
.A1(n_1605),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1757)
);

OAI21x1_ASAP7_75t_SL g1758 ( 
.A1(n_1635),
.A2(n_128),
.B(n_130),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1689),
.B(n_131),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1587),
.Y(n_1760)
);

OAI21xp33_ASAP7_75t_L g1761 ( 
.A1(n_1683),
.A2(n_132),
.B(n_133),
.Y(n_1761)
);

AO31x2_ASAP7_75t_L g1762 ( 
.A1(n_1713),
.A2(n_1705),
.A3(n_1679),
.B(n_1686),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1564),
.A2(n_516),
.B(n_514),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1717),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1625),
.Y(n_1765)
);

BUFx10_ASAP7_75t_L g1766 ( 
.A(n_1576),
.Y(n_1766)
);

NAND3xp33_ASAP7_75t_L g1767 ( 
.A(n_1658),
.B(n_132),
.C(n_133),
.Y(n_1767)
);

OAI21x1_ASAP7_75t_L g1768 ( 
.A1(n_1721),
.A2(n_523),
.B(n_518),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1562),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1551),
.A2(n_526),
.B(n_525),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1579),
.B(n_134),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1698),
.B(n_1595),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1670),
.Y(n_1773)
);

OAI21x1_ASAP7_75t_L g1774 ( 
.A1(n_1586),
.A2(n_529),
.B(n_527),
.Y(n_1774)
);

OA21x2_ASAP7_75t_L g1775 ( 
.A1(n_1592),
.A2(n_532),
.B(n_530),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1551),
.A2(n_1561),
.B(n_1728),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1695),
.A2(n_134),
.B(n_135),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1619),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1623),
.Y(n_1779)
);

AO31x2_ASAP7_75t_L g1780 ( 
.A1(n_1711),
.A2(n_135),
.A3(n_136),
.B(n_137),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1556),
.B(n_534),
.Y(n_1781)
);

OAI21x1_ASAP7_75t_L g1782 ( 
.A1(n_1599),
.A2(n_536),
.B(n_535),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1709),
.B(n_136),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1590),
.A2(n_137),
.B(n_138),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1728),
.A2(n_539),
.B(n_537),
.Y(n_1785)
);

AOI21x1_ASAP7_75t_L g1786 ( 
.A1(n_1720),
.A2(n_542),
.B(n_541),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1624),
.B(n_139),
.Y(n_1787)
);

NAND2x1_ASAP7_75t_L g1788 ( 
.A(n_1628),
.B(n_543),
.Y(n_1788)
);

AOI211x1_ASAP7_75t_L g1789 ( 
.A1(n_1584),
.A2(n_139),
.B(n_140),
.C(n_142),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1591),
.A2(n_140),
.B(n_142),
.Y(n_1790)
);

AO31x2_ASAP7_75t_L g1791 ( 
.A1(n_1703),
.A2(n_143),
.A3(n_144),
.B(n_145),
.Y(n_1791)
);

INVxp67_ASAP7_75t_L g1792 ( 
.A(n_1560),
.Y(n_1792)
);

NOR2xp67_ASAP7_75t_L g1793 ( 
.A(n_1697),
.B(n_545),
.Y(n_1793)
);

OAI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1714),
.A2(n_547),
.B(n_546),
.Y(n_1794)
);

A2O1A1Ixp33_ASAP7_75t_L g1795 ( 
.A1(n_1648),
.A2(n_143),
.B(n_146),
.C(n_147),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1647),
.B(n_146),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1573),
.B(n_147),
.Y(n_1797)
);

OA21x2_ASAP7_75t_L g1798 ( 
.A1(n_1727),
.A2(n_549),
.B(n_548),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1639),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1640),
.A2(n_1575),
.B(n_1652),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1656),
.A2(n_553),
.B(n_552),
.Y(n_1801)
);

INVx1_ASAP7_75t_SL g1802 ( 
.A(n_1585),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1580),
.A2(n_148),
.B(n_150),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1664),
.A2(n_556),
.B(n_554),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1684),
.B(n_148),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1665),
.B(n_1631),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1578),
.A2(n_150),
.B(n_151),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_SL g1808 ( 
.A1(n_1675),
.A2(n_559),
.B(n_557),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1667),
.B(n_151),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1642),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_L g1811 ( 
.A(n_1663),
.B(n_152),
.Y(n_1811)
);

OAI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1716),
.A2(n_153),
.B(n_154),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1630),
.B(n_153),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1710),
.A2(n_154),
.B(n_155),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1617),
.B(n_155),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1572),
.A2(n_156),
.B1(n_158),
.B2(n_161),
.Y(n_1816)
);

OAI21x1_ASAP7_75t_L g1817 ( 
.A1(n_1710),
.A2(n_156),
.B(n_162),
.Y(n_1817)
);

OAI21x1_ASAP7_75t_L g1818 ( 
.A1(n_1601),
.A2(n_162),
.B(n_163),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1730),
.A2(n_163),
.B(n_164),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1632),
.B(n_164),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1664),
.A2(n_312),
.B(n_165),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1606),
.B(n_165),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1615),
.B(n_1618),
.Y(n_1823)
);

OA21x2_ASAP7_75t_L g1824 ( 
.A1(n_1719),
.A2(n_166),
.B(n_167),
.Y(n_1824)
);

AND2x2_ASAP7_75t_SL g1825 ( 
.A(n_1690),
.B(n_168),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1682),
.A2(n_169),
.B(n_170),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1690),
.B(n_170),
.Y(n_1827)
);

AOI21x1_ASAP7_75t_L g1828 ( 
.A1(n_1725),
.A2(n_171),
.B(n_172),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1628),
.A2(n_171),
.B(n_172),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1629),
.Y(n_1830)
);

AOI21xp33_ASAP7_75t_L g1831 ( 
.A1(n_1691),
.A2(n_173),
.B(n_174),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1650),
.A2(n_173),
.B(n_175),
.Y(n_1832)
);

OAI21x1_ASAP7_75t_L g1833 ( 
.A1(n_1650),
.A2(n_1699),
.B(n_1676),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1644),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1588),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1582),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1702),
.B(n_176),
.Y(n_1837)
);

OAI21x1_ASAP7_75t_L g1838 ( 
.A1(n_1704),
.A2(n_177),
.B(n_178),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_SL g1839 ( 
.A(n_1620),
.B(n_177),
.C(n_178),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1653),
.B(n_179),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1715),
.A2(n_1693),
.B(n_1589),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1687),
.A2(n_1608),
.B(n_1669),
.Y(n_1842)
);

AOI221x1_ASAP7_75t_L g1843 ( 
.A1(n_1600),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.C(n_184),
.Y(n_1843)
);

OAI21x1_ASAP7_75t_L g1844 ( 
.A1(n_1673),
.A2(n_180),
.B(n_182),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1649),
.B(n_185),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1712),
.A2(n_311),
.B(n_186),
.Y(n_1846)
);

O2A1O1Ixp5_ASAP7_75t_L g1847 ( 
.A1(n_1571),
.A2(n_1680),
.B(n_1645),
.C(n_1636),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1626),
.A2(n_310),
.B(n_187),
.Y(n_1848)
);

AO31x2_ASAP7_75t_L g1849 ( 
.A1(n_1598),
.A2(n_1701),
.A3(n_1694),
.B(n_1696),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1567),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1668),
.A2(n_188),
.B(n_189),
.C(n_190),
.Y(n_1851)
);

OAI22x1_ASAP7_75t_L g1852 ( 
.A1(n_1570),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1597),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1613),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1627),
.B(n_191),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1646),
.B(n_192),
.Y(n_1856)
);

NOR2xp67_ASAP7_75t_L g1857 ( 
.A(n_1565),
.B(n_193),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1609),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1568),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1616),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_SL g1861 ( 
.A1(n_1602),
.A2(n_194),
.B(n_195),
.C(n_196),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1678),
.A2(n_310),
.B(n_199),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1587),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1708),
.A2(n_198),
.B(n_199),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1613),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1643),
.B(n_198),
.Y(n_1866)
);

OAI21x1_ASAP7_75t_L g1867 ( 
.A1(n_1581),
.A2(n_200),
.B(n_201),
.Y(n_1867)
);

NOR2xp67_ASAP7_75t_SL g1868 ( 
.A(n_1634),
.B(n_201),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1688),
.B(n_202),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1613),
.B(n_202),
.Y(n_1870)
);

BUFx12f_ASAP7_75t_L g1871 ( 
.A(n_1609),
.Y(n_1871)
);

A2O1A1Ixp33_ASAP7_75t_L g1872 ( 
.A1(n_1723),
.A2(n_1594),
.B(n_1659),
.C(n_1677),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1558),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1706),
.B(n_203),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1633),
.Y(n_1875)
);

OAI21x1_ASAP7_75t_L g1876 ( 
.A1(n_1722),
.A2(n_204),
.B(n_205),
.Y(n_1876)
);

OAI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1722),
.A2(n_206),
.B(n_207),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1552),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1674),
.Y(n_1879)
);

AOI21x1_ASAP7_75t_SL g1880 ( 
.A1(n_1616),
.A2(n_206),
.B(n_207),
.Y(n_1880)
);

NOR2xp67_ASAP7_75t_SL g1881 ( 
.A(n_1622),
.B(n_208),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1681),
.A2(n_309),
.B(n_210),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1622),
.Y(n_1883)
);

OAI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1707),
.A2(n_1611),
.B(n_1655),
.Y(n_1884)
);

OAI21x1_ASAP7_75t_L g1885 ( 
.A1(n_1722),
.A2(n_209),
.B(n_210),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1661),
.B(n_209),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1854),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1733),
.Y(n_1888)
);

AO21x2_ASAP7_75t_L g1889 ( 
.A1(n_1776),
.A2(n_1612),
.B(n_1638),
.Y(n_1889)
);

OAI21x1_ASAP7_75t_L g1890 ( 
.A1(n_1747),
.A2(n_1722),
.B(n_1654),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1733),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1800),
.A2(n_1616),
.B(n_1641),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1732),
.A2(n_1622),
.B(n_1569),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1749),
.B(n_1583),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1823),
.B(n_1604),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1740),
.A2(n_1569),
.B(n_1637),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1734),
.Y(n_1897)
);

OAI21x1_ASAP7_75t_L g1898 ( 
.A1(n_1738),
.A2(n_1736),
.B(n_1753),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1731),
.A2(n_1637),
.B(n_1604),
.Y(n_1899)
);

AND2x2_ASAP7_75t_SL g1900 ( 
.A(n_1860),
.B(n_1825),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1772),
.B(n_1841),
.Y(n_1901)
);

OAI21x1_ASAP7_75t_L g1902 ( 
.A1(n_1768),
.A2(n_1604),
.B(n_1685),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1875),
.B(n_1685),
.Y(n_1903)
);

NOR2xp67_ASAP7_75t_L g1904 ( 
.A(n_1859),
.B(n_1685),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1735),
.A2(n_1741),
.B(n_1756),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1839),
.A2(n_1761),
.B1(n_1803),
.B2(n_1790),
.Y(n_1906)
);

OA21x2_ASAP7_75t_L g1907 ( 
.A1(n_1814),
.A2(n_211),
.B(n_212),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1737),
.Y(n_1908)
);

AOI21xp33_ASAP7_75t_L g1909 ( 
.A1(n_1847),
.A2(n_212),
.B(n_213),
.Y(n_1909)
);

CKINVDCx20_ASAP7_75t_R g1910 ( 
.A(n_1766),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1879),
.B(n_213),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1737),
.Y(n_1912)
);

NAND3xp33_ASAP7_75t_L g1913 ( 
.A(n_1784),
.B(n_214),
.C(n_215),
.Y(n_1913)
);

OAI21x1_ASAP7_75t_L g1914 ( 
.A1(n_1763),
.A2(n_214),
.B(n_215),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1836),
.Y(n_1915)
);

OA21x2_ASAP7_75t_L g1916 ( 
.A1(n_1817),
.A2(n_216),
.B(n_217),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1787),
.B(n_217),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1746),
.Y(n_1918)
);

OAI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1767),
.A2(n_1843),
.B1(n_1850),
.B2(n_1837),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1764),
.Y(n_1920)
);

OAI21x1_ASAP7_75t_L g1921 ( 
.A1(n_1770),
.A2(n_218),
.B(n_219),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1807),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.C(n_221),
.Y(n_1922)
);

OAI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1804),
.A2(n_221),
.B(n_222),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1854),
.B(n_223),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1873),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1766),
.Y(n_1926)
);

OAI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1774),
.A2(n_223),
.B(n_224),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1806),
.B(n_224),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1765),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1778),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1764),
.Y(n_1931)
);

O2A1O1Ixp5_ASAP7_75t_L g1932 ( 
.A1(n_1821),
.A2(n_225),
.B(n_226),
.C(n_227),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1773),
.Y(n_1933)
);

OAI21x1_ASAP7_75t_L g1934 ( 
.A1(n_1782),
.A2(n_225),
.B(n_226),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1778),
.Y(n_1935)
);

CKINVDCx11_ASAP7_75t_R g1936 ( 
.A(n_1871),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1779),
.Y(n_1937)
);

OAI21x1_ASAP7_75t_L g1938 ( 
.A1(n_1751),
.A2(n_1794),
.B(n_1812),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1769),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1865),
.B(n_228),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1826),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_1941)
);

OAI21x1_ASAP7_75t_L g1942 ( 
.A1(n_1833),
.A2(n_231),
.B(n_232),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1779),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_L g1944 ( 
.A1(n_1785),
.A2(n_231),
.B(n_232),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1883),
.B(n_233),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1799),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1810),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1757),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1834),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1872),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1757),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_1951)
);

AOI21xp33_ASAP7_75t_L g1952 ( 
.A1(n_1884),
.A2(n_240),
.B(n_242),
.Y(n_1952)
);

INVx1_ASAP7_75t_SL g1953 ( 
.A(n_1835),
.Y(n_1953)
);

O2A1O1Ixp33_ASAP7_75t_SL g1954 ( 
.A1(n_1795),
.A2(n_240),
.B(n_242),
.C(n_243),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1762),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1883),
.B(n_244),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1801),
.A2(n_244),
.B(n_245),
.Y(n_1957)
);

AOI21x1_ASAP7_75t_L g1958 ( 
.A1(n_1828),
.A2(n_245),
.B(n_246),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1743),
.B(n_309),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1745),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1750),
.A2(n_246),
.B(n_247),
.Y(n_1961)
);

O2A1O1Ixp33_ASAP7_75t_SL g1962 ( 
.A1(n_1777),
.A2(n_247),
.B(n_248),
.C(n_249),
.Y(n_1962)
);

OA21x2_ASAP7_75t_L g1963 ( 
.A1(n_1818),
.A2(n_248),
.B(n_249),
.Y(n_1963)
);

OAI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1842),
.A2(n_250),
.B(n_251),
.Y(n_1964)
);

NOR2xp67_ASAP7_75t_L g1965 ( 
.A(n_1792),
.B(n_251),
.Y(n_1965)
);

O2A1O1Ixp33_ASAP7_75t_SL g1966 ( 
.A1(n_1748),
.A2(n_252),
.B(n_253),
.C(n_254),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1866),
.B(n_1771),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1830),
.Y(n_1968)
);

OAI21x1_ASAP7_75t_L g1969 ( 
.A1(n_1786),
.A2(n_252),
.B(n_253),
.Y(n_1969)
);

INVx4_ASAP7_75t_L g1970 ( 
.A(n_1746),
.Y(n_1970)
);

OAI21x1_ASAP7_75t_L g1971 ( 
.A1(n_1775),
.A2(n_254),
.B(n_255),
.Y(n_1971)
);

BUFx4_ASAP7_75t_SL g1972 ( 
.A(n_1878),
.Y(n_1972)
);

OAI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1852),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1762),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1746),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1809),
.B(n_257),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1744),
.B(n_1856),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1802),
.B(n_308),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1798),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1853),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1838),
.A2(n_258),
.B(n_259),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1760),
.Y(n_1982)
);

OAI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1846),
.A2(n_260),
.B(n_261),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1754),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1762),
.Y(n_1985)
);

AOI21xp33_ASAP7_75t_L g1986 ( 
.A1(n_1797),
.A2(n_260),
.B(n_261),
.Y(n_1986)
);

OA21x2_ASAP7_75t_L g1987 ( 
.A1(n_1844),
.A2(n_262),
.B(n_263),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1796),
.B(n_262),
.Y(n_1988)
);

AO21x2_ASAP7_75t_L g1989 ( 
.A1(n_1905),
.A2(n_1758),
.B(n_1860),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1901),
.B(n_1977),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1955),
.B(n_1791),
.Y(n_1991)
);

OA21x2_ASAP7_75t_L g1992 ( 
.A1(n_1898),
.A2(n_1979),
.B(n_1892),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1946),
.B(n_1815),
.Y(n_1993)
);

OAI21x1_ASAP7_75t_SL g1994 ( 
.A1(n_1983),
.A2(n_1848),
.B(n_1862),
.Y(n_1994)
);

AO21x2_ASAP7_75t_L g1995 ( 
.A1(n_1979),
.A2(n_1984),
.B(n_1974),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1897),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1922),
.A2(n_1845),
.B(n_1831),
.C(n_1851),
.Y(n_1997)
);

OAI21x1_ASAP7_75t_L g1998 ( 
.A1(n_1938),
.A2(n_1832),
.B(n_1829),
.Y(n_1998)
);

OA21x2_ASAP7_75t_L g1999 ( 
.A1(n_1971),
.A2(n_1877),
.B(n_1885),
.Y(n_1999)
);

OAI21x1_ASAP7_75t_L g2000 ( 
.A1(n_1942),
.A2(n_1876),
.B(n_1775),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1920),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1906),
.A2(n_1868),
.B1(n_1755),
.B2(n_1857),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1893),
.A2(n_1808),
.B(n_1798),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1888),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1929),
.Y(n_2005)
);

AOI21x1_ASAP7_75t_L g2006 ( 
.A1(n_1958),
.A2(n_1824),
.B(n_1867),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1931),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1888),
.B(n_1754),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1891),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1891),
.B(n_1754),
.Y(n_2010)
);

OAI21x1_ASAP7_75t_L g2011 ( 
.A1(n_1964),
.A2(n_1880),
.B(n_1819),
.Y(n_2011)
);

A2O1A1Ixp33_ASAP7_75t_L g2012 ( 
.A1(n_1913),
.A2(n_1882),
.B(n_1864),
.C(n_1881),
.Y(n_2012)
);

AOI21xp33_ASAP7_75t_L g2013 ( 
.A1(n_1919),
.A2(n_1813),
.B(n_1820),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1929),
.Y(n_2014)
);

OAI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1950),
.A2(n_1919),
.B1(n_1973),
.B2(n_1917),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1908),
.B(n_1791),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1946),
.Y(n_2017)
);

AOI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1961),
.A2(n_1889),
.B(n_1906),
.Y(n_2018)
);

AOI222xp33_ASAP7_75t_L g2019 ( 
.A1(n_1941),
.A2(n_1816),
.B1(n_1822),
.B2(n_1855),
.C1(n_1805),
.C2(n_1874),
.Y(n_2019)
);

AO21x2_ASAP7_75t_L g2020 ( 
.A1(n_1985),
.A2(n_1861),
.B(n_1783),
.Y(n_2020)
);

OAI21x1_ASAP7_75t_L g2021 ( 
.A1(n_1890),
.A2(n_1788),
.B(n_1742),
.Y(n_2021)
);

BUFx2_ASAP7_75t_L g2022 ( 
.A(n_1912),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1918),
.Y(n_2023)
);

OA21x2_ASAP7_75t_L g2024 ( 
.A1(n_1921),
.A2(n_1886),
.B(n_1759),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1980),
.B(n_1781),
.Y(n_2025)
);

OAI21x1_ASAP7_75t_L g2026 ( 
.A1(n_1927),
.A2(n_1824),
.B(n_1870),
.Y(n_2026)
);

AOI21x1_ASAP7_75t_L g2027 ( 
.A1(n_1899),
.A2(n_1793),
.B(n_1752),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1935),
.Y(n_2028)
);

AOI21x1_ASAP7_75t_L g2029 ( 
.A1(n_1894),
.A2(n_1827),
.B(n_1840),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1930),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1930),
.B(n_1780),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1895),
.B(n_1849),
.Y(n_2032)
);

OAI21x1_ASAP7_75t_L g2033 ( 
.A1(n_1914),
.A2(n_1934),
.B(n_1923),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1937),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1902),
.A2(n_1739),
.B(n_1869),
.Y(n_2035)
);

OA21x2_ASAP7_75t_L g2036 ( 
.A1(n_1981),
.A2(n_1811),
.B(n_1849),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1889),
.A2(n_1849),
.B(n_1755),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2022),
.Y(n_2038)
);

OA21x2_ASAP7_75t_L g2039 ( 
.A1(n_2000),
.A2(n_1932),
.B(n_1969),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1992),
.B(n_2016),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2022),
.Y(n_2041)
);

INVx1_ASAP7_75t_SL g2042 ( 
.A(n_2005),
.Y(n_2042)
);

OAI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_2018),
.A2(n_1941),
.B(n_1909),
.Y(n_2043)
);

OR2x6_ASAP7_75t_L g2044 ( 
.A(n_2003),
.B(n_1943),
.Y(n_2044)
);

AO21x2_ASAP7_75t_L g2045 ( 
.A1(n_2037),
.A2(n_1962),
.B(n_1952),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_2004),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_2009),
.B(n_1947),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_2032),
.B(n_1949),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1992),
.B(n_1900),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_2030),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1992),
.B(n_1900),
.Y(n_2051)
);

BUFx6f_ASAP7_75t_L g2052 ( 
.A(n_2035),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1996),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2028),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_1995),
.Y(n_2055)
);

OAI21x1_ASAP7_75t_L g2056 ( 
.A1(n_2000),
.A2(n_1944),
.B(n_1957),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2034),
.Y(n_2057)
);

OR2x6_ASAP7_75t_L g2058 ( 
.A(n_2035),
.B(n_1896),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2017),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2017),
.Y(n_2060)
);

INVx4_ASAP7_75t_L g2061 ( 
.A(n_2023),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2016),
.B(n_1907),
.Y(n_2062)
);

AO21x2_ASAP7_75t_L g2063 ( 
.A1(n_1995),
.A2(n_2006),
.B(n_1994),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2031),
.B(n_1907),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_2043),
.A2(n_2015),
.B1(n_1994),
.B2(n_2013),
.Y(n_2065)
);

OAI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_2043),
.A2(n_2002),
.B1(n_1997),
.B2(n_1948),
.C(n_1951),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_2045),
.A2(n_2012),
.B(n_1962),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_SL g2068 ( 
.A1(n_2045),
.A2(n_2036),
.B1(n_1917),
.B2(n_1988),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2050),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2050),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_2045),
.A2(n_1948),
.B1(n_1951),
.B2(n_2036),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2049),
.B(n_2008),
.Y(n_2072)
);

AOI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_2045),
.A2(n_2036),
.B1(n_1973),
.B2(n_2019),
.Y(n_2073)
);

OAI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_2056),
.A2(n_2012),
.B(n_1997),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2050),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2050),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2046),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2049),
.B(n_2008),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2049),
.B(n_2010),
.Y(n_2079)
);

OAI33xp33_ASAP7_75t_L g2080 ( 
.A1(n_2048),
.A2(n_1990),
.A3(n_1959),
.B1(n_1993),
.B2(n_1978),
.B3(n_2001),
.Y(n_2080)
);

OAI211xp5_ASAP7_75t_SL g2081 ( 
.A1(n_2042),
.A2(n_1986),
.B(n_1988),
.C(n_1953),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_SL g2082 ( 
.A1(n_2045),
.A2(n_1755),
.B1(n_1989),
.B2(n_2024),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2046),
.Y(n_2083)
);

OA21x2_ASAP7_75t_L g2084 ( 
.A1(n_2055),
.A2(n_2033),
.B(n_1998),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2042),
.B(n_2014),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2048),
.B(n_2007),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2040),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2087),
.Y(n_2088)
);

OAI221xp5_ASAP7_75t_L g2089 ( 
.A1(n_2065),
.A2(n_2025),
.B1(n_2029),
.B2(n_2058),
.C(n_1933),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2087),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2077),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_2072),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2072),
.B(n_2051),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2077),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_2074),
.B(n_2047),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2083),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2087),
.B(n_2038),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2095),
.B(n_2092),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2095),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2091),
.B(n_2078),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2095),
.B(n_2078),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2093),
.B(n_2068),
.Y(n_2102)
);

OAI221xp5_ASAP7_75t_L g2103 ( 
.A1(n_2089),
.A2(n_2074),
.B1(n_2066),
.B2(n_2073),
.C(n_2071),
.Y(n_2103)
);

AOI31xp33_ASAP7_75t_L g2104 ( 
.A1(n_2103),
.A2(n_2080),
.A3(n_2067),
.B(n_2082),
.Y(n_2104)
);

OAI211xp5_ASAP7_75t_L g2105 ( 
.A1(n_2102),
.A2(n_2081),
.B(n_1966),
.C(n_1954),
.Y(n_2105)
);

OAI21x1_ASAP7_75t_L g2106 ( 
.A1(n_2099),
.A2(n_2094),
.B(n_2090),
.Y(n_2106)
);

AOI211xp5_ASAP7_75t_L g2107 ( 
.A1(n_2098),
.A2(n_1966),
.B(n_1954),
.C(n_1965),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_2100),
.Y(n_2108)
);

OAI31xp33_ASAP7_75t_L g2109 ( 
.A1(n_2101),
.A2(n_2051),
.A3(n_2085),
.B(n_2093),
.Y(n_2109)
);

OAI21xp33_ASAP7_75t_L g2110 ( 
.A1(n_2100),
.A2(n_2051),
.B(n_2086),
.Y(n_2110)
);

NOR2xp67_ASAP7_75t_L g2111 ( 
.A(n_2098),
.B(n_2096),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2099),
.B(n_2079),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2112),
.B(n_2088),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_2108),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2106),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2111),
.B(n_2088),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2108),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_2106),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2105),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2104),
.B(n_2079),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2109),
.B(n_2110),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2107),
.B(n_2094),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2104),
.B(n_1915),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2114),
.B(n_2117),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2119),
.B(n_1936),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2114),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2122),
.B(n_2090),
.Y(n_2127)
);

INVx1_ASAP7_75t_SL g2128 ( 
.A(n_2123),
.Y(n_2128)
);

INVxp67_ASAP7_75t_L g2129 ( 
.A(n_2120),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2113),
.B(n_2121),
.Y(n_2130)
);

INVx1_ASAP7_75t_SL g2131 ( 
.A(n_2118),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_2125),
.B(n_1936),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2129),
.B(n_2113),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2126),
.Y(n_2134)
);

OAI22xp33_ASAP7_75t_L g2135 ( 
.A1(n_2128),
.A2(n_2115),
.B1(n_2116),
.B2(n_2058),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2134),
.B(n_2130),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2133),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_2135),
.B(n_2131),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2132),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2136),
.Y(n_2140)
);

XNOR2xp5_ASAP7_75t_L g2141 ( 
.A(n_2139),
.B(n_2124),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2137),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2138),
.Y(n_2143)
);

OAI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_2138),
.A2(n_2124),
.B(n_2127),
.Y(n_2144)
);

OAI21xp33_ASAP7_75t_L g2145 ( 
.A1(n_2143),
.A2(n_2115),
.B(n_2116),
.Y(n_2145)
);

OAI322xp33_ASAP7_75t_L g2146 ( 
.A1(n_2141),
.A2(n_1903),
.A3(n_1910),
.B1(n_1858),
.B2(n_2097),
.C1(n_1926),
.C2(n_1976),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2144),
.A2(n_1939),
.B(n_1928),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2142),
.B(n_1967),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2140),
.B(n_1903),
.Y(n_2149)
);

OA21x2_ASAP7_75t_L g2150 ( 
.A1(n_2144),
.A2(n_2097),
.B(n_1928),
.Y(n_2150)
);

NOR2xp33_ASAP7_75t_L g2151 ( 
.A(n_2143),
.B(n_1925),
.Y(n_2151)
);

AOI211xp5_ASAP7_75t_L g2152 ( 
.A1(n_2143),
.A2(n_1911),
.B(n_1925),
.C(n_1945),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_2143),
.B(n_1972),
.Y(n_2153)
);

NAND3xp33_ASAP7_75t_L g2154 ( 
.A(n_2143),
.B(n_1911),
.C(n_1956),
.Y(n_2154)
);

OAI211xp5_ASAP7_75t_L g2155 ( 
.A1(n_2145),
.A2(n_1972),
.B(n_1789),
.C(n_1970),
.Y(n_2155)
);

OAI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_2153),
.A2(n_2061),
.B1(n_2058),
.B2(n_2052),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2148),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2149),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2154),
.A2(n_2061),
.B1(n_2058),
.B2(n_2052),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_2147),
.B(n_2052),
.Y(n_2160)
);

OAI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2151),
.A2(n_2061),
.B1(n_2058),
.B2(n_2052),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2152),
.B(n_2083),
.Y(n_2162)
);

AOI22x1_ASAP7_75t_L g2163 ( 
.A1(n_2146),
.A2(n_2150),
.B1(n_1956),
.B2(n_1945),
.Y(n_2163)
);

A2O1A1Ixp33_ASAP7_75t_L g2164 ( 
.A1(n_2153),
.A2(n_1924),
.B(n_1940),
.C(n_1904),
.Y(n_2164)
);

OAI32xp33_ASAP7_75t_L g2165 ( 
.A1(n_2153),
.A2(n_2061),
.A3(n_1970),
.B1(n_1975),
.B2(n_1982),
.Y(n_2165)
);

OAI21xp33_ASAP7_75t_SL g2166 ( 
.A1(n_2153),
.A2(n_2069),
.B(n_2075),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2145),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2167),
.A2(n_1924),
.B1(n_1940),
.B2(n_1755),
.Y(n_2168)
);

AOI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_2158),
.A2(n_2061),
.B1(n_2058),
.B2(n_2052),
.Y(n_2169)
);

AOI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_2160),
.A2(n_1963),
.B(n_2024),
.Y(n_2170)
);

NOR2x1_ASAP7_75t_L g2171 ( 
.A(n_2157),
.B(n_263),
.Y(n_2171)
);

O2A1O1Ixp33_ASAP7_75t_L g2172 ( 
.A1(n_2165),
.A2(n_264),
.B(n_265),
.C(n_266),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2163),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_2166),
.A2(n_1963),
.B(n_2024),
.Y(n_2174)
);

NAND2xp33_ASAP7_75t_R g2175 ( 
.A(n_2162),
.B(n_266),
.Y(n_2175)
);

OAI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2156),
.A2(n_2027),
.B(n_2021),
.Y(n_2176)
);

A2O1A1Ixp33_ASAP7_75t_L g2177 ( 
.A1(n_2164),
.A2(n_1975),
.B(n_1982),
.C(n_2056),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2155),
.Y(n_2178)
);

AOI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_2159),
.A2(n_2161),
.B(n_1963),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2167),
.A2(n_2058),
.B1(n_2052),
.B2(n_2084),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2173),
.B(n_2171),
.Y(n_2181)
);

OAI31xp33_ASAP7_75t_L g2182 ( 
.A1(n_2178),
.A2(n_267),
.A3(n_268),
.B(n_269),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2175),
.A2(n_2052),
.B1(n_1918),
.B2(n_2084),
.Y(n_2183)
);

AOI221xp5_ASAP7_75t_L g2184 ( 
.A1(n_2172),
.A2(n_2052),
.B1(n_1863),
.B2(n_1760),
.C(n_274),
.Y(n_2184)
);

OAI22xp33_ASAP7_75t_L g2185 ( 
.A1(n_2180),
.A2(n_1918),
.B1(n_2023),
.B2(n_1760),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2168),
.B(n_2084),
.Y(n_2186)
);

NOR2x1_ASAP7_75t_L g2187 ( 
.A(n_2177),
.B(n_270),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2169),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2179),
.B(n_2070),
.Y(n_2189)
);

AOI211xp5_ASAP7_75t_L g2190 ( 
.A1(n_2176),
.A2(n_270),
.B(n_272),
.C(n_273),
.Y(n_2190)
);

AOI221xp5_ASAP7_75t_L g2191 ( 
.A1(n_2170),
.A2(n_1863),
.B1(n_273),
.B2(n_274),
.C(n_275),
.Y(n_2191)
);

AOI221xp5_ASAP7_75t_L g2192 ( 
.A1(n_2174),
.A2(n_1863),
.B1(n_275),
.B2(n_276),
.C(n_277),
.Y(n_2192)
);

NOR2x1_ASAP7_75t_L g2193 ( 
.A(n_2181),
.B(n_272),
.Y(n_2193)
);

AO22x2_ASAP7_75t_L g2194 ( 
.A1(n_2188),
.A2(n_2182),
.B1(n_2189),
.B2(n_2184),
.Y(n_2194)
);

INVx1_ASAP7_75t_SL g2195 ( 
.A(n_2187),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2190),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2186),
.Y(n_2197)
);

NOR2xp67_ASAP7_75t_L g2198 ( 
.A(n_2183),
.B(n_276),
.Y(n_2198)
);

INVxp33_ASAP7_75t_SL g2199 ( 
.A(n_2192),
.Y(n_2199)
);

AO22x2_ASAP7_75t_L g2200 ( 
.A1(n_2191),
.A2(n_2076),
.B1(n_2069),
.B2(n_2075),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2185),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2181),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2181),
.Y(n_2203)
);

AOI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_2181),
.A2(n_1918),
.B1(n_2023),
.B2(n_2084),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2181),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_2181),
.B(n_277),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_2202),
.A2(n_2023),
.B1(n_2063),
.B2(n_2076),
.Y(n_2207)
);

NOR4xp75_ASAP7_75t_L g2208 ( 
.A(n_2199),
.B(n_278),
.C(n_279),
.D(n_280),
.Y(n_2208)
);

BUFx2_ASAP7_75t_L g2209 ( 
.A(n_2193),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2203),
.B(n_2070),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2195),
.B(n_281),
.Y(n_2211)
);

NAND4xp75_ASAP7_75t_L g2212 ( 
.A(n_2206),
.B(n_281),
.C(n_282),
.D(n_283),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2205),
.B(n_2062),
.Y(n_2213)
);

OAI322xp33_ASAP7_75t_L g2214 ( 
.A1(n_2201),
.A2(n_282),
.A3(n_283),
.B1(n_284),
.B2(n_285),
.C1(n_287),
.C2(n_288),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2194),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2196),
.B(n_287),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2198),
.B(n_290),
.Y(n_2217)
);

INVxp67_ASAP7_75t_L g2218 ( 
.A(n_2197),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2204),
.B(n_290),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2200),
.B(n_291),
.Y(n_2220)
);

AOI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_2202),
.A2(n_2023),
.B1(n_2063),
.B2(n_2020),
.Y(n_2221)
);

NOR3xp33_ASAP7_75t_L g2222 ( 
.A(n_2202),
.B(n_291),
.C(n_293),
.Y(n_2222)
);

NOR4xp25_ASAP7_75t_L g2223 ( 
.A(n_2195),
.B(n_294),
.C(n_295),
.D(n_296),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2193),
.Y(n_2224)
);

NAND2x1_ASAP7_75t_L g2225 ( 
.A(n_2193),
.B(n_1987),
.Y(n_2225)
);

AOI22xp33_ASAP7_75t_L g2226 ( 
.A1(n_2215),
.A2(n_2063),
.B1(n_1887),
.B2(n_2020),
.Y(n_2226)
);

AOI22x1_ASAP7_75t_L g2227 ( 
.A1(n_2209),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_2227)
);

OAI221xp5_ASAP7_75t_L g2228 ( 
.A1(n_2223),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.C(n_301),
.Y(n_2228)
);

NOR3xp33_ASAP7_75t_L g2229 ( 
.A(n_2211),
.B(n_298),
.C(n_299),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_2224),
.B(n_300),
.Y(n_2230)
);

AOI211xp5_ASAP7_75t_L g2231 ( 
.A1(n_2218),
.A2(n_301),
.B(n_302),
.C(n_303),
.Y(n_2231)
);

AOI221xp5_ASAP7_75t_L g2232 ( 
.A1(n_2220),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.C(n_305),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2216),
.Y(n_2233)
);

NAND3xp33_ASAP7_75t_SL g2234 ( 
.A(n_2208),
.B(n_304),
.C(n_306),
.Y(n_2234)
);

OAI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_2217),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.C(n_1987),
.Y(n_2235)
);

NOR3xp33_ASAP7_75t_SL g2236 ( 
.A(n_2214),
.B(n_307),
.C(n_1960),
.Y(n_2236)
);

AO221x1_ASAP7_75t_L g2237 ( 
.A1(n_2212),
.A2(n_1887),
.B1(n_2038),
.B2(n_2041),
.C(n_2054),
.Y(n_2237)
);

NAND4xp75_ASAP7_75t_L g2238 ( 
.A(n_2233),
.B(n_2210),
.C(n_2213),
.D(n_2207),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_2229),
.B(n_2222),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2230),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_2234),
.B(n_2228),
.Y(n_2241)
);

OAI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2236),
.A2(n_2219),
.B(n_2225),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2230),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2227),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2232),
.B(n_2221),
.Y(n_2245)
);

XOR2x1_ASAP7_75t_L g2246 ( 
.A(n_2231),
.B(n_1987),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2237),
.B(n_2064),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2235),
.Y(n_2248)
);

XNOR2xp5_ASAP7_75t_L g2249 ( 
.A(n_2226),
.B(n_1907),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2230),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2236),
.B(n_2064),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2240),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2250),
.Y(n_2253)
);

OR3x2_ASAP7_75t_L g2254 ( 
.A(n_2243),
.B(n_2006),
.C(n_1991),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2241),
.A2(n_2063),
.B1(n_2020),
.B2(n_2041),
.Y(n_2255)
);

AOI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_2242),
.A2(n_2063),
.B(n_1916),
.Y(n_2256)
);

NOR2xp67_ASAP7_75t_L g2257 ( 
.A(n_2244),
.B(n_2054),
.Y(n_2257)
);

OAI22x1_ASAP7_75t_L g2258 ( 
.A1(n_2239),
.A2(n_1916),
.B1(n_2055),
.B2(n_2060),
.Y(n_2258)
);

AOI21xp5_ASAP7_75t_L g2259 ( 
.A1(n_2245),
.A2(n_1916),
.B(n_2021),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2251),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2246),
.Y(n_2261)
);

XNOR2xp5_ASAP7_75t_L g2262 ( 
.A(n_2238),
.B(n_2026),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2239),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2253),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2252),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2260),
.Y(n_2266)
);

XNOR2xp5_ASAP7_75t_L g2267 ( 
.A(n_2263),
.B(n_2248),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2257),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2261),
.Y(n_2269)
);

OAI221xp5_ASAP7_75t_L g2270 ( 
.A1(n_2262),
.A2(n_2249),
.B1(n_2247),
.B2(n_2057),
.C(n_2053),
.Y(n_2270)
);

XOR2x1_ASAP7_75t_L g2271 ( 
.A(n_2254),
.B(n_2039),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_2259),
.B(n_2053),
.Y(n_2272)
);

OAI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2256),
.A2(n_2026),
.B(n_2056),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2264),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2265),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2267),
.Y(n_2276)
);

OAI21x1_ASAP7_75t_L g2277 ( 
.A1(n_2268),
.A2(n_2266),
.B(n_2269),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2272),
.B(n_2255),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2270),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2271),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2273),
.Y(n_2281)
);

BUFx2_ASAP7_75t_L g2282 ( 
.A(n_2275),
.Y(n_2282)
);

AOI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2274),
.A2(n_2258),
.B(n_2039),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2276),
.B(n_1968),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2277),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2280),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2279),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2278),
.A2(n_2281),
.B1(n_2057),
.B2(n_2059),
.Y(n_2288)
);

AOI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2287),
.A2(n_2064),
.B1(n_2062),
.B2(n_2060),
.Y(n_2289)
);

NOR2x1_ASAP7_75t_L g2290 ( 
.A(n_2285),
.B(n_1999),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_2282),
.B(n_2039),
.Y(n_2291)
);

OAI221xp5_ASAP7_75t_SL g2292 ( 
.A1(n_2286),
.A2(n_2060),
.B1(n_2059),
.B2(n_2044),
.C(n_1991),
.Y(n_2292)
);

OA21x2_ASAP7_75t_L g2293 ( 
.A1(n_2291),
.A2(n_2283),
.B(n_2284),
.Y(n_2293)
);

AOI22xp33_ASAP7_75t_SL g2294 ( 
.A1(n_2293),
.A2(n_2288),
.B1(n_2290),
.B2(n_2292),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_SL g2295 ( 
.A1(n_2294),
.A2(n_2289),
.B1(n_1999),
.B2(n_2039),
.Y(n_2295)
);

AOI22xp33_ASAP7_75t_L g2296 ( 
.A1(n_2294),
.A2(n_2039),
.B1(n_1999),
.B2(n_1989),
.Y(n_2296)
);

OAI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_2295),
.A2(n_2011),
.B(n_2033),
.Y(n_2297)
);

OAI22xp5_ASAP7_75t_L g2298 ( 
.A1(n_2297),
.A2(n_2296),
.B1(n_2044),
.B2(n_2059),
.Y(n_2298)
);

AOI211xp5_ASAP7_75t_L g2299 ( 
.A1(n_2298),
.A2(n_2011),
.B(n_1998),
.C(n_2062),
.Y(n_2299)
);


endmodule