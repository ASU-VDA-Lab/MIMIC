module fake_jpeg_8504_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_40),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_37),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_33),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_60),
.Y(n_92)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_29),
.Y(n_77)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_33),
.B1(n_23),
.B2(n_34),
.Y(n_66)
);

OAI22x1_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_73),
.B1(n_76),
.B2(n_80),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_33),
.B1(n_37),
.B2(n_23),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_37),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_17),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_33),
.B1(n_23),
.B2(n_34),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_23),
.B1(n_34),
.B2(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_29),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_43),
.B1(n_37),
.B2(n_29),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_30),
.B1(n_25),
.B2(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_36),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_19),
.B1(n_32),
.B2(n_30),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_46),
.B(n_37),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_36),
.C(n_35),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_39),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_99),
.Y(n_126)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_96),
.B(n_101),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_79),
.B1(n_86),
.B2(n_72),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_83),
.B1(n_92),
.B2(n_74),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_112),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_110),
.B1(n_82),
.B2(n_89),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_46),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_35),
.C(n_61),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_63),
.C(n_59),
.Y(n_117)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_69),
.A2(n_19),
.A3(n_32),
.B1(n_25),
.B2(n_30),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_17),
.A3(n_67),
.B1(n_27),
.B2(n_31),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_26),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_83),
.B1(n_69),
.B2(n_92),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_129),
.B(n_144),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_146),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_17),
.B(n_19),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_110),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_138),
.A2(n_122),
.B1(n_136),
.B2(n_137),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_74),
.B1(n_67),
.B2(n_81),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_68),
.B1(n_64),
.B2(n_87),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_65),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_26),
.B(n_20),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_21),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_103),
.A2(n_98),
.A3(n_99),
.B1(n_112),
.B2(n_100),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_96),
.A2(n_89),
.B1(n_49),
.B2(n_48),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_105),
.B1(n_87),
.B2(n_113),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_26),
.B(n_20),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_26),
.B(n_20),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_104),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_151),
.B(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_161),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_156),
.B1(n_178),
.B2(n_144),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_104),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_16),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_163),
.C(n_173),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_128),
.B(n_18),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_172),
.B(n_148),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_109),
.C(n_108),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_122),
.B1(n_139),
.B2(n_133),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_24),
.Y(n_165)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_18),
.B1(n_28),
.B2(n_64),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_167),
.A2(n_168),
.B1(n_165),
.B2(n_171),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_28),
.B1(n_31),
.B2(n_27),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_95),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_170),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_24),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_175),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_1),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_16),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_95),
.C(n_24),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_95),
.C(n_88),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_126),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_177),
.Y(n_207)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_16),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_145),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_185),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_149),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_7),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_162),
.B1(n_166),
.B2(n_152),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_191),
.C(n_193),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_150),
.A2(n_166),
.B1(n_156),
.B2(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_190),
.A2(n_167),
.B1(n_124),
.B2(n_139),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_125),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_125),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_197),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_121),
.B(n_31),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_155),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_204),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_138),
.B1(n_129),
.B2(n_135),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_206),
.B1(n_200),
.B2(n_205),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_125),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_152),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_130),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_121),
.B1(n_135),
.B2(n_27),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_214),
.B(n_215),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_213),
.C(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_153),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_153),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_228),
.C(n_189),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_208),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_225),
.B1(n_229),
.B2(n_232),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_224),
.B(n_207),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_124),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_233),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_199),
.B1(n_198),
.B2(n_204),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_26),
.Y(n_226)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_26),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_195),
.A2(n_88),
.B1(n_31),
.B2(n_27),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_230),
.A2(n_206),
.B1(n_184),
.B2(n_182),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_228),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_216),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_222),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_202),
.B(n_206),
.C(n_188),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_211),
.B(n_232),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_182),
.C(n_2),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_248),
.C(n_249),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_1),
.C(n_2),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_2),
.C(n_3),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_251),
.Y(n_258)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_220),
.A2(n_8),
.B1(n_14),
.B2(n_12),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_3),
.C(n_4),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_4),
.C(n_5),
.Y(n_269)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_261),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_233),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_249),
.C(n_234),
.Y(n_271)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_8),
.Y(n_267)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_240),
.B(n_8),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_263),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_256),
.A2(n_235),
.B1(n_253),
.B2(n_238),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_254),
.B1(n_268),
.B2(n_238),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_234),
.C(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_283),
.C(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_238),
.C(n_10),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_292),
.Y(n_299)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_295),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_283),
.B1(n_274),
.B2(n_279),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_262),
.B(n_269),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_290),
.A2(n_291),
.B(n_294),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_262),
.B(n_10),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_7),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_10),
.B(n_12),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_278),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_300),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_281),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_272),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_295),
.C(n_301),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_298),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_15),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_285),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_310),
.A2(n_284),
.B(n_279),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_313),
.B(n_309),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_314),
.A2(n_312),
.B(n_310),
.Y(n_315)
);

OAI321xp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_308),
.A3(n_306),
.B1(n_305),
.B2(n_15),
.C(n_6),
.Y(n_316)
);

AOI21x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_4),
.B(n_5),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_4),
.B(n_5),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_5),
.B1(n_6),
.B2(n_317),
.Y(n_319)
);


endmodule