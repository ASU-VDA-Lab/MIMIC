module fake_jpeg_28598_n_508 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_508);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_508;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_68),
.Y(n_107)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_61),
.Y(n_120)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_65),
.B(n_67),
.Y(n_122)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_14),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g151 ( 
.A(n_70),
.Y(n_151)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_75),
.Y(n_125)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_32),
.B(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_79),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_80),
.B(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_81),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_32),
.B(n_0),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_103),
.B(n_44),
.Y(n_105)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_105),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_62),
.A2(n_44),
.B1(n_43),
.B2(n_49),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_116),
.A2(n_150),
.B1(n_155),
.B2(n_157),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_87),
.A2(n_26),
.B1(n_33),
.B2(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_88),
.B1(n_64),
.B2(n_77),
.Y(n_166)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_101),
.B(n_26),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_100),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_56),
.B(n_35),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_161),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_81),
.A2(n_43),
.B1(n_49),
.B2(n_35),
.Y(n_150)
);

INVx6_ASAP7_75t_SL g154 ( 
.A(n_69),
.Y(n_154)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_72),
.A2(n_49),
.B1(n_33),
.B2(n_45),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_63),
.A2(n_28),
.B(n_46),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_105),
.C(n_120),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_83),
.A2(n_46),
.B1(n_41),
.B2(n_39),
.Y(n_157)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_84),
.B(n_41),
.Y(n_161)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

INVx4_ASAP7_75t_SL g207 ( 
.A(n_163),
.Y(n_207)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_165),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_113),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_171),
.B(n_184),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_106),
.B(n_52),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_173),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_107),
.B(n_34),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_120),
.B(n_39),
.C(n_34),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_183),
.Y(n_221)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

CKINVDCx12_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

BUFx24_ASAP7_75t_L g250 ( 
.A(n_181),
.Y(n_250)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_146),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_122),
.B(n_48),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_151),
.A2(n_104),
.B1(n_55),
.B2(n_99),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_185),
.A2(n_210),
.B1(n_211),
.B2(n_220),
.Y(n_227)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_122),
.B(n_37),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_199),
.Y(n_230)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_113),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_200),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_52),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_153),
.B(n_48),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_130),
.B(n_37),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_209),
.Y(n_251)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

BUFx24_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_137),
.Y(n_206)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_133),
.A2(n_102),
.B1(n_89),
.B2(n_74),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_128),
.A2(n_74),
.B1(n_82),
.B2(n_45),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_212),
.B(n_213),
.Y(n_259)
);

CKINVDCx12_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_136),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_116),
.A2(n_98),
.B1(n_96),
.B2(n_92),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_124),
.B1(n_123),
.B2(n_126),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_114),
.B(n_33),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_216),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_114),
.B(n_45),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_125),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_139),
.B(n_82),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_218),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_124),
.Y(n_240)
);

AO22x1_ASAP7_75t_SL g220 ( 
.A1(n_155),
.A2(n_90),
.B1(n_86),
.B2(n_85),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_225),
.B(n_145),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_255),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_178),
.B(n_204),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_237),
.A2(n_211),
.B(n_185),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_240),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_169),
.B(n_138),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_167),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_126),
.B1(n_138),
.B2(n_142),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_117),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_179),
.C(n_195),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_194),
.A2(n_152),
.B1(n_66),
.B2(n_91),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_207),
.B1(n_206),
.B2(n_208),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_266),
.Y(n_332)
);

OR2x4_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_177),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g304 ( 
.A1(n_267),
.A2(n_274),
.B(n_291),
.Y(n_304)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_269),
.Y(n_334)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_270),
.B(n_271),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_165),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_259),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_276),
.Y(n_305)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_279),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_L g274 ( 
.A1(n_232),
.A2(n_229),
.B(n_225),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_275),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_186),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_186),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_278),
.Y(n_306)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_189),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_282),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_281),
.B(n_287),
.Y(n_335)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_245),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_221),
.B(n_191),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_286),
.Y(n_318)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_284),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_260),
.A2(n_166),
.B1(n_188),
.B2(n_180),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_285),
.A2(n_233),
.B1(n_286),
.B2(n_299),
.Y(n_311)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_292),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_296),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_236),
.A2(n_111),
.B1(n_207),
.B2(n_201),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_290),
.A2(n_261),
.B(n_253),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_222),
.B(n_0),
.Y(n_291)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_247),
.B(n_0),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_294),
.Y(n_321)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_228),
.B(n_191),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_301),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_230),
.B(n_212),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_254),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_233),
.A2(n_210),
.B1(n_149),
.B2(n_205),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_299),
.A2(n_261),
.B(n_243),
.Y(n_326)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_231),
.B(n_1),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_302),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_230),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_310),
.C(n_314),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_230),
.C(n_281),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_317),
.B1(n_325),
.B2(n_328),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_227),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_297),
.A2(n_227),
.B1(n_255),
.B2(n_240),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_316),
.A2(n_278),
.B1(n_235),
.B2(n_168),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_297),
.A2(n_234),
.B1(n_240),
.B2(n_258),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_252),
.C(n_256),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_320),
.B(n_331),
.C(n_333),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_258),
.Y(n_324)
);

OA22x2_ASAP7_75t_L g344 ( 
.A1(n_324),
.A2(n_243),
.B1(n_287),
.B2(n_279),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_297),
.A2(n_267),
.B1(n_293),
.B2(n_266),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_283),
.A2(n_242),
.B1(n_219),
.B2(n_197),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_269),
.B(n_301),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_273),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_270),
.B(n_250),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_268),
.B(n_250),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_337),
.B(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_321),
.B(n_291),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_245),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_351),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_319),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_341),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_318),
.A2(n_282),
.B(n_294),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_342),
.A2(n_343),
.B(n_353),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_344),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_345),
.A2(n_354),
.B1(n_364),
.B2(n_343),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_275),
.Y(n_347)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_350),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_336),
.B(n_250),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_313),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_352),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_292),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_316),
.A2(n_314),
.B1(n_332),
.B2(n_318),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_326),
.A2(n_288),
.B(n_249),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_355),
.A2(n_324),
.B(n_329),
.Y(n_372)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_357),
.Y(n_390)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_322),
.Y(n_358)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_305),
.A2(n_265),
.B1(n_246),
.B2(n_248),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_359),
.A2(n_328),
.B1(n_345),
.B2(n_317),
.Y(n_370)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_360),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_327),
.B(n_288),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_361),
.B(n_352),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_325),
.B(n_288),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_365),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_306),
.B(n_248),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_368),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_310),
.A2(n_246),
.B1(n_249),
.B2(n_164),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_1),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_334),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_312),
.B(n_284),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_307),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_312),
.B(n_164),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_370),
.A2(n_397),
.B1(n_344),
.B2(n_308),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_372),
.A2(n_348),
.B(n_347),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_361),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_391),
.Y(n_406)
);

NAND2x1_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_324),
.Y(n_374)
);

OAI21xp33_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_344),
.B(n_338),
.Y(n_410)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_376),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_315),
.Y(n_380)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_380),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_381),
.B(n_144),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_341),
.B(n_320),
.Y(n_386)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_333),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_356),
.Y(n_402)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_389),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_303),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_349),
.A2(n_311),
.B1(n_304),
.B2(n_303),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_393),
.A2(n_344),
.B1(n_358),
.B2(n_357),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_334),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_395),
.B(n_396),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_393),
.Y(n_398)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_346),
.C(n_367),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_404),
.C(n_405),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_356),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_400),
.B(n_408),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_417),
.Y(n_436)
);

AO22x2_ASAP7_75t_SL g403 ( 
.A1(n_382),
.A2(n_354),
.B1(n_342),
.B2(n_353),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_410),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_364),
.C(n_337),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_350),
.C(n_362),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_407),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_331),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_349),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_414),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_416),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_365),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_422),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_308),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_129),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_144),
.C(n_2),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_387),
.C(n_394),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_420),
.B(n_397),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_373),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_406),
.Y(n_424)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_424),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_426),
.B(n_441),
.Y(n_457)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_429),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_419),
.Y(n_458)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_431),
.Y(n_452)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_437),
.Y(n_447)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_403),
.A2(n_372),
.B(n_396),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_439),
.Y(n_446)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_418),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_383),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_420),
.B(n_384),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_402),
.B(n_384),
.C(n_378),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_442),
.B(n_404),
.C(n_405),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_399),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_445),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_403),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_453),
.C(n_454),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_387),
.C(n_392),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_458),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_423),
.A2(n_392),
.B1(n_398),
.B2(n_382),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_450),
.A2(n_370),
.B1(n_427),
.B2(n_383),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_417),
.C(n_379),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_371),
.C(n_369),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_439),
.Y(n_455)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_455),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

MAJx2_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_435),
.C(n_441),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_467),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_432),
.C(n_434),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_466),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_434),
.C(n_426),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_430),
.C(n_438),
.Y(n_467)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_468),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_425),
.C(n_435),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_457),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_446),
.A2(n_435),
.B(n_427),
.Y(n_470)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_470),
.Y(n_478)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_471),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_452),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g482 ( 
.A(n_472),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_371),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_473),
.A2(n_369),
.B1(n_394),
.B2(n_390),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_465),
.Y(n_475)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_475),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_447),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_477),
.B(n_479),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_457),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_473),
.Y(n_481)
);

AOI31xp67_ASAP7_75t_L g492 ( 
.A1(n_481),
.A2(n_422),
.A3(n_374),
.B(n_6),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_483),
.B(n_459),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_484),
.A2(n_374),
.B(n_390),
.Y(n_488)
);

AOI321xp33_ASAP7_75t_L g486 ( 
.A1(n_482),
.A2(n_461),
.A3(n_410),
.B1(n_462),
.B2(n_460),
.C(n_467),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_486),
.B(n_489),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_492),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_491),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_459),
.C(n_464),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_466),
.C(n_469),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_474),
.C(n_478),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_498),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_476),
.C(n_484),
.Y(n_498)
);

OAI21xp33_ASAP7_75t_L g499 ( 
.A1(n_497),
.A2(n_488),
.B(n_4),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_499),
.A2(n_8),
.B(n_4),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_497),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_495),
.B1(n_496),
.B2(n_6),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_503),
.C(n_500),
.Y(n_504)
);

A2O1A1Ixp33_ASAP7_75t_SL g505 ( 
.A1(n_504),
.A2(n_1),
.B(n_6),
.C(n_7),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_505),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_6),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_7),
.C(n_387),
.Y(n_508)
);


endmodule