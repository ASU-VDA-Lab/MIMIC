module fake_jpeg_2609_n_580 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_580);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_61),
.Y(n_159)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_66),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_30),
.B(n_10),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_75),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_78),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_35),
.B(n_8),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_79),
.Y(n_191)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_82),
.Y(n_187)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_29),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_98),
.Y(n_153)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_42),
.B(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_117),
.Y(n_160)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_19),
.Y(n_111)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx5_ASAP7_75t_SL g139 ( 
.A(n_114),
.Y(n_139)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_33),
.Y(n_115)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_116),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_42),
.B(n_49),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_56),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_122),
.B(n_140),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_41),
.B1(n_52),
.B2(n_50),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_127),
.A2(n_151),
.B1(n_158),
.B2(n_170),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_40),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_72),
.A2(n_44),
.B1(n_33),
.B2(n_39),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_81),
.B(n_56),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_152),
.B(n_154),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_40),
.Y(n_154)
);

INVx5_ASAP7_75t_SL g155 ( 
.A(n_61),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_155),
.B(n_182),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_72),
.A2(n_44),
.B1(n_33),
.B2(n_39),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_94),
.B(n_37),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_164),
.B(n_173),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_83),
.A2(n_41),
.B1(n_52),
.B2(n_50),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_109),
.B(n_37),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_98),
.B(n_39),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_185),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_60),
.A2(n_26),
.B1(n_36),
.B2(n_24),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_184),
.B1(n_84),
.B2(n_38),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_89),
.B(n_55),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_64),
.A2(n_26),
.B1(n_36),
.B2(n_45),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_99),
.B(n_49),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_89),
.B(n_55),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_106),
.B(n_45),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_135),
.Y(n_193)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_195),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_196),
.Y(n_313)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_198),
.Y(n_278)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_199),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_128),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_200),
.B(n_211),
.Y(n_263)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_201),
.Y(n_298)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_202),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_130),
.B(n_77),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_206),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_108),
.B1(n_86),
.B2(n_79),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_207),
.A2(n_224),
.B1(n_228),
.B2(n_139),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_SL g208 ( 
.A(n_160),
.B(n_53),
.C(n_27),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_208),
.B(n_232),
.C(n_172),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_135),
.A2(n_53),
.B1(n_52),
.B2(n_50),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_209),
.A2(n_212),
.B1(n_241),
.B2(n_248),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_119),
.B(n_39),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_210),
.B(n_244),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_120),
.A2(n_38),
.B1(n_39),
.B2(n_27),
.Y(n_212)
);

INVx3_ASAP7_75t_SL g213 ( 
.A(n_142),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_213),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_148),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_214),
.B(n_215),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_216),
.B(n_220),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_73),
.B1(n_67),
.B2(n_75),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_218),
.A2(n_229),
.B1(n_237),
.B2(n_251),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_151),
.A2(n_101),
.B(n_115),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_219),
.A2(n_221),
.B(n_230),
.Y(n_308)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_221),
.B(n_226),
.Y(n_285)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_130),
.B(n_27),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_223),
.B(n_234),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_160),
.A2(n_113),
.B1(n_112),
.B2(n_38),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_225),
.A2(n_260),
.B1(n_237),
.B2(n_194),
.Y(n_286)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_184),
.A2(n_27),
.B1(n_48),
.B2(n_21),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_143),
.A2(n_147),
.B1(n_166),
.B2(n_162),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_126),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_230),
.B(n_231),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_129),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_27),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_233),
.B(n_235),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_186),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_180),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_236),
.B(n_252),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_120),
.A2(n_21),
.B1(n_11),
.B2(n_12),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_145),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_238),
.Y(n_282)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_175),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_239),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_134),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_240),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_123),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_150),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_243),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_124),
.B(n_0),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_158),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_245),
.A2(n_4),
.B1(n_249),
.B2(n_193),
.Y(n_304)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_153),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_246),
.B(n_250),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_125),
.B(n_1),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_259),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_163),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_159),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_153),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_132),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_187),
.B(n_6),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_121),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_183),
.B(n_1),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_255),
.B(n_169),
.Y(n_275)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_144),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_169),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_258),
.B1(n_137),
.B2(n_176),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_136),
.A2(n_5),
.B1(n_6),
.B2(n_12),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_179),
.B(n_3),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_131),
.A2(n_5),
.B1(n_6),
.B2(n_13),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_264),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_197),
.B(n_191),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_271),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_197),
.B(n_217),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_217),
.B(n_191),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_274),
.B(n_279),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_275),
.B(n_293),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_277),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_156),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_227),
.C(n_211),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_280),
.B(n_257),
.C(n_293),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_156),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_281),
.B(n_290),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_296),
.B1(n_299),
.B2(n_301),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_208),
.B(n_259),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_219),
.A2(n_228),
.B1(n_189),
.B2(n_167),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_225),
.A2(n_157),
.B1(n_189),
.B2(n_167),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_242),
.A2(n_141),
.B1(n_169),
.B2(n_3),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_207),
.A2(n_4),
.B1(n_13),
.B2(n_17),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_242),
.A2(n_4),
.B1(n_13),
.B2(n_17),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_255),
.B(n_13),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_308),
.B(n_299),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_244),
.A2(n_4),
.B1(n_255),
.B2(n_256),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_244),
.B(n_200),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_311),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_210),
.A2(n_4),
.B1(n_216),
.B2(n_214),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_318),
.B1(n_201),
.B2(n_235),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_304),
.A2(n_305),
.B1(n_310),
.B2(n_222),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_215),
.A2(n_213),
.B1(n_254),
.B2(n_198),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_210),
.A2(n_213),
.B1(n_202),
.B2(n_220),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_309),
.B1(n_253),
.B2(n_240),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_246),
.A2(n_250),
.B1(n_226),
.B2(n_243),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_196),
.A2(n_205),
.B1(n_206),
.B2(n_195),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_204),
.B(n_206),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_199),
.A2(n_239),
.B1(n_233),
.B2(n_238),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_321),
.Y(n_370)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_322),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_262),
.B(n_241),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_311),
.B(n_231),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_327),
.B(n_347),
.Y(n_369)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_328),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_329),
.B(n_335),
.C(n_344),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_330),
.Y(n_400)
);

INVx8_ASAP7_75t_L g331 ( 
.A(n_284),
.Y(n_331)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_262),
.B(n_273),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_271),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_298),
.Y(n_338)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_338),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_290),
.A2(n_264),
.B1(n_291),
.B2(n_269),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_339),
.A2(n_346),
.B1(n_323),
.B2(n_353),
.Y(n_403)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_342),
.Y(n_382)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_283),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_343),
.B(n_345),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_280),
.B(n_287),
.C(n_263),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_265),
.B(n_274),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_275),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_348),
.A2(n_351),
.B(n_268),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_285),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_354),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_287),
.B(n_263),
.C(n_265),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_350),
.B(n_357),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_308),
.A2(n_302),
.B(n_267),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_285),
.Y(n_354)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_358),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g357 ( 
.A(n_275),
.B(n_279),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_297),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_289),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_367),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_287),
.B(n_281),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_360),
.B(n_362),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_287),
.B(n_301),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_368),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_295),
.B(n_319),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_286),
.A2(n_294),
.B1(n_316),
.B2(n_296),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_363),
.A2(n_366),
.B1(n_314),
.B2(n_317),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_289),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_364),
.B(n_365),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_300),
.B(n_303),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_318),
.A2(n_315),
.B1(n_288),
.B2(n_314),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_297),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_307),
.B(n_270),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_351),
.A2(n_304),
.B(n_288),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_372),
.A2(n_375),
.B(n_376),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_315),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_373),
.B(n_387),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_321),
.A2(n_282),
.B(n_292),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_328),
.A2(n_282),
.B(n_292),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_330),
.A2(n_270),
.B(n_305),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_379),
.A2(n_388),
.B(n_389),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_361),
.B(n_309),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_386),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_332),
.B(n_307),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_348),
.A2(n_298),
.B(n_310),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_393),
.A2(n_399),
.B1(n_404),
.B2(n_378),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_362),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_401),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_363),
.A2(n_323),
.B1(n_353),
.B2(n_352),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_366),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_403),
.A2(n_313),
.B1(n_331),
.B2(n_312),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_352),
.A2(n_355),
.B1(n_339),
.B2(n_348),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_355),
.A2(n_314),
.B1(n_313),
.B2(n_312),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_407),
.A2(n_278),
.B1(n_381),
.B2(n_401),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_336),
.A2(n_341),
.B(n_344),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_408),
.A2(n_278),
.B(n_266),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_336),
.C(n_350),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_410),
.B(n_426),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_342),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_411),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_343),
.Y(n_413)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_413),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_370),
.B(n_359),
.Y(n_414)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_415),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_329),
.C(n_335),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_418),
.C(n_422),
.Y(n_447)
);

XOR2x1_ASAP7_75t_SL g417 ( 
.A(n_400),
.B(n_336),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_417),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_360),
.C(n_347),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_388),
.A2(n_357),
.B(n_322),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_382),
.Y(n_420)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_420),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_364),
.C(n_365),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_334),
.Y(n_423)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_423),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_340),
.C(n_337),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_425),
.C(n_442),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_405),
.B(n_345),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_400),
.A2(n_326),
.B(n_338),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g427 ( 
.A(n_374),
.B(n_338),
.CI(n_266),
.CON(n_427),
.SN(n_427)
);

OAI32xp33_ASAP7_75t_L g462 ( 
.A1(n_427),
.A2(n_371),
.A3(n_391),
.B1(n_384),
.B2(n_394),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_356),
.Y(n_429)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_429),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_430),
.A2(n_439),
.B1(n_389),
.B2(n_398),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_372),
.A2(n_266),
.B(n_313),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_433),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_383),
.A2(n_400),
.B1(n_381),
.B2(n_393),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_432),
.A2(n_441),
.B1(n_386),
.B2(n_403),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_375),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_435),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_436),
.B(n_379),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_372),
.A2(n_408),
.B(n_379),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_407),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_438),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_370),
.B(n_384),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_440),
.B(n_392),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_374),
.B(n_405),
.C(n_406),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_375),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_443),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_444),
.B(n_437),
.Y(n_482)
);

AOI22x1_ASAP7_75t_L g448 ( 
.A1(n_434),
.A2(n_378),
.B1(n_404),
.B2(n_399),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_448),
.A2(n_452),
.B1(n_453),
.B2(n_454),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_406),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_459),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_441),
.A2(n_409),
.B1(n_434),
.B2(n_426),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_369),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_409),
.A2(n_386),
.B1(n_371),
.B2(n_373),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_461),
.A2(n_465),
.B1(n_410),
.B2(n_424),
.Y(n_480)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_462),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_432),
.A2(n_369),
.B1(n_391),
.B2(n_394),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_416),
.B(n_376),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_472),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_439),
.A2(n_389),
.B1(n_376),
.B2(n_392),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_470),
.A2(n_412),
.B1(n_433),
.B2(n_431),
.Y(n_478)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_471),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_458),
.A2(n_415),
.B1(n_420),
.B2(n_435),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_474),
.A2(n_478),
.B1(n_480),
.B2(n_487),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_454),
.A2(n_419),
.B1(n_421),
.B2(n_443),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_489),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_482),
.B(n_486),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_442),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_485),
.Y(n_499)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_484),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_447),
.B(n_425),
.Y(n_485)
);

MAJx2_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_450),
.C(n_447),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_465),
.A2(n_421),
.B1(n_430),
.B2(n_423),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_445),
.A2(n_457),
.B1(n_464),
.B2(n_449),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_488),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_470),
.A2(n_413),
.B1(n_411),
.B2(n_427),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_473),
.A2(n_414),
.B(n_440),
.Y(n_490)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_490),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_461),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_492),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_472),
.A2(n_427),
.B1(n_429),
.B2(n_412),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_463),
.B(n_398),
.Y(n_494)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_494),
.Y(n_514)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_446),
.Y(n_495)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_495),
.Y(n_517)
);

FAx1_ASAP7_75t_SL g497 ( 
.A(n_466),
.B(n_417),
.CI(n_427),
.CON(n_497),
.SN(n_497)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_497),
.B(n_469),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_448),
.A2(n_412),
.B1(n_407),
.B2(n_438),
.Y(n_498)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_498),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_450),
.C(n_468),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_500),
.B(n_507),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_462),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_505),
.B(n_506),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_444),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_436),
.C(n_455),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_428),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_511),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_483),
.B(n_448),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_497),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_455),
.C(n_417),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_518),
.C(n_520),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_460),
.C(n_453),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_489),
.B(n_477),
.Y(n_520)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_501),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_528),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_494),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_529),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_506),
.B(n_482),
.Y(n_526)
);

XNOR2x1_ASAP7_75t_L g550 ( 
.A(n_526),
.B(n_537),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_503),
.A2(n_475),
.B1(n_479),
.B2(n_487),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_527),
.A2(n_530),
.B1(n_531),
.B2(n_533),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_508),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_446),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_519),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_500),
.B(n_492),
.C(n_495),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_532),
.B(n_536),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_504),
.B(n_484),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_502),
.A2(n_479),
.B(n_428),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_534),
.A2(n_510),
.B(n_507),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_499),
.B(n_467),
.C(n_385),
.Y(n_536)
);

XNOR2x1_ASAP7_75t_L g537 ( 
.A(n_509),
.B(n_497),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_536),
.B(n_511),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_539),
.B(n_542),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_540),
.A2(n_549),
.B(n_522),
.Y(n_556)
);

INVx11_ASAP7_75t_L g541 ( 
.A(n_533),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_547),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_499),
.C(n_518),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_523),
.B(n_476),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_544),
.B(n_545),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_521),
.B(n_505),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_535),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_527),
.A2(n_515),
.B1(n_520),
.B2(n_513),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_529),
.A2(n_515),
.B(n_516),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_534),
.A2(n_385),
.B1(n_402),
.B2(n_380),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_551),
.B(n_549),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_543),
.C(n_532),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_553),
.B(n_554),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_546),
.A2(n_530),
.B1(n_525),
.B2(n_537),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_555),
.B(n_558),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_559),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_539),
.B(n_535),
.C(n_522),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_560),
.B(n_561),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_540),
.A2(n_516),
.B(n_526),
.Y(n_561)
);

NOR2x1_ASAP7_75t_SL g562 ( 
.A(n_553),
.B(n_550),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_562),
.A2(n_567),
.B(n_568),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_552),
.B(n_550),
.C(n_548),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_554),
.B(n_538),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_564),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_569),
.A2(n_570),
.B(n_563),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_565),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_566),
.A2(n_557),
.B(n_556),
.Y(n_572)
);

AOI21xp33_ASAP7_75t_L g574 ( 
.A1(n_572),
.A2(n_567),
.B(n_541),
.Y(n_574)
);

AOI31xp33_ASAP7_75t_L g576 ( 
.A1(n_573),
.A2(n_558),
.A3(n_559),
.B(n_402),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_574),
.A2(n_571),
.B(n_548),
.Y(n_575)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_575),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_577),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_576),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_579),
.B(n_380),
.Y(n_580)
);


endmodule