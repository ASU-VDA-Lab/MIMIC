module fake_netlist_1_2911_n_552 (n_117, n_44, n_133, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_130, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_16, n_13, n_113, n_95, n_124, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_122, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_136, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_134, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_132, n_51, n_96, n_39, n_552);
input n_117;
input n_44;
input n_133;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_16;
input n_13;
input n_113;
input n_95;
input n_124;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_122;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_51;
input n_96;
input n_39;
output n_552;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_141;
wire n_517;
wire n_479;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_475;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_178;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_158;
wire n_524;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g137 ( .A(n_45), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_103), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_104), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_73), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_134), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_96), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_26), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_100), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_68), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_59), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_53), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_8), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_63), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_17), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_76), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_125), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_56), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_32), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_113), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_77), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_91), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_129), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_24), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_136), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_26), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_12), .Y(n_163) );
INVxp33_ASAP7_75t_L g164 ( .A(n_105), .Y(n_164) );
BUFx10_ASAP7_75t_L g165 ( .A(n_88), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_27), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_79), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_21), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_7), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_16), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_41), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_70), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_17), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_31), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_20), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_60), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_120), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_74), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_71), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_15), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_94), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_106), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_9), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_128), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_61), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_23), .Y(n_187) );
BUFx10_ASAP7_75t_L g188 ( .A(n_87), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_51), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_69), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_99), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_89), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_112), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_34), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_75), .Y(n_195) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_133), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_58), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_15), .Y(n_198) );
NOR2xp67_ASAP7_75t_L g199 ( .A(n_78), .B(n_102), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_64), .Y(n_200) );
NOR2xp67_ASAP7_75t_L g201 ( .A(n_18), .B(n_62), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_126), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_57), .Y(n_203) );
INVxp67_ASAP7_75t_L g204 ( .A(n_93), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_84), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_95), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_86), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_80), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_131), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_101), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_121), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_24), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_111), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_130), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_135), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_36), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_92), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_116), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_65), .Y(n_219) );
INVxp67_ASAP7_75t_L g220 ( .A(n_12), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_25), .Y(n_221) );
INVxp67_ASAP7_75t_L g222 ( .A(n_98), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_54), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_81), .Y(n_224) );
OR2x2_ASAP7_75t_L g225 ( .A(n_66), .B(n_85), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_72), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_127), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_11), .B(n_117), .Y(n_228) );
CKINVDCx14_ASAP7_75t_R g229 ( .A(n_37), .Y(n_229) );
XNOR2x2_ASAP7_75t_R g230 ( .A(n_31), .B(n_90), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_19), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_97), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_165), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_138), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_137), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_180), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_206), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_206), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_164), .B(n_0), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_180), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_206), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_137), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_141), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_164), .B(n_1), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_200), .B(n_1), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_206), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_140), .Y(n_247) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_140), .A2(n_47), .B(n_46), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_188), .B(n_2), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_154), .B(n_2), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_174), .B(n_3), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_146), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_143), .B(n_3), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_138), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_158), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_148), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_158), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_175), .B(n_4), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_165), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_198), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_196), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_229), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_229), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_142), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_237), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_237), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_247), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_247), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_233), .B(n_204), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_239), .A2(n_172), .B1(n_184), .B2(n_169), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_260), .B(n_165), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_237), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_263), .B(n_188), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_237), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_236), .Y(n_276) );
INVx6_ASAP7_75t_L g277 ( .A(n_259), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_243), .B(n_213), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_243), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_252), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_237), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_252), .Y(n_282) );
INVx5_ASAP7_75t_L g283 ( .A(n_254), .Y(n_283) );
INVx5_ASAP7_75t_L g284 ( .A(n_254), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_237), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_254), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_240), .Y(n_287) );
BUFx4f_ASAP7_75t_L g288 ( .A(n_259), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_244), .A2(n_231), .B1(n_216), .B2(n_220), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_262), .A2(n_153), .B1(n_179), .B2(n_157), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_244), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_234), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_259), .B(n_162), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_234), .Y(n_294) );
NAND2xp33_ASAP7_75t_L g295 ( .A(n_265), .B(n_139), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_259), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_251), .B(n_150), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_272), .B(n_245), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_288), .A2(n_257), .B(n_261), .C(n_256), .Y(n_299) );
AND2x2_ASAP7_75t_SL g300 ( .A(n_288), .B(n_250), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_287), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_297), .B(n_251), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_297), .B(n_253), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_270), .B(n_253), .Y(n_304) );
NOR2xp33_ASAP7_75t_SL g305 ( .A(n_290), .B(n_157), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_293), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_296), .B(n_258), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_291), .B(n_249), .Y(n_308) );
INVxp33_ASAP7_75t_SL g309 ( .A(n_279), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_294), .Y(n_310) );
NAND2xp33_ASAP7_75t_L g311 ( .A(n_296), .B(n_225), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_289), .A2(n_195), .B1(n_224), .B2(n_179), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_271), .B(n_155), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_274), .B(n_235), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_295), .B(n_242), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_293), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_293), .Y(n_317) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_268), .A2(n_145), .B(n_147), .C(n_144), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_277), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_277), .Y(n_320) );
OR2x6_ASAP7_75t_L g321 ( .A(n_268), .B(n_230), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_269), .B(n_160), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_276), .B(n_161), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_269), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_280), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_282), .B(n_163), .Y(n_326) );
INVx4_ASAP7_75t_L g327 ( .A(n_292), .Y(n_327) );
OR2x6_ASAP7_75t_L g328 ( .A(n_286), .B(n_228), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_283), .B(n_170), .Y(n_329) );
NOR2xp33_ASAP7_75t_SL g330 ( .A(n_283), .B(n_226), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_283), .B(n_222), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_283), .B(n_171), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_283), .B(n_187), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_284), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_284), .A2(n_254), .B1(n_255), .B2(n_248), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_266), .B(n_223), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_266), .B(n_212), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_267), .B(n_173), .Y(n_338) );
O2A1O1Ixp5_ASAP7_75t_L g339 ( .A1(n_273), .A2(n_149), .B(n_152), .C(n_151), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_273), .A2(n_254), .B1(n_255), .B2(n_248), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_275), .B(n_227), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_275), .B(n_178), .Y(n_342) );
NAND2xp33_ASAP7_75t_L g343 ( .A(n_281), .B(n_182), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_285), .B(n_156), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_303), .Y(n_345) );
BUFx12f_ASAP7_75t_L g346 ( .A(n_321), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_307), .A2(n_248), .B(n_159), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_302), .A2(n_176), .B(n_181), .C(n_167), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_324), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_307), .A2(n_248), .B(n_166), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_L g351 ( .A1(n_318), .A2(n_221), .B(n_168), .C(n_177), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_304), .B(n_183), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_308), .B(n_201), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_322), .B(n_186), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_L g355 ( .A1(n_299), .A2(n_189), .B(n_190), .C(n_185), .Y(n_355) );
O2A1O1Ixp33_ASAP7_75t_L g356 ( .A1(n_311), .A2(n_193), .B(n_202), .C(n_192), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
BUFx12f_ASAP7_75t_L g358 ( .A(n_321), .Y(n_358) );
INVxp33_ASAP7_75t_L g359 ( .A(n_305), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_325), .A2(n_207), .B(n_205), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_326), .B(n_203), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_306), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_298), .A2(n_209), .B(n_210), .C(n_208), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_316), .A2(n_194), .B1(n_255), .B2(n_211), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_298), .A2(n_215), .B1(n_218), .B2(n_214), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_319), .Y(n_366) );
BUFx12f_ASAP7_75t_L g367 ( .A(n_328), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_314), .B(n_217), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_315), .B(n_219), .Y(n_369) );
NOR3xp33_ASAP7_75t_L g370 ( .A(n_313), .B(n_197), .C(n_191), .Y(n_370) );
BUFx10_ASAP7_75t_L g371 ( .A(n_315), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g372 ( .A1(n_301), .A2(n_199), .B(n_246), .C(n_255), .Y(n_372) );
BUFx4f_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_337), .B(n_232), .Y(n_374) );
AO22x1_ASAP7_75t_L g375 ( .A1(n_332), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_375) );
O2A1O1Ixp5_ASAP7_75t_L g376 ( .A1(n_339), .A2(n_327), .B(n_341), .C(n_336), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_320), .A2(n_241), .B1(n_238), .B2(n_13), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_333), .B(n_10), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_323), .B(n_14), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_331), .B(n_14), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_340), .A2(n_241), .B(n_48), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_340), .A2(n_50), .B(n_49), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_344), .A2(n_18), .B1(n_19), .B2(n_20), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_310), .Y(n_384) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_334), .B(n_22), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_335), .A2(n_55), .B(n_52), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_338), .A2(n_342), .B(n_343), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_303), .B(n_27), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_317), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_303), .B(n_28), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_317), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_317), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_324), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_302), .B(n_29), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_324), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_324), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_324), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_302), .B(n_29), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_303), .B(n_30), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_303), .B(n_30), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_302), .B(n_32), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_305), .Y(n_402) );
AO21x1_ASAP7_75t_L g403 ( .A1(n_311), .A2(n_33), .B(n_35), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_317), .Y(n_404) );
AO22x1_ASAP7_75t_L g405 ( .A1(n_309), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_405) );
CKINVDCx10_ASAP7_75t_R g406 ( .A(n_321), .Y(n_406) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_393), .B(n_42), .Y(n_407) );
CKINVDCx6p67_ASAP7_75t_R g408 ( .A(n_406), .Y(n_408) );
AND3x1_ASAP7_75t_L g409 ( .A(n_406), .B(n_42), .C(n_43), .Y(n_409) );
BUFx12f_ASAP7_75t_L g410 ( .A(n_346), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_394), .B(n_44), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_396), .Y(n_412) );
NAND2xp33_ASAP7_75t_R g413 ( .A(n_357), .B(n_44), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_388), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_358), .Y(n_416) );
INVx4_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_349), .B(n_67), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_366), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_400), .B(n_82), .Y(n_420) );
OR2x6_ASAP7_75t_L g421 ( .A(n_348), .B(n_83), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_365), .A2(n_107), .B1(n_108), .B2(n_110), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_366), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_389), .Y(n_424) );
AO31x2_ASAP7_75t_L g425 ( .A1(n_363), .A2(n_114), .A3(n_115), .B(n_118), .Y(n_425) );
AO32x2_ASAP7_75t_L g426 ( .A1(n_377), .A2(n_119), .A3(n_122), .B1(n_123), .B2(n_124), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_352), .A2(n_374), .B(n_368), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_351), .B(n_371), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_373), .A2(n_383), .B1(n_395), .B2(n_397), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_371), .B(n_353), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_361), .A2(n_369), .B(n_354), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_370), .B(n_362), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_391), .B(n_404), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_392), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_379), .B(n_378), .Y(n_435) );
OAI22x1_ASAP7_75t_L g436 ( .A1(n_385), .A2(n_405), .B1(n_375), .B2(n_380), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_364), .A2(n_376), .B(n_350), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_384), .A2(n_288), .B(n_387), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_376), .A2(n_350), .B(n_347), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_387), .A2(n_288), .B(n_347), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_345), .B(n_309), .Y(n_441) );
AO31x2_ASAP7_75t_L g442 ( .A1(n_372), .A2(n_403), .A3(n_347), .B(n_350), .Y(n_442) );
AOI21xp33_ASAP7_75t_L g443 ( .A1(n_359), .A2(n_309), .B(n_278), .Y(n_443) );
INVx5_ASAP7_75t_L g444 ( .A(n_393), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_345), .B(n_303), .Y(n_445) );
NOR2xp67_ASAP7_75t_L g446 ( .A(n_346), .B(n_358), .Y(n_446) );
AND2x6_ASAP7_75t_L g447 ( .A(n_393), .B(n_396), .Y(n_447) );
AO31x2_ASAP7_75t_L g448 ( .A1(n_372), .A2(n_403), .A3(n_347), .B(n_350), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_345), .B(n_303), .Y(n_449) );
AO31x2_ASAP7_75t_L g450 ( .A1(n_372), .A2(n_403), .A3(n_347), .B(n_350), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_356), .A2(n_401), .B(n_398), .C(n_355), .Y(n_451) );
AO21x1_ASAP7_75t_L g452 ( .A1(n_381), .A2(n_382), .B(n_386), .Y(n_452) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_357), .B(n_330), .Y(n_453) );
OAI21x1_ASAP7_75t_SL g454 ( .A1(n_360), .A2(n_403), .B(n_356), .Y(n_454) );
AO31x2_ASAP7_75t_L g455 ( .A1(n_372), .A2(n_403), .A3(n_347), .B(n_350), .Y(n_455) );
OAI22x1_ASAP7_75t_L g456 ( .A1(n_402), .A2(n_312), .B1(n_357), .B2(n_264), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_399), .A2(n_288), .B1(n_300), .B2(n_325), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_376), .A2(n_350), .B(n_347), .Y(n_458) );
NAND2x1_ASAP7_75t_L g459 ( .A(n_447), .B(n_418), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_410), .B(n_446), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_408), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_445), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_427), .A2(n_437), .B(n_431), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_449), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_452), .A2(n_438), .B(n_451), .Y(n_465) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_444), .B(n_417), .Y(n_466) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_436), .A2(n_454), .B(n_429), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_434), .Y(n_468) );
INVx4_ASAP7_75t_L g469 ( .A(n_444), .Y(n_469) );
NOR2x1_ASAP7_75t_SL g470 ( .A(n_444), .B(n_421), .Y(n_470) );
BUFx10_ASAP7_75t_L g471 ( .A(n_416), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_414), .B(n_415), .Y(n_472) );
BUFx4f_ASAP7_75t_L g473 ( .A(n_453), .Y(n_473) );
INVx5_ASAP7_75t_L g474 ( .A(n_447), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_412), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_428), .A2(n_411), .B(n_420), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_443), .B(n_430), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_424), .Y(n_478) );
OAI21x1_ASAP7_75t_L g479 ( .A1(n_407), .A2(n_433), .B(n_422), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_432), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_456), .B(n_421), .Y(n_481) );
OAI21x1_ASAP7_75t_SL g482 ( .A1(n_426), .A2(n_413), .B(n_423), .Y(n_482) );
AO31x2_ASAP7_75t_L g483 ( .A1(n_442), .A2(n_455), .A3(n_448), .B(n_450), .Y(n_483) );
OAI21x1_ASAP7_75t_SL g484 ( .A1(n_426), .A2(n_419), .B(n_425), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_409), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_439), .A2(n_458), .B(n_440), .Y(n_486) );
AND2x6_ASAP7_75t_L g487 ( .A(n_418), .B(n_399), .Y(n_487) );
AOI21xp33_ASAP7_75t_SL g488 ( .A1(n_413), .A2(n_321), .B(n_421), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_427), .A2(n_431), .B(n_435), .C(n_451), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_445), .B(n_345), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_445), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_441), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_439), .A2(n_458), .B(n_440), .Y(n_493) );
NOR2x1_ASAP7_75t_SL g494 ( .A(n_457), .B(n_367), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_439), .A2(n_458), .B(n_440), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_445), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_468), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_466), .Y(n_498) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_484), .A2(n_465), .B(n_463), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_466), .Y(n_500) );
OAI21x1_ASAP7_75t_L g501 ( .A1(n_486), .A2(n_493), .B(n_495), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_475), .B(n_470), .Y(n_502) );
AO21x1_ASAP7_75t_SL g503 ( .A1(n_467), .A2(n_487), .B(n_481), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_460), .Y(n_504) );
NAND2x1p5_ASAP7_75t_L g505 ( .A(n_459), .B(n_474), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_478), .B(n_480), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_472), .Y(n_507) );
OR2x6_ASAP7_75t_L g508 ( .A(n_482), .B(n_476), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_483), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_462), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_487), .B(n_489), .Y(n_511) );
INVx3_ASAP7_75t_L g512 ( .A(n_469), .Y(n_512) );
NOR2x1_ASAP7_75t_SL g513 ( .A(n_469), .B(n_460), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_464), .B(n_491), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_514), .B(n_496), .Y(n_515) );
NOR2x1_ASAP7_75t_SL g516 ( .A(n_503), .B(n_460), .Y(n_516) );
INVx8_ASAP7_75t_L g517 ( .A(n_512), .Y(n_517) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_510), .A2(n_488), .B1(n_477), .B2(n_485), .C(n_492), .Y(n_518) );
INVx6_ASAP7_75t_L g519 ( .A(n_498), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_509), .B(n_494), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_497), .B(n_473), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_507), .B(n_490), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_498), .Y(n_523) );
AND2x4_ASAP7_75t_SL g524 ( .A(n_502), .B(n_471), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_511), .B(n_479), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_525), .B(n_508), .Y(n_526) );
INVx5_ASAP7_75t_L g527 ( .A(n_517), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_520), .Y(n_528) );
INVxp67_ASAP7_75t_SL g529 ( .A(n_516), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_528), .Y(n_530) );
AND3x2_ASAP7_75t_L g531 ( .A(n_529), .B(n_518), .C(n_516), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_527), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_528), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_526), .B(n_499), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_526), .B(n_501), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_528), .Y(n_536) );
INVxp33_ASAP7_75t_L g537 ( .A(n_532), .Y(n_537) );
XNOR2x1_ASAP7_75t_L g538 ( .A(n_531), .B(n_461), .Y(n_538) );
OAI31xp33_ASAP7_75t_L g539 ( .A1(n_538), .A2(n_524), .A3(n_534), .B(n_535), .Y(n_539) );
NAND3xp33_ASAP7_75t_SL g540 ( .A(n_539), .B(n_537), .C(n_504), .Y(n_540) );
OAI21xp5_ASAP7_75t_SL g541 ( .A1(n_540), .A2(n_521), .B(n_523), .Y(n_541) );
NAND4xp25_ASAP7_75t_L g542 ( .A(n_541), .B(n_521), .C(n_522), .D(n_500), .Y(n_542) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_542), .B(n_512), .Y(n_543) );
XOR2x2_ASAP7_75t_L g544 ( .A(n_543), .B(n_513), .Y(n_544) );
XNOR2xp5_ASAP7_75t_L g545 ( .A(n_544), .B(n_515), .Y(n_545) );
XNOR2xp5_ASAP7_75t_L g546 ( .A(n_545), .B(n_506), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_546), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_547), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_548), .A2(n_505), .B(n_512), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_549), .B(n_506), .Y(n_550) );
OR2x6_ASAP7_75t_L g551 ( .A(n_550), .B(n_519), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_551), .A2(n_533), .B1(n_530), .B2(n_536), .Y(n_552) );
endmodule