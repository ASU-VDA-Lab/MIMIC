module real_jpeg_32953_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_178;
wire n_67;
wire n_76;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_244;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

AND2x2_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_0),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_0),
.B(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_0),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_1),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_1),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_61),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_1),
.B(n_175),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_3),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_35),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_6),
.B(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_6),
.B(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_6),
.B(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_7),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_8),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_8),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_8),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_8),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_8),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_8),
.B(n_247),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_9),
.B(n_95),
.Y(n_94)
);

NAND2x1p5_ASAP7_75t_L g119 ( 
.A(n_9),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_9),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_10),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_10),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_10),
.B(n_211),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_10),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_11),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_13),
.Y(n_113)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_14),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_14),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_15),
.B(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_178),
.Y(n_16)
);

NAND2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_177),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp67_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_130),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_20),
.B(n_130),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_64),
.C(n_89),
.Y(n_20)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_21),
.B(n_90),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_22),
.B(n_39),
.C(n_62),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_28),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_23),
.B(n_32),
.C(n_36),
.Y(n_142)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_27),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_27),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_31),
.Y(n_168)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_38)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

MAJx2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.C(n_48),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_48),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_41),
.Y(n_218)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_42),
.Y(n_160)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_42),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_58),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_55),
.B(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_57),
.Y(n_198)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_57),
.Y(n_253)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_61),
.Y(n_239)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_65),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.C(n_85),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_66),
.B(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_70),
.B(n_85),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.C(n_82),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_71),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_74),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_75),
.A2(n_76),
.B1(n_82),
.B2(n_83),
.Y(n_222)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_77),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2x1_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_107),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_146),
.C(n_147),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_101),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_92),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_94),
.Y(n_199)
);

AO22x1_ASAP7_75t_SL g281 ( 
.A1(n_94),
.A2(n_196),
.B1(n_199),
.B2(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_95),
.Y(n_271)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_97),
.B(n_102),
.Y(n_202)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_123),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_118),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_117),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_117),
.C(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_113),
.Y(n_264)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx4f_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_126),
.B(n_129),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_126),
.Y(n_129)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_148),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_145),
.Y(n_131)
);

XOR2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_176),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_163),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_162),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_156),
.B1(n_157),
.B2(n_161),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_173),
.B2(n_174),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_203),
.B(n_292),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_181),
.B(n_183),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_200),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_201),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.C(n_195),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_191),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_192),
.B(n_239),
.Y(n_250)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_196),
.Y(n_282)
);

BUFx4f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_225),
.B(n_291),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_223),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_205),
.B(n_223),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.C(n_219),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_207),
.B(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_209),
.A2(n_220),
.B1(n_221),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_209),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.C(n_216),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_210),
.B(n_213),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_252),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_285),
.B(n_290),
.Y(n_225)
);

OAI21x1_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_273),
.B(n_284),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_254),
.B(n_272),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_240),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_231),
.A2(n_232),
.B1(n_236),
.B2(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_231),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_248),
.B2(n_249),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_246),
.C(n_248),
.Y(n_283)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_251),
.Y(n_279)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_266),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_265),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_265),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_283),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_278),
.C(n_281),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);


endmodule