module fake_jpeg_13920_n_378 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_0),
.B(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx8_ASAP7_75t_SL g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

OR2x4_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_64),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_65),
.B(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_18),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_8),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_70),
.Y(n_171)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_40),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_73),
.B(n_100),
.Y(n_175)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_16),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_79),
.Y(n_125)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_77),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_5),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_5),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_11),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_95),
.Y(n_130)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_32),
.B(n_11),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_32),
.B(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_102),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_36),
.B(n_9),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_9),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_24),
.Y(n_142)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_110),
.Y(n_124)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_108),
.B(n_109),
.Y(n_172)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_39),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_63),
.A2(n_45),
.B1(n_27),
.B2(n_52),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_115),
.A2(n_119),
.B1(n_162),
.B2(n_140),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_63),
.A2(n_45),
.B1(n_27),
.B2(n_39),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_59),
.A2(n_53),
.B(n_48),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_122),
.B(n_167),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_53),
.B(n_48),
.C(n_47),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_128),
.A2(n_134),
.A3(n_124),
.B1(n_158),
.B2(n_173),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_94),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_141),
.B(n_163),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_87),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_96),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_86),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_24),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_153),
.B(n_155),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_107),
.A2(n_61),
.B1(n_70),
.B2(n_81),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_85),
.B1(n_99),
.B2(n_56),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_69),
.B(n_30),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_69),
.B(n_30),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_157),
.B(n_164),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_73),
.A2(n_44),
.B1(n_34),
.B2(n_3),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_158),
.A2(n_138),
.B(n_115),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_66),
.A2(n_44),
.B1(n_2),
.B2(n_3),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_88),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_80),
.B(n_2),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_82),
.B(n_3),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_72),
.B(n_83),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_168),
.B(n_151),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_177),
.B(n_191),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_111),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_179),
.B(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_180),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_71),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_185),
.Y(n_233)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_92),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_184),
.B(n_193),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_172),
.Y(n_185)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_123),
.B(n_103),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_198),
.Y(n_236)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_195),
.A2(n_225),
.B1(n_191),
.B2(n_192),
.Y(n_240)
);

AOI32xp33_ASAP7_75t_L g196 ( 
.A1(n_122),
.A2(n_75),
.A3(n_125),
.B1(n_128),
.B2(n_113),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_SL g267 ( 
.A(n_196),
.B(n_224),
.C(n_227),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_150),
.A2(n_159),
.B1(n_166),
.B2(n_146),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_199),
.A2(n_195),
.B1(n_214),
.B2(n_197),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_116),
.B(n_120),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_202),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_135),
.B(n_143),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_201),
.Y(n_256)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_212),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_169),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_205),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_134),
.B(n_152),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_207),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_131),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_209),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_131),
.B(n_148),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_198),
.B(n_221),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_173),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_216),
.Y(n_253)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_119),
.A2(n_162),
.B1(n_146),
.B2(n_160),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_229),
.B1(n_114),
.B2(n_147),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_112),
.B(n_160),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_215),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_118),
.B(n_171),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_222),
.Y(n_257)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_221),
.Y(n_252)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_137),
.B(n_132),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_127),
.B(n_140),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_228),
.Y(n_242)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_127),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_144),
.B(n_151),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g239 ( 
.A(n_226),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_126),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_144),
.B(n_151),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_171),
.A2(n_114),
.B1(n_126),
.B2(n_132),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_232),
.A2(n_248),
.B1(n_262),
.B2(n_266),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_251),
.B1(n_255),
.B2(n_260),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_182),
.B1(n_186),
.B2(n_197),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_185),
.B(n_200),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_264),
.C(n_242),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_186),
.A2(n_225),
.B1(n_205),
.B2(n_196),
.Y(n_255)
);

O2A1O1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_258),
.A2(n_259),
.B(n_261),
.C(n_252),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_181),
.A2(n_199),
.B1(n_215),
.B2(n_210),
.Y(n_260)
);

OAI22x1_ASAP7_75t_SL g261 ( 
.A1(n_193),
.A2(n_184),
.B1(n_217),
.B2(n_203),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_263),
.B1(n_268),
.B2(n_259),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_184),
.A2(n_202),
.B1(n_194),
.B2(n_222),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_178),
.A2(n_230),
.B1(n_188),
.B2(n_212),
.Y(n_263)
);

AO22x1_ASAP7_75t_SL g265 ( 
.A1(n_184),
.A2(n_219),
.B1(n_180),
.B2(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_223),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_184),
.A2(n_223),
.B1(n_227),
.B2(n_183),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_187),
.A2(n_189),
.B1(n_216),
.B2(n_218),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_271),
.Y(n_316)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_269),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_224),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_276),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_220),
.Y(n_276)
);

AND2x6_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_267),
.Y(n_277)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_277),
.A2(n_296),
.A3(n_235),
.B1(n_249),
.B2(n_250),
.C1(n_256),
.C2(n_293),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_260),
.A2(n_251),
.B1(n_259),
.B2(n_231),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_278),
.A2(n_295),
.B(n_299),
.Y(n_315)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_284),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_280),
.B(n_285),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_233),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_283),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_238),
.B(n_233),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_282),
.B(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_234),
.B(n_237),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_245),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_245),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_288),
.Y(n_310)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_234),
.B(n_252),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_293),
.Y(n_317)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_248),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_294),
.C(n_281),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_292),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_258),
.A2(n_232),
.B1(n_236),
.B2(n_267),
.Y(n_293)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_265),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_253),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_298),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_256),
.B(n_241),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_246),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_274),
.A2(n_266),
.B1(n_262),
.B2(n_265),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_300),
.A2(n_286),
.B1(n_316),
.B2(n_317),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_304),
.B(n_277),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_271),
.A2(n_250),
.B(n_235),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_308),
.A2(n_312),
.B(n_314),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_309),
.B(n_320),
.Y(n_326)
);

OR2x6_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_295),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_278),
.A2(n_280),
.B(n_274),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_283),
.A2(n_275),
.B(n_276),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_289),
.C(n_272),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_306),
.B(n_285),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_321),
.B(n_323),
.Y(n_340)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_R g338 ( 
.A(n_327),
.B(n_334),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_303),
.B(n_287),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_329),
.Y(n_347)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_310),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_307),
.Y(n_330)
);

BUFx12_ASAP7_75t_L g345 ( 
.A(n_330),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_331),
.A2(n_332),
.B1(n_335),
.B2(n_319),
.Y(n_341)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

AO221x1_ASAP7_75t_L g334 ( 
.A1(n_313),
.A2(n_279),
.B1(n_288),
.B2(n_284),
.C(n_296),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_303),
.B(n_286),
.Y(n_336)
);

A2O1A1O1Ixp25_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_319),
.B(n_318),
.C(n_317),
.D(n_302),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_309),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_339),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_309),
.C(n_320),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_341),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_343),
.A2(n_312),
.B1(n_316),
.B2(n_346),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_320),
.C(n_314),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_344),
.B(n_346),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_315),
.C(n_302),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_338),
.A2(n_331),
.B1(n_329),
.B2(n_333),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_350),
.A2(n_341),
.B1(n_300),
.B2(n_312),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g351 ( 
.A1(n_347),
.A2(n_311),
.B(n_306),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_351),
.B(n_352),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_345),
.Y(n_352)
);

AOI321xp33_ASAP7_75t_L g353 ( 
.A1(n_340),
.A2(n_311),
.A3(n_332),
.B1(n_330),
.B2(n_304),
.C(n_312),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_353),
.B(n_357),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_344),
.A2(n_315),
.B(n_333),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_355),
.A2(n_312),
.B(n_308),
.Y(n_359)
);

OAI322xp33_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_347),
.A3(n_312),
.B1(n_337),
.B2(n_339),
.C1(n_338),
.C2(n_335),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_358),
.A2(n_359),
.B(n_312),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_363),
.Y(n_369)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_301),
.C(n_345),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_354),
.Y(n_367)
);

NAND4xp25_ASAP7_75t_SL g365 ( 
.A(n_360),
.B(n_345),
.C(n_364),
.D(n_343),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_365),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_362),
.B(n_342),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_366),
.A2(n_367),
.B(n_368),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_361),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_371),
.B(n_356),
.C(n_301),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_372),
.A2(n_366),
.B(n_356),
.C(n_348),
.Y(n_373)
);

OAI21x1_ASAP7_75t_SL g375 ( 
.A1(n_373),
.A2(n_359),
.B(n_348),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_374),
.B(n_370),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_375),
.B(n_376),
.C(n_322),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_325),
.Y(n_378)
);


endmodule