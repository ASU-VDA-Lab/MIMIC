module real_jpeg_30916_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_0),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_0),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_468),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_1),
.B(n_469),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_2),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_2),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_3),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_3),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_4),
.Y(n_398)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_5),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_5),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_6),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_7),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_8),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_8),
.A2(n_146),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_L g352 ( 
.A1(n_8),
.A2(n_146),
.B1(n_205),
.B2(n_353),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_8),
.A2(n_146),
.B1(n_426),
.B2(n_428),
.Y(n_425)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22x1_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_10),
.A2(n_29),
.B1(n_88),
.B2(n_92),
.Y(n_87)
);

AO22x2_ASAP7_75t_SL g130 ( 
.A1(n_10),
.A2(n_29),
.B1(n_131),
.B2(n_135),
.Y(n_130)
);

OAI22x1_ASAP7_75t_SL g216 ( 
.A1(n_10),
.A2(n_29),
.B1(n_217),
.B2(n_220),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_11),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_11),
.A2(n_61),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_11),
.A2(n_61),
.B1(n_231),
.B2(n_235),
.Y(n_230)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_12),
.A2(n_73),
.B1(n_76),
.B2(n_78),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_12),
.Y(n_78)
);

AOI22x1_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_78),
.B1(n_98),
.B2(n_102),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_12),
.A2(n_78),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g367 ( 
.A(n_12),
.B(n_368),
.Y(n_367)
);

OAI32xp33_ASAP7_75t_L g392 ( 
.A1(n_12),
.A2(n_393),
.A3(n_399),
.B1(n_401),
.B2(n_405),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_12),
.B(n_129),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_13),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_256),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_254),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_224),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_19),
.B(n_224),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_179),
.C(n_187),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_21),
.B(n_179),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_94),
.Y(n_21)
);

INVxp33_ASAP7_75t_SL g252 ( 
.A(n_22),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_54),
.B(n_67),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_23),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_23),
.B(n_54),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_23),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

AO22x2_ASAP7_75t_L g184 ( 
.A1(n_24),
.A2(n_35),
.B1(n_55),
.B2(n_66),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_24),
.B(n_66),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_27),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_28),
.Y(n_360)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_34),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_35),
.B(n_203),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_35),
.A2(n_66),
.B(n_203),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_35),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_45),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_42),
.Y(n_413)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_44),
.Y(n_369)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_49),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_49),
.Y(n_404)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_66),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_66),
.B(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_66),
.B(n_352),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g441 ( 
.A(n_66),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_67),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_79),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_68),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AO21x2_ASAP7_75t_L g181 ( 
.A1(n_70),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_72),
.B(n_80),
.Y(n_336)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21x1_ASAP7_75t_SL g170 ( 
.A1(n_78),
.A2(n_171),
.B(n_175),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_78),
.B(n_176),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_78),
.B(n_178),
.Y(n_334)
);

AOI32xp33_ASAP7_75t_L g357 ( 
.A1(n_78),
.A2(n_358),
.A3(n_361),
.B1(n_366),
.B2(n_367),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_78),
.B(n_402),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_78),
.B(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_78),
.B(n_81),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_79),
.A2(n_191),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_79),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_87),
.Y(n_79)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_80),
.B(n_425),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_87),
.B(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_91),
.Y(n_193)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_139),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_95),
.Y(n_253)
);

NOR2x1p5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_128),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_96),
.Y(n_383)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_105),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_97),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_97),
.Y(n_290)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_101),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_104),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_105),
.Y(n_241)
);

AO21x2_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_113),
.B(n_121),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_106),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_121)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_122),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_128),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_129),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_129),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_129),
.B(n_292),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_130),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_133),
.Y(n_272)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_133),
.Y(n_294)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp33_ASAP7_75t_SL g251 ( 
.A(n_139),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_169),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_140),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_151),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_141),
.B(n_161),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_145),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_145),
.Y(n_280)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_151),
.B(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_151),
.A2(n_170),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_151),
.B(n_170),
.Y(n_321)
);

NOR2x1p5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_161),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_159),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_156),
.Y(n_276)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_156),
.Y(n_285)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

AO22x2_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_175),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_177),
.B(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_181),
.A2(n_185),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_SL g356 ( 
.A(n_181),
.B(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_181),
.A2(n_185),
.B1(n_357),
.B2(n_380),
.Y(n_379)
);

OAI21xp33_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_191),
.B(n_197),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_185),
.Y(n_249)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_188),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_210),
.C(n_214),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_189),
.B(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_201),
.Y(n_189)
);

XOR2x2_ASAP7_75t_L g322 ( 
.A(n_190),
.B(n_201),
.Y(n_322)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_193),
.Y(n_427)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_197),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_SL g442 ( 
.A(n_197),
.B(n_424),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_198),
.Y(n_268)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_202),
.B(n_386),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_207),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_208),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_209),
.B(n_351),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_211),
.B(n_214),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_223),
.B(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_250),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_244),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_242),
.Y(n_226)
);

NAND2x1_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_238),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_236),
.A2(n_282),
.B(n_286),
.Y(n_281)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_240),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_243),
.B(n_351),
.Y(n_350)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.C(n_253),
.Y(n_250)
);

INVxp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21x1_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_307),
.B(n_467),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_305),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_259),
.B(n_305),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.C(n_302),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_260),
.A2(n_261),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_265),
.B(n_303),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_287),
.C(n_299),
.Y(n_265)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_267),
.B(n_269),
.Y(n_330)
);

OAI31xp33_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_273),
.A3(n_277),
.B(n_281),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_287),
.A2(n_288),
.B1(n_300),
.B2(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_339),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_343),
.B(n_461),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_326),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_310),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_323),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_311),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.C(n_322),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

XOR2x1_ASAP7_75t_SL g342 ( 
.A(n_316),
.B(n_322),
.Y(n_342)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.C(n_320),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_383),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_329),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_323),
.Y(n_466)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_341),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_327),
.B(n_341),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.C(n_331),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_371),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_332),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_338),
.B(n_340),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_333),
.A2(n_334),
.B(n_335),
.Y(n_349)
);

NOR2x1_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_SL g340 ( 
.A(n_334),
.B(n_335),
.Y(n_340)
);

NOR2x1p5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_336),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_349),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_372),
.B(n_460),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_370),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_346),
.B(n_370),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.C(n_356),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_348),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_356),
.Y(n_376)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx6f_ASAP7_75t_SL g368 ( 
.A(n_369),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_387),
.B(n_459),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_377),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_374),
.B(n_377),
.Y(n_459)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.C(n_384),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_379),
.B(n_455),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_381),
.A2(n_382),
.B1(n_384),
.B2(n_385),
.Y(n_455)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_453),
.B(n_458),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_389),
.A2(n_431),
.B(n_452),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_416),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_390),
.B(n_416),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_414),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_391),
.A2(n_392),
.B1(n_414),
.B2(n_415),
.Y(n_437)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_398),
.Y(n_430)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_422),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_423),
.C(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_421),
.Y(n_457)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AOI21x1_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_438),
.B(n_451),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_437),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_437),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_445),
.Y(n_444)
);

BUFx4f_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_443),
.B(n_450),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_442),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_442),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_446),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_449),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_454),
.B(n_456),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);


endmodule