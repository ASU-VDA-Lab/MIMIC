module real_jpeg_12076_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_1),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_1),
.A2(n_29),
.B1(n_33),
.B2(n_46),
.Y(n_156)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_5),
.A2(n_74),
.B1(n_75),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_5),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_5),
.A2(n_73),
.B(n_74),
.C(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_5),
.B(n_84),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_145),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_5),
.A2(n_102),
.B1(n_103),
.B2(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_5),
.B(n_90),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_6),
.A2(n_74),
.B1(n_75),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_6),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_147),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_147),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_6),
.A2(n_29),
.B1(n_33),
.B2(n_147),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_10),
.A2(n_74),
.B1(n_75),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_10),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_135),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_135),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_10),
.A2(n_29),
.B1(n_33),
.B2(n_135),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_11),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_11),
.A2(n_29),
.B1(n_33),
.B2(n_55),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_12),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_12),
.A2(n_37),
.B1(n_61),
.B2(n_62),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_12),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_12),
.A2(n_37),
.B1(n_74),
.B2(n_75),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_13),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_13),
.A2(n_32),
.B1(n_74),
.B2(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_13),
.A2(n_32),
.B1(n_61),
.B2(n_62),
.Y(n_131)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_15),
.A2(n_74),
.B1(n_75),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_82),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_15),
.A2(n_43),
.B1(n_44),
.B2(n_82),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_15),
.A2(n_29),
.B1(n_33),
.B2(n_82),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_138),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_19),
.B(n_116),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_86),
.B2(n_115),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.C(n_69),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_22),
.A2(n_23),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_26),
.A2(n_102),
.B(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_27),
.A2(n_38),
.B1(n_126),
.B2(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_27),
.A2(n_38),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_28),
.A2(n_38),
.B(n_128),
.Y(n_197)
);

CKINVDCx6p67_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_29),
.A2(n_33),
.B1(n_49),
.B2(n_50),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_33),
.B(n_50),
.C(n_145),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_33),
.B(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_34),
.A2(n_103),
.B(n_156),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_36),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_42),
.A2(n_52),
.B(n_95),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g193 ( 
.A1(n_43),
.A2(n_58),
.B(n_194),
.C(n_196),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_43),
.B(n_216),
.Y(n_215)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

NOR3xp33_ASAP7_75t_L g196 ( 
.A(n_44),
.B(n_59),
.C(n_61),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_47),
.A2(n_54),
.B(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_47),
.A2(n_94),
.B(n_107),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_47),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_47),
.A2(n_53),
.B1(n_201),
.B2(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_47),
.A2(n_53),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_47),
.A2(n_53),
.B1(n_209),
.B2(n_219),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_52),
.B(n_145),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_69),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_64),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_68),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_57),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_66)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_62),
.B1(n_73),
.B2(n_78),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_61),
.A2(n_78),
.B(n_145),
.Y(n_158)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g195 ( 
.A(n_62),
.B(n_145),
.CON(n_195),
.SN(n_195)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_65),
.A2(n_90),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_65),
.A2(n_90),
.B1(n_167),
.B2(n_195),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_80),
.B(n_83),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_70),
.A2(n_79),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_71),
.A2(n_81),
.B1(n_84),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_71),
.A2(n_84),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_72)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_99),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B(n_98),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_90),
.B(n_131),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_93),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_108),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_102),
.A2(n_103),
.B1(n_224),
.B2(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_103),
.B(n_145),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_122),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_121),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_122),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.C(n_133),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_123),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_129),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_130),
.B(n_133),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_268),
.B(n_273),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_185),
.B(n_259),
.C(n_267),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_170),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_141),
.B(n_170),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_153),
.C(n_161),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_142),
.B(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_149),
.C(n_152),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_153),
.B(n_161),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_159),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.C(n_165),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_165),
.B(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_179),
.B(n_180),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_182),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_171),
.B(n_183),
.C(n_184),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_181),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_175),
.B(n_178),
.C(n_181),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_254),
.B(n_258),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_210),
.B(n_253),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_205),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_205),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_202),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_192),
.B(n_198),
.C(n_202),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_197),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.C(n_208),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_208),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_248),
.B(n_252),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_238),
.B(n_247),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_227),
.B(n_237),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_222),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_220),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_236),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_235),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_240),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_243),
.C(n_246),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_266),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_263),
.C(n_264),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);


endmodule