module real_jpeg_21498_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_249;
wire n_286;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_150;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_0),
.A2(n_66),
.B1(n_67),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_0),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_0),
.A2(n_28),
.B1(n_37),
.B2(n_111),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_111),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_111),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_1),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_1),
.B(n_72),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_1),
.A2(n_16),
.B(n_45),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_136),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_81),
.B1(n_82),
.B2(n_194),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_1),
.B(n_59),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_1),
.A2(n_37),
.B(n_225),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_66),
.B1(n_67),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_2),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_90),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_2),
.A2(n_28),
.B1(n_37),
.B2(n_90),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_90),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_3),
.A2(n_36),
.B1(n_66),
.B2(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_3),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_4),
.A2(n_66),
.B1(n_67),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_4),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_4),
.A2(n_28),
.B1(n_37),
.B2(n_138),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_138),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_138),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_5),
.A2(n_28),
.B1(n_37),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_5),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_132),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_132),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_132),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_6),
.A2(n_28),
.B1(n_37),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_6),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_122)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_8),
.A2(n_28),
.B1(n_37),
.B2(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_101)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_13),
.A2(n_28),
.B1(n_37),
.B2(n_65),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_65),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_65),
.Y(n_169)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_14),
.A2(n_33),
.A3(n_37),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_16),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_16),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_91),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_91),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_78),
.B2(n_79),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_51),
.B2(n_52),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_25),
.A2(n_26),
.B(n_40),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_26)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_27),
.A2(n_31),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_27),
.A2(n_31),
.B1(n_133),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_27),
.A2(n_31),
.B1(n_164),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_27),
.A2(n_31),
.B1(n_107),
.B2(n_146),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.Y(n_30)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_28),
.A2(n_37),
.B1(n_70),
.B2(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_28),
.A2(n_71),
.B1(n_135),
.B2(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_28),
.B(n_136),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_29),
.B(n_32),
.Y(n_220)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_33),
.A2(n_43),
.B(n_136),
.C(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_35),
.A2(n_57),
.B1(n_59),
.B2(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_37),
.B(n_70),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_44),
.B(n_49),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_41),
.A2(n_44),
.B1(n_47),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_41),
.A2(n_44),
.B1(n_86),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_41),
.A2(n_44),
.B1(n_104),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_41),
.A2(n_44),
.B1(n_124),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_41),
.A2(n_44),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_41),
.A2(n_44),
.B1(n_190),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_41),
.A2(n_44),
.B1(n_210),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_41),
.A2(n_44),
.B1(n_128),
.B2(n_228),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_44),
.B(n_136),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_46),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_62),
.B1(n_76),
.B2(n_77),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_57),
.A2(n_59),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_68),
.B1(n_74),
.B2(n_75),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_69),
.B1(n_72),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_66),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_70),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_66),
.B(n_136),
.CON(n_135),
.SN(n_135)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_75),
.B1(n_89),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_68),
.A2(n_75),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_68),
.A2(n_75),
.B1(n_110),
.B2(n_144),
.Y(n_266)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_69),
.A2(n_72),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_84),
.B(n_87),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_87),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_80),
.A2(n_85),
.B1(n_95),
.B2(n_281),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_83),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_81),
.A2(n_82),
.B1(n_101),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_81),
.A2(n_122),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_81),
.A2(n_82),
.B1(n_152),
.B2(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_81),
.A2(n_153),
.B1(n_180),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_81),
.A2(n_82),
.B1(n_182),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_81),
.A2(n_82),
.B1(n_169),
.B2(n_212),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_82),
.B(n_136),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_85),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_97),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_92),
.B(n_96),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_97),
.A2(n_98),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.C(n_108),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_99),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_100),
.B(n_103),
.Y(n_260)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_105),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_284),
.B(n_289),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_271),
.B(n_283),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_170),
.B(n_253),
.C(n_270),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_155),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_118),
.B(n_155),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_139),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_120),
.B(n_125),
.C(n_139),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_121),
.B(n_123),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_134),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_137),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_148),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_147),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_141),
.B(n_147),
.C(n_148),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_145),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_151),
.Y(n_159)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_178),
.B1(n_179),
.B2(n_181),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_156),
.B(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_167),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_162),
.B(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_166),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_252),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_247),
.B(n_251),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_233),
.B(n_246),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_214),
.B(n_232),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_202),
.B(n_213),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_191),
.B(n_201),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_183),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_183),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_187),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_196),
.B(n_200),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_195),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_204),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_211),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_209),
.C(n_211),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_216),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_222),
.B1(n_230),
.B2(n_231),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_217),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_219),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_221),
.Y(n_225)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_226),
.B1(n_227),
.B2(n_229),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_223),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_234),
.B(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_240),
.B2(n_241),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_243),
.C(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_243),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_249),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_254),
.B(n_255),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_269),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_262),
.C(n_269),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_265),
.C(n_268),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_273),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_282),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_280),
.C(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);


endmodule