module fake_jpeg_90_n_525 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_14),
.B(n_13),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_51),
.B(n_89),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_52),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_31),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_88),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_55),
.Y(n_138)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_72),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_34),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_1),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_39),
.Y(n_88)
);

BUFx12f_ASAP7_75t_SL g89 ( 
.A(n_39),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_96),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

BUFx4f_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_97),
.B(n_96),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_99),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_36),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_38),
.B1(n_20),
.B2(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_109),
.A2(n_112),
.B1(n_124),
.B2(n_137),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_38),
.B1(n_47),
.B2(n_34),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_126),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_118),
.A2(n_44),
.B(n_40),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_80),
.A2(n_38),
.B1(n_47),
.B2(n_43),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_42),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_127),
.B(n_131),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_63),
.B(n_36),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_85),
.A2(n_28),
.B1(n_25),
.B2(n_33),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_55),
.A2(n_33),
.B1(n_28),
.B2(n_46),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_139),
.A2(n_86),
.B1(n_87),
.B2(n_91),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_54),
.B(n_2),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_74),
.B(n_2),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_48),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_66),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_97),
.B(n_46),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_95),
.B(n_46),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_70),
.Y(n_185)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_162),
.Y(n_240)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_164),
.Y(n_214)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_167),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_157),
.A2(n_112),
.B1(n_118),
.B2(n_115),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_197),
.B1(n_125),
.B2(n_128),
.Y(n_210)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_192),
.Y(n_221)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_157),
.A2(n_107),
.B1(n_148),
.B2(n_146),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_176),
.A2(n_199),
.B1(n_205),
.B2(n_207),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_64),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_190),
.Y(n_211)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_21),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_194),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_150),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_195),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_196),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_244)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_198),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_146),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

O2A1O1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_124),
.A2(n_44),
.B(n_24),
.C(n_17),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_151),
.B(n_161),
.Y(n_219)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_132),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_132),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_121),
.Y(n_228)
);

CKINVDCx6p67_ASAP7_75t_R g207 ( 
.A(n_137),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_148),
.A2(n_84),
.B1(n_82),
.B2(n_79),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_209),
.B1(n_161),
.B2(n_145),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_168),
.B1(n_183),
.B2(n_212),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_101),
.C(n_105),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_201),
.C(n_180),
.Y(n_259)
);

OA22x2_ASAP7_75t_SL g218 ( 
.A1(n_207),
.A2(n_130),
.B1(n_158),
.B2(n_151),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_218),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_219),
.A2(n_203),
.B1(n_194),
.B2(n_182),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_228),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_123),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_238),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_138),
.B1(n_155),
.B2(n_149),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_188),
.B1(n_133),
.B2(n_142),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_184),
.B(n_114),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_247),
.A2(n_260),
.B1(n_268),
.B2(n_273),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_207),
.B1(n_170),
.B2(n_164),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_248),
.A2(n_262),
.B1(n_213),
.B2(n_243),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_175),
.C(n_179),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_272),
.C(n_243),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_242),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_172),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_265),
.Y(n_282)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_SL g280 ( 
.A1(n_256),
.A2(n_248),
.B(n_257),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_163),
.B(n_172),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_266),
.B(n_218),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_165),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_233),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_228),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_264),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_214),
.A2(n_166),
.B1(n_178),
.B2(n_200),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_SL g264 ( 
.A1(n_230),
.A2(n_178),
.B(n_181),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_122),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_219),
.A2(n_177),
.B(n_209),
.Y(n_266)
);

OR2x2_ASAP7_75t_SL g267 ( 
.A(n_218),
.B(n_167),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_267),
.A2(n_213),
.B(n_223),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_210),
.A2(n_102),
.B1(n_133),
.B2(n_142),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_229),
.B(n_169),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_271),
.Y(n_283)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_270),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_221),
.B(n_173),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_221),
.B(n_186),
.C(n_204),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_231),
.A2(n_102),
.B1(n_160),
.B2(n_154),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_227),
.B(n_193),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_236),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_280),
.A2(n_250),
.B(n_261),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_274),
.Y(n_281)
);

BUFx4f_ASAP7_75t_SL g334 ( 
.A(n_281),
.Y(n_334)
);

OAI21xp33_ASAP7_75t_SL g284 ( 
.A1(n_256),
.A2(n_218),
.B(n_244),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_288),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_285),
.A2(n_294),
.B(n_304),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_258),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_247),
.A2(n_240),
.B1(n_224),
.B2(n_227),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_290),
.B1(n_268),
.B2(n_272),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_224),
.B1(n_240),
.B2(n_246),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_305),
.B1(n_270),
.B2(n_263),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_266),
.A2(n_276),
.B(n_253),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_306),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_296),
.A2(n_261),
.B(n_267),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_249),
.B(n_224),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_299),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_249),
.B(n_235),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_261),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_309),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_266),
.A2(n_216),
.B(n_237),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_264),
.A2(n_246),
.B1(n_237),
.B2(n_216),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_233),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_226),
.C(n_232),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_250),
.A2(n_222),
.B1(n_236),
.B2(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_294),
.A2(n_300),
.B1(n_285),
.B2(n_302),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_313),
.A2(n_316),
.B1(n_324),
.B2(n_331),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_326),
.B(n_337),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_300),
.A2(n_262),
.B1(n_267),
.B2(n_250),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_307),
.Y(n_318)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_321),
.A2(n_291),
.B1(n_289),
.B2(n_278),
.Y(n_343)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_323),
.A2(n_336),
.B(n_326),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_292),
.A2(n_299),
.B1(n_281),
.B2(n_288),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_251),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_332),
.Y(n_349)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_327),
.Y(n_353)
);

A2O1A1O1Ixp25_ASAP7_75t_L g328 ( 
.A1(n_292),
.A2(n_269),
.B(n_259),
.C(n_265),
.D(n_272),
.Y(n_328)
);

OAI211xp5_ASAP7_75t_L g374 ( 
.A1(n_328),
.A2(n_341),
.B(n_192),
.C(n_234),
.Y(n_374)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_303),
.Y(n_329)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_279),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_330),
.B(n_308),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_292),
.A2(n_305),
.B1(n_282),
.B2(n_280),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_275),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_297),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_292),
.A2(n_255),
.B(n_254),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_298),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_279),
.A2(n_260),
.B1(n_273),
.B2(n_217),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_340),
.A2(n_198),
.B1(n_222),
.B2(n_239),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_290),
.A2(n_222),
.B1(n_195),
.B2(n_189),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_295),
.C(n_308),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_343),
.A2(n_350),
.B1(n_355),
.B2(n_363),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_327),
.A2(n_304),
.B1(n_309),
.B2(n_282),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_345),
.A2(n_368),
.B1(n_373),
.B2(n_331),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_334),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_346),
.B(n_352),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_372),
.C(n_319),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_348),
.A2(n_371),
.B(n_374),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_313),
.A2(n_284),
.B1(n_283),
.B2(n_295),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_312),
.B(n_283),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_310),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_316),
.A2(n_296),
.B1(n_286),
.B2(n_309),
.Y(n_355)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_226),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_375),
.Y(n_388)
);

OA21x2_ASAP7_75t_L g361 ( 
.A1(n_315),
.A2(n_234),
.B(n_239),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_339),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_217),
.Y(n_366)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_366),
.Y(n_389)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_315),
.A2(n_217),
.B1(n_160),
.B2(n_154),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_317),
.B(n_202),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_369),
.B(n_323),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_232),
.Y(n_370)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_342),
.C(n_332),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_315),
.A2(n_239),
.B1(n_155),
.B2(n_149),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_324),
.B(n_199),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_377),
.A2(n_385),
.B1(n_392),
.B2(n_400),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_386),
.C(n_375),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_320),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_381),
.B(n_393),
.Y(n_409)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_384),
.B(n_401),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_310),
.B1(n_337),
.B2(n_320),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_372),
.C(n_359),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_314),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_395),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_370),
.Y(n_391)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_391),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_353),
.A2(n_337),
.B1(n_336),
.B2(n_329),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_328),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_341),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_343),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_344),
.B(n_322),
.Y(n_395)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_344),
.B(n_225),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_373),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_225),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_399),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_366),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_348),
.B(n_196),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_225),
.Y(n_402)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_402),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_355),
.A2(n_205),
.B1(n_76),
.B2(n_78),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_404),
.A2(n_356),
.B1(n_77),
.B2(n_73),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_145),
.Y(n_405)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_418),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_379),
.A2(n_371),
.B(n_361),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_413),
.A2(n_424),
.B(n_394),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_386),
.B(n_361),
.C(n_345),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_419),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_421),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_377),
.A2(n_351),
.B1(n_367),
.B2(n_358),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_422),
.A2(n_404),
.B1(n_380),
.B2(n_69),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_379),
.A2(n_368),
.B(n_358),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_378),
.B(n_351),
.C(n_364),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_431),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_362),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_401),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_356),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_376),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_395),
.Y(n_429)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_429),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_430),
.A2(n_65),
.B1(n_60),
.B2(n_24),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_396),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_435),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_388),
.C(n_390),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_439),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_407),
.B(n_426),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_434),
.B(n_443),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_413),
.A2(n_392),
.B(n_385),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_436),
.A2(n_442),
.B(n_414),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_415),
.Y(n_437)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_437),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_388),
.C(n_397),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_441),
.B(n_410),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_389),
.B(n_398),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_389),
.C(n_384),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_398),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_444),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_446),
.A2(n_430),
.B1(n_445),
.B2(n_424),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_416),
.B(n_2),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_449),
.B(n_2),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_409),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_SL g454 ( 
.A(n_450),
.B(n_453),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_452),
.A2(n_419),
.B1(n_422),
.B2(n_414),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_35),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_450),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_420),
.C(n_421),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_466),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_458),
.A2(n_460),
.B1(n_462),
.B2(n_463),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_412),
.Y(n_459)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_459),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_442),
.A2(n_423),
.B1(n_411),
.B2(n_406),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_406),
.C(n_44),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_447),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_468),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_451),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_446),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_433),
.B(n_2),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_471),
.B(n_470),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_436),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_472),
.A2(n_453),
.B1(n_4),
.B2(n_5),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_460),
.A2(n_432),
.B(n_440),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_473),
.A2(n_488),
.B(n_5),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_477),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_463),
.A2(n_443),
.B(n_444),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_480),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_457),
.B(n_435),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_466),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_440),
.C(n_441),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_484),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_459),
.A2(n_461),
.B(n_456),
.Y(n_480)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_481),
.Y(n_491)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_482),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_3),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_4),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_489),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_462),
.A2(n_4),
.B(n_5),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_35),
.C(n_6),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_6),
.C(n_7),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_458),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_493),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_480),
.B(n_486),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_487),
.B(n_454),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_499),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_479),
.B(n_472),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_501),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_474),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_482),
.Y(n_508)
);

NOR2x1_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_497),
.Y(n_505)
);

NAND3xp33_ASAP7_75t_SL g514 ( 
.A(n_505),
.B(n_510),
.C(n_501),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_474),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_507),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_494),
.A2(n_476),
.B(n_478),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_508),
.B(n_509),
.Y(n_516)
);

OAI321xp33_ASAP7_75t_L g509 ( 
.A1(n_494),
.A2(n_481),
.A3(n_473),
.B1(n_488),
.B2(n_489),
.C(n_35),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_503),
.A2(n_490),
.B(n_500),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_SL g518 ( 
.A(n_512),
.B(n_514),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_504),
.B(n_498),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_515),
.B(n_517),
.C(n_7),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_502),
.C(n_35),
.Y(n_517)
);

AOI321xp33_ASAP7_75t_L g519 ( 
.A1(n_513),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_519),
.A2(n_8),
.B(n_12),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_520),
.A2(n_516),
.B1(n_10),
.B2(n_11),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_521),
.A2(n_522),
.B(n_518),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g524 ( 
.A(n_523),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_12),
.Y(n_525)
);


endmodule