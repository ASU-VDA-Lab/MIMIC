module fake_jpeg_27322_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_55),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_25),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_28),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_39),
.B2(n_38),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_72),
.B1(n_17),
.B2(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_16),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_29),
.Y(n_69)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_88),
.B1(n_89),
.B2(n_94),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_41),
.C(n_46),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_90),
.C(n_109),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_39),
.B1(n_38),
.B2(n_42),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_98),
.B1(n_64),
.B2(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_101),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_45),
.B1(n_36),
.B2(n_43),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_84),
.A2(n_64),
.B1(n_74),
.B2(n_54),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_87),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g87 ( 
.A(n_48),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_23),
.B1(n_27),
.B2(n_32),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_19),
.B1(n_34),
.B2(n_33),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_43),
.C(n_45),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_91),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_49),
.A2(n_23),
.B1(n_27),
.B2(n_32),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_47),
.A2(n_17),
.B1(n_21),
.B2(n_26),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_111),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_54),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_104),
.A2(n_61),
.B1(n_55),
.B2(n_60),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_30),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_43),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_49),
.A2(n_45),
.B1(n_36),
.B2(n_34),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_51),
.A2(n_30),
.B1(n_33),
.B2(n_31),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_113),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_48),
.B(n_36),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_126),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_128),
.B1(n_106),
.B2(n_103),
.Y(n_154)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_105),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_90),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_80),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_131),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_30),
.C(n_33),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_99),
.C(n_109),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_137),
.B1(n_140),
.B2(n_113),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_95),
.A2(n_74),
.B(n_34),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_111),
.B(n_86),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_31),
.B1(n_24),
.B2(n_19),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_31),
.B1(n_24),
.B2(n_19),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_143),
.Y(n_166)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_144),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_105),
.B(n_95),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_164),
.B(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_146),
.B(n_150),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_152),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_155),
.B1(n_168),
.B2(n_5),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_83),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_172),
.B(n_5),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_75),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_102),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_159),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_156),
.B1(n_160),
.B2(n_167),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_120),
.B1(n_123),
.B2(n_138),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_111),
.B1(n_84),
.B2(n_81),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_109),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_120),
.B1(n_135),
.B2(n_139),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_161),
.B(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_111),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_120),
.A2(n_113),
.B(n_82),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_175),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_139),
.B1(n_132),
.B2(n_141),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_110),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_96),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_143),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_93),
.B1(n_106),
.B2(n_24),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_91),
.B(n_2),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_116),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_130),
.B1(n_126),
.B2(n_8),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_116),
.B(n_5),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_142),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_7),
.Y(n_195)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_180),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_192),
.B1(n_200),
.B2(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_187),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_159),
.C(n_153),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_201),
.C(n_149),
.Y(n_220)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_7),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_7),
.Y(n_199)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_8),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_10),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_171),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_12),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_13),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_209),
.B(n_219),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_214),
.B1(n_221),
.B2(n_225),
.Y(n_241)
);

AOI22x1_ASAP7_75t_SL g213 ( 
.A1(n_207),
.A2(n_151),
.B1(n_167),
.B2(n_168),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_213),
.A2(n_228),
.B1(n_198),
.B2(n_193),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_148),
.B1(n_145),
.B2(n_144),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_224),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_180),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_172),
.B1(n_164),
.B2(n_161),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_179),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_183),
.B(n_182),
.C(n_184),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_173),
.B(n_176),
.C(n_15),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_232),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_190),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_225),
.B1(n_181),
.B2(n_186),
.Y(n_247)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_191),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_191),
.B(n_182),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_226),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_226),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_217),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_187),
.Y(n_242)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_189),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_229),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_255),
.B1(n_224),
.B2(n_208),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_248),
.A2(n_251),
.B1(n_254),
.B2(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_201),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_215),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_252),
.B(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_198),
.B1(n_208),
.B2(n_223),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_256),
.A2(n_245),
.B1(n_234),
.B2(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_210),
.C(n_233),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_261),
.C(n_272),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_220),
.C(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_249),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_211),
.C(n_222),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_227),
.C(n_249),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_279),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_260),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_240),
.B1(n_236),
.B2(n_235),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_282),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_268),
.Y(n_298)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_284),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_243),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_286),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_254),
.B(n_269),
.C(n_259),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_267),
.B(n_265),
.Y(n_296)
);

INVx11_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_272),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_298),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_275),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_300),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_285),
.C(n_261),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_287),
.B(n_270),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_305),
.B(n_290),
.Y(n_309)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_287),
.B(n_282),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_298),
.B(n_296),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_287),
.B(n_262),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_303),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_309),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_289),
.B(n_291),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_312),
.B1(n_293),
.B2(n_291),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_310),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_294),
.C(n_301),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_317),
.Y(n_318)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_306),
.B(n_314),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_262),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_257),
.Y(n_321)
);


endmodule