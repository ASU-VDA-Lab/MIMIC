module fake_netlist_6_806_n_2180 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2180);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2180;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_162),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_101),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_115),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_11),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_118),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_41),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_117),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_97),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_85),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_110),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_98),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_50),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_119),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_179),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_10),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_132),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_32),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_40),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_129),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_45),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_124),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_76),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_51),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_37),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_42),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_5),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_33),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_57),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_15),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_214),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_100),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_193),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_194),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_174),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_113),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_71),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_186),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_9),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_172),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_107),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_63),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_196),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_161),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_24),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_158),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_15),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_91),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_136),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_165),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_182),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_84),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_89),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_66),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_75),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_190),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_45),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_133),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_63),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_8),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_178),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_173),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_57),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_140),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_68),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_163),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_92),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_90),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_35),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_77),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_183),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_58),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_42),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_147),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_82),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_87),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_41),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_34),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_58),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_65),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_37),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_134),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_112),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_111),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_105),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_122),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_114),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_71),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_167),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_192),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_146),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_171),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_52),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_99),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_39),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_130),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_185),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_120),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_102),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_166),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_187),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_80),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_2),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_141),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_152),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_26),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_189),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_128),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_75),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_34),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_143),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_198),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_24),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_177),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_126),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_212),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_176),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_72),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_44),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_144),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_10),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_66),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_9),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_205),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_145),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_199),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_1),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_70),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_67),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_17),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_27),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_78),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_31),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_195),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_206),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_28),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_46),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_209),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_61),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_46),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_109),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_86),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_121),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_6),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_26),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_74),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_169),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_44),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_11),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_211),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_153),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_188),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_139),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_65),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_61),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_123),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_48),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_81),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_88),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_215),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_43),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_40),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_25),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_168),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_68),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_52),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_135),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_28),
.Y(n_387)
);

BUFx2_ASAP7_75t_SL g388 ( 
.A(n_20),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_48),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_148),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_150),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_191),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_204),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_0),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_43),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_104),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_72),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_216),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_149),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_49),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_156),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_8),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_47),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_64),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_95),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_125),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_33),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_106),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_94),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_18),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_23),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_54),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_67),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_69),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_55),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_55),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_7),
.Y(n_417)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_180),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_0),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_137),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_2),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_56),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_5),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_6),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_108),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_12),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_31),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_223),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_325),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_232),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_325),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_382),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_382),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_266),
.B(n_1),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_240),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_382),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_279),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_296),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_249),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_281),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_322),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_311),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_348),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_264),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_283),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_220),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_264),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_337),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_302),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_353),
.B(n_305),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_344),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_410),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_299),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_327),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_267),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_410),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_414),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_269),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_3),
.Y(n_463)
);

BUFx6f_ASAP7_75t_SL g464 ( 
.A(n_310),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_310),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_273),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_271),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_276),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_305),
.B(n_3),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_282),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_278),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_304),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_291),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_220),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_274),
.B(n_4),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_272),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_222),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_287),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_289),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_292),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_297),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_299),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_290),
.B(n_4),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_244),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_307),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_222),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_328),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_329),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_290),
.B(n_7),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_350),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_301),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_356),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_363),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_389),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_298),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_391),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_394),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_300),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_312),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_303),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_299),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_244),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_341),
.B(n_12),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_314),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_332),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_338),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_L g510 ( 
.A(n_338),
.B(n_13),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_226),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_306),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_371),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_342),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_374),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_226),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_346),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_374),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_400),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_308),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_404),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_313),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_347),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_315),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_419),
.B(n_13),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_316),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_391),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_424),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_218),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_326),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_340),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_317),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_374),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_326),
.B(n_333),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_340),
.B(n_14),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_349),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_454),
.B(n_217),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_513),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_513),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_513),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_432),
.B(n_333),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_513),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_446),
.B(n_217),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_433),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_531),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_433),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_434),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_513),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_463),
.B(n_339),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_438),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_536),
.A2(n_474),
.B(n_449),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_432),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_474),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_438),
.B(n_339),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_449),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_430),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_484),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_453),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_468),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_456),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_456),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_460),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_466),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_477),
.B(n_380),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_532),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_467),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_486),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_532),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_463),
.B(n_370),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_532),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_439),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_486),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_450),
.B(n_370),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_505),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_498),
.B(n_409),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_471),
.B(n_219),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_505),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_509),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_509),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_533),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_533),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_531),
.B(n_409),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_485),
.B(n_491),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_487),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_489),
.Y(n_592)
);

BUFx8_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_510),
.B(n_371),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_490),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_492),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_465),
.B(n_368),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_494),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_465),
.B(n_368),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_495),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_496),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_499),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_529),
.B(n_219),
.Y(n_603)
);

INVx6_ASAP7_75t_L g604 ( 
.A(n_529),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_468),
.B(n_470),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_504),
.B(n_371),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_519),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_448),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_521),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_522),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_428),
.A2(n_427),
.B1(n_242),
.B2(n_284),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_526),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_470),
.B(n_401),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_530),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_429),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_431),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_435),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_436),
.B(n_371),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_461),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_537),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_451),
.B(n_221),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_435),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_473),
.B(n_221),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_506),
.B(n_371),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_440),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_451),
.B(n_225),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_572),
.Y(n_627)
);

BUFx4f_ASAP7_75t_L g628 ( 
.A(n_554),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_572),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_572),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_590),
.B(n_444),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_572),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_604),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_547),
.B(n_224),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_558),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_541),
.Y(n_636)
);

INVx6_ASAP7_75t_L g637 ( 
.A(n_604),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_543),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_543),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_558),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_554),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_575),
.B(n_420),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_543),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_543),
.Y(n_644)
);

INVx6_ASAP7_75t_L g645 ( 
.A(n_604),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_613),
.B(n_458),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_541),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_613),
.B(n_430),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_623),
.B(n_535),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_617),
.B(n_473),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_558),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_590),
.B(n_459),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_541),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_539),
.B(n_462),
.Y(n_654)
);

AND2x2_ASAP7_75t_SL g655 ( 
.A(n_554),
.B(n_420),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_539),
.B(n_469),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_547),
.B(n_227),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_558),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_561),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_570),
.A2(n_352),
.B1(n_402),
.B2(n_288),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_608),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_559),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_623),
.B(n_478),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_617),
.B(n_475),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_543),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_617),
.B(n_476),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_617),
.A2(n_575),
.B1(n_552),
.B2(n_579),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_621),
.B(n_479),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_559),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_559),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_582),
.B(n_480),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_543),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_608),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_595),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_617),
.B(n_604),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_604),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_559),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_604),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_563),
.Y(n_679)
);

AND2x2_ASAP7_75t_SL g680 ( 
.A(n_554),
.B(n_420),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_575),
.B(n_475),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_595),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_618),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_563),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_564),
.B(n_482),
.Y(n_685)
);

OR2x6_ASAP7_75t_L g686 ( 
.A(n_604),
.B(n_527),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_564),
.B(n_482),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_621),
.B(n_488),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_605),
.B(n_483),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_541),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_563),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_603),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_541),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_605),
.B(n_483),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_541),
.Y(n_695)
);

OR2x6_ASAP7_75t_L g696 ( 
.A(n_603),
.B(n_570),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_626),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_626),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_575),
.A2(n_527),
.B1(n_387),
.B2(n_403),
.Y(n_699)
);

INVx11_ASAP7_75t_L g700 ( 
.A(n_593),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_545),
.B(n_497),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_541),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_545),
.B(n_497),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_595),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_579),
.B(n_388),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_575),
.B(n_500),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_563),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_575),
.B(n_500),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_595),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_552),
.B(n_501),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_547),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_552),
.B(n_501),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_595),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_565),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_565),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_565),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_565),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_579),
.B(n_507),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_541),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_561),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_560),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_567),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_581),
.A2(n_387),
.B1(n_403),
.B2(n_373),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_560),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_556),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_567),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_571),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_581),
.B(n_507),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_596),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_596),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_582),
.B(n_481),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_581),
.B(n_511),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_567),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_567),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_568),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_596),
.Y(n_736)
);

INVxp33_ASAP7_75t_L g737 ( 
.A(n_611),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_593),
.B(n_508),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_568),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_622),
.B(n_538),
.Y(n_740)
);

AND2x6_ASAP7_75t_L g741 ( 
.A(n_624),
.B(n_420),
.Y(n_741)
);

AND2x6_ASAP7_75t_L g742 ( 
.A(n_624),
.B(n_420),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_596),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_547),
.B(n_493),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_624),
.B(n_508),
.Y(n_745)
);

BUFx10_ASAP7_75t_L g746 ( 
.A(n_622),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_589),
.B(n_239),
.C(n_228),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_597),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_554),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_624),
.B(n_514),
.Y(n_750)
);

BUFx6f_ASAP7_75t_SL g751 ( 
.A(n_624),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_620),
.B(n_373),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_554),
.A2(n_421),
.B1(n_445),
.B2(n_516),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_596),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_589),
.B(n_514),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_597),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_597),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_611),
.B(n_503),
.C(n_457),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_593),
.B(n_517),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_612),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_624),
.A2(n_421),
.B1(n_321),
.B2(n_425),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_568),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_599),
.B(n_268),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_568),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_599),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_546),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_599),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_612),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_556),
.Y(n_769)
);

OR2x6_ASAP7_75t_L g770 ( 
.A(n_616),
.B(n_270),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_612),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_540),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_546),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_546),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_612),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_589),
.B(n_275),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_616),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_R g778 ( 
.A(n_562),
.B(n_577),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_551),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_612),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_551),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_675),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_746),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_692),
.A2(n_594),
.B1(n_557),
.B2(n_592),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_692),
.B(n_594),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_667),
.B(n_594),
.Y(n_786)
);

OAI221xp5_ASAP7_75t_L g787 ( 
.A1(n_699),
.A2(n_619),
.B1(n_588),
.B2(n_600),
.C(n_601),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_652),
.B(n_631),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_721),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_766),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_697),
.B(n_594),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_698),
.B(n_594),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_661),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_655),
.B(n_593),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_696),
.A2(n_512),
.B1(n_520),
.B2(n_502),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_655),
.B(n_680),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_765),
.B(n_592),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_766),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_748),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_655),
.B(n_593),
.Y(n_800)
);

OAI22xp33_ASAP7_75t_L g801 ( 
.A1(n_696),
.A2(n_577),
.B1(n_625),
.B2(n_562),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_671),
.B(n_523),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_680),
.B(n_592),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_748),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_680),
.B(n_592),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_SL g806 ( 
.A(n_660),
.B(n_441),
.C(n_437),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_675),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_650),
.B(n_664),
.Y(n_808)
);

INVxp33_ASAP7_75t_L g809 ( 
.A(n_661),
.Y(n_809)
);

NAND2x1_ASAP7_75t_L g810 ( 
.A(n_675),
.B(n_637),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_666),
.B(n_619),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_628),
.B(n_593),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_696),
.A2(n_528),
.B1(n_534),
.B2(n_525),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_731),
.B(n_654),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_773),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_642),
.B(n_304),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_773),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_774),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_628),
.B(n_562),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_656),
.B(n_625),
.C(n_577),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_628),
.B(n_625),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_666),
.B(n_615),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_756),
.B(n_592),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_756),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_757),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_675),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_757),
.A2(n_557),
.B1(n_609),
.B2(n_592),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_767),
.B(n_592),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_641),
.B(n_304),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_767),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_638),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_774),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_779),
.Y(n_833)
);

AOI221xp5_ASAP7_75t_L g834 ( 
.A1(n_737),
.A2(n_238),
.B1(n_397),
.B2(n_229),
.C(n_365),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_711),
.B(n_609),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_638),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_641),
.B(n_304),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_639),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_779),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_781),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_639),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_643),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_644),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_641),
.B(n_304),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_749),
.B(n_304),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_749),
.B(n_304),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_711),
.B(n_609),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_749),
.B(n_304),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_705),
.B(n_620),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_696),
.B(n_609),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_665),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_665),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_777),
.B(n_615),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_732),
.B(n_615),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_L g855 ( 
.A(n_646),
.B(n_524),
.C(n_517),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_777),
.B(n_615),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_781),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_696),
.B(n_609),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_672),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_681),
.B(n_418),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_689),
.B(n_440),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_753),
.A2(n_447),
.B1(n_452),
.B2(n_442),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_672),
.B(n_609),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_694),
.B(n_443),
.Y(n_864)
);

NOR2x1p5_ASAP7_75t_L g865 ( 
.A(n_721),
.B(n_724),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_674),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_776),
.A2(n_557),
.B1(n_609),
.B2(n_280),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_706),
.A2(n_455),
.B1(n_538),
.B2(n_524),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_718),
.B(n_609),
.Y(n_869)
);

AO21x1_ASAP7_75t_L g870 ( 
.A1(n_776),
.A2(n_285),
.B(n_277),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_674),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_728),
.B(n_557),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_708),
.B(n_557),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_701),
.A2(n_703),
.B1(n_750),
.B2(n_745),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_776),
.B(n_556),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_648),
.B(n_443),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_732),
.B(n_588),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_776),
.B(n_710),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_673),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_635),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_723),
.A2(n_607),
.B(n_601),
.C(n_600),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_712),
.B(n_556),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_682),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_772),
.B(n_556),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_668),
.B(n_515),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_682),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_704),
.Y(n_887)
);

BUFx10_ASAP7_75t_L g888 ( 
.A(n_663),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_725),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_740),
.B(n_518),
.C(n_607),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_755),
.B(n_746),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_634),
.B(n_548),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_668),
.B(n_464),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_688),
.B(n_418),
.Y(n_894)
);

AND2x2_ASAP7_75t_SL g895 ( 
.A(n_758),
.B(n_286),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_634),
.B(n_548),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_704),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_634),
.B(n_549),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_635),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_634),
.B(n_549),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_640),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_640),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_651),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_651),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_658),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_658),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_688),
.B(n_649),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_709),
.B(n_418),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_709),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_642),
.A2(n_379),
.B1(n_294),
.B2(n_295),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_657),
.B(n_553),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_657),
.B(n_553),
.Y(n_912)
);

AND2x6_ASAP7_75t_SL g913 ( 
.A(n_744),
.B(n_293),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_657),
.B(n_566),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_675),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_755),
.B(n_591),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_657),
.B(n_566),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_713),
.B(n_729),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_713),
.B(n_574),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_746),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_705),
.B(n_591),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_729),
.B(n_730),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_662),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_705),
.A2(n_318),
.B1(n_319),
.B2(n_324),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_685),
.B(n_464),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_730),
.B(n_574),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_736),
.B(n_743),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_705),
.A2(n_331),
.B1(n_334),
.B2(n_336),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_736),
.B(n_574),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_687),
.B(n_225),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_705),
.B(n_591),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_673),
.B(n_235),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_L g933 ( 
.A(n_659),
.B(n_376),
.C(n_355),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_743),
.B(n_574),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_754),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_754),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_760),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_686),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_760),
.B(n_574),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_727),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_686),
.A2(n_396),
.B1(n_377),
.B2(n_369),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_778),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_768),
.B(n_551),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_768),
.B(n_576),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_771),
.B(n_418),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_662),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_720),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_771),
.B(n_576),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_686),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_775),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_669),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_790),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_814),
.A2(n_763),
.B1(n_686),
.B2(n_642),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_790),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_788),
.B(n_686),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_796),
.A2(n_676),
.B(n_633),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_891),
.B(n_659),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_796),
.A2(n_780),
.B(n_775),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_808),
.A2(n_660),
.B1(n_761),
.B2(n_763),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_822),
.B(n_763),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_786),
.A2(n_763),
.B1(n_642),
.B2(n_747),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_793),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_803),
.A2(n_676),
.B(n_633),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_822),
.B(n_763),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_819),
.A2(n_752),
.B(n_747),
.C(n_738),
.Y(n_965)
);

AO21x1_ASAP7_75t_L g966 ( 
.A1(n_850),
.A2(n_780),
.B(n_320),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_878),
.A2(n_759),
.B(n_769),
.C(n_725),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_916),
.A2(n_642),
.B1(n_770),
.B2(n_751),
.Y(n_968)
);

NAND2xp33_ASAP7_75t_L g969 ( 
.A(n_782),
.B(n_724),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_782),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_SL g971 ( 
.A1(n_829),
.A2(n_323),
.B(n_330),
.C(n_309),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_916),
.B(n_725),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_891),
.B(n_769),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_854),
.B(n_769),
.Y(n_974)
);

NOR3xp33_ASAP7_75t_L g975 ( 
.A(n_802),
.B(n_231),
.C(n_230),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_819),
.A2(n_752),
.B(n_770),
.C(n_343),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_854),
.B(n_752),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_885),
.B(n_752),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_798),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_805),
.A2(n_678),
.B(n_690),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_829),
.A2(n_678),
.B(n_670),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_932),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_785),
.B(n_770),
.Y(n_983)
);

AO22x1_ASAP7_75t_L g984 ( 
.A1(n_930),
.A2(n_257),
.B1(n_255),
.B2(n_248),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_831),
.Y(n_985)
);

OAI21xp33_ASAP7_75t_L g986 ( 
.A1(n_834),
.A2(n_236),
.B(n_235),
.Y(n_986)
);

AND2x2_ASAP7_75t_SL g987 ( 
.A(n_947),
.B(n_335),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_907),
.A2(n_241),
.B(n_236),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_869),
.A2(n_693),
.B(n_690),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_872),
.B(n_770),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_798),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_783),
.B(n_573),
.Y(n_992)
);

BUFx5_ASAP7_75t_L g993 ( 
.A(n_866),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_810),
.A2(n_693),
.B(n_690),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_811),
.B(n_770),
.Y(n_995)
);

NAND3xp33_ASAP7_75t_SL g996 ( 
.A(n_820),
.B(n_243),
.C(n_241),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_783),
.B(n_230),
.Y(n_997)
);

AOI21xp33_ASAP7_75t_L g998 ( 
.A1(n_861),
.A2(n_384),
.B(n_381),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_811),
.B(n_636),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_836),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_815),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_821),
.A2(n_614),
.B(n_591),
.C(n_598),
.Y(n_1002)
);

INVx5_ASAP7_75t_L g1003 ( 
.A(n_782),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_873),
.A2(n_647),
.B(n_636),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_877),
.B(n_380),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_791),
.B(n_636),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_920),
.B(n_231),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_807),
.A2(n_751),
.B1(n_700),
.B2(n_645),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_837),
.A2(n_653),
.B(n_647),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_932),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_789),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_837),
.A2(n_653),
.B(n_647),
.Y(n_1012)
);

O2A1O1Ixp5_ASAP7_75t_L g1013 ( 
.A1(n_860),
.A2(n_695),
.B(n_702),
.C(n_653),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_821),
.A2(n_614),
.B(n_610),
.C(n_598),
.Y(n_1014)
);

AND2x6_ASAP7_75t_L g1015 ( 
.A(n_807),
.B(n_727),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_942),
.B(n_751),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_815),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_838),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_920),
.B(n_233),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_SL g1020 ( 
.A(n_789),
.B(n_233),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_792),
.B(n_695),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_844),
.A2(n_702),
.B(n_695),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_844),
.A2(n_719),
.B(n_702),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_877),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_882),
.B(n_719),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_782),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_807),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_826),
.A2(n_700),
.B1(n_637),
.B2(n_645),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_845),
.A2(n_719),
.B(n_629),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_809),
.B(n_888),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_826),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_826),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_845),
.A2(n_848),
.B(n_846),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_841),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_799),
.B(n_642),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_809),
.B(n_234),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_915),
.A2(n_645),
.B1(n_637),
.B2(n_251),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_846),
.A2(n_670),
.B(n_669),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_848),
.A2(n_629),
.B(n_627),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_915),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_915),
.A2(n_637),
.B1(n_645),
.B2(n_234),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_817),
.Y(n_1042)
);

AOI21x1_ASAP7_75t_L g1043 ( 
.A1(n_927),
.A2(n_679),
.B(n_677),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_874),
.B(n_237),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_879),
.B(n_237),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_894),
.A2(n_598),
.B(n_602),
.C(n_610),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_860),
.A2(n_679),
.B(n_677),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_823),
.A2(n_828),
.B(n_875),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_842),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_804),
.B(n_642),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_927),
.A2(n_691),
.B(n_684),
.Y(n_1051)
);

AND2x2_ASAP7_75t_SL g1052 ( 
.A(n_895),
.B(n_380),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_801),
.B(n_250),
.Y(n_1053)
);

AO21x1_ASAP7_75t_L g1054 ( 
.A1(n_858),
.A2(n_630),
.B(n_627),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_797),
.A2(n_632),
.B(n_630),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_824),
.B(n_727),
.Y(n_1056)
);

BUFx12f_ASAP7_75t_L g1057 ( 
.A(n_865),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_888),
.B(n_250),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_843),
.A2(n_632),
.B(n_602),
.C(n_610),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_888),
.B(n_251),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_894),
.A2(n_598),
.B(n_602),
.C(n_610),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_825),
.B(n_727),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_817),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_863),
.A2(n_691),
.B(n_684),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_864),
.B(n_876),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_884),
.A2(n_714),
.B(n_707),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_830),
.B(n_727),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_851),
.A2(n_602),
.B(n_614),
.C(n_739),
.Y(n_1068)
);

BUFx8_ASAP7_75t_L g1069 ( 
.A(n_921),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_892),
.A2(n_714),
.B(n_707),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_896),
.A2(n_716),
.B(n_715),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_938),
.B(n_252),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_898),
.A2(n_716),
.B(n_715),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_818),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_853),
.Y(n_1075)
);

AND2x6_ASAP7_75t_SL g1076 ( 
.A(n_925),
.B(n_573),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_938),
.B(n_683),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_900),
.A2(n_764),
.B(n_722),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_949),
.B(n_252),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_911),
.A2(n_722),
.B(n_717),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_852),
.A2(n_859),
.B(n_931),
.C(n_921),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_853),
.B(n_690),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_881),
.A2(n_614),
.B(n_762),
.C(n_726),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_835),
.A2(n_693),
.B(n_683),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_853),
.B(n_693),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_856),
.B(n_693),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_871),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_847),
.A2(n_683),
.B(n_717),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_L g1089 ( 
.A(n_949),
.B(n_741),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_856),
.B(n_726),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_918),
.A2(n_734),
.B(n_733),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_889),
.A2(n_683),
.B(n_733),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_856),
.B(n_735),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_849),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_912),
.A2(n_683),
.B(n_735),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_931),
.B(n_739),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_784),
.B(n_762),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_870),
.A2(n_742),
.B1(n_741),
.B2(n_418),
.Y(n_1098)
);

NOR2x1_ASAP7_75t_L g1099 ( 
.A(n_890),
.B(n_764),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_914),
.A2(n_917),
.B(n_922),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_827),
.A2(n_571),
.B(n_540),
.Y(n_1101)
);

OAI321xp33_ASAP7_75t_L g1102 ( 
.A1(n_806),
.A2(n_586),
.A3(n_585),
.B1(n_587),
.B2(n_576),
.C(n_255),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_940),
.A2(n_571),
.B(n_540),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_883),
.B(n_741),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_886),
.A2(n_741),
.B(n_742),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_895),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_868),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_887),
.B(n_741),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_897),
.B(n_741),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_940),
.A2(n_571),
.B(n_540),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_909),
.B(n_741),
.Y(n_1111)
);

NOR2x1p5_ASAP7_75t_L g1112 ( 
.A(n_913),
.B(n_243),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_935),
.B(n_742),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_818),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_936),
.A2(n_742),
.B(n_542),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_940),
.A2(n_571),
.B(n_540),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_919),
.A2(n_542),
.B(n_550),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_926),
.A2(n_542),
.B(n_550),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_937),
.A2(n_742),
.B(n_542),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_929),
.A2(n_939),
.B(n_934),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_950),
.B(n_742),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_893),
.A2(n_366),
.B(n_375),
.C(n_372),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_862),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_832),
.B(n_833),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_944),
.A2(n_544),
.B(n_550),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_849),
.Y(n_1126)
);

OAI321xp33_ASAP7_75t_L g1127 ( 
.A1(n_787),
.A2(n_585),
.A3(n_587),
.B1(n_586),
.B2(n_247),
.C(n_246),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_794),
.A2(n_366),
.B1(n_253),
.B2(n_254),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_832),
.B(n_742),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_849),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_795),
.B(n_253),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_833),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_948),
.A2(n_544),
.B(n_550),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_813),
.B(n_254),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_908),
.A2(n_544),
.B(n_571),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_839),
.B(n_569),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_849),
.B(n_256),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_839),
.B(n_569),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_840),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_840),
.B(n_569),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_857),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_881),
.A2(n_569),
.B(n_555),
.C(n_544),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1100),
.A2(n_800),
.B(n_794),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1033),
.A2(n_800),
.B(n_812),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1123),
.A2(n_867),
.B1(n_812),
.B2(n_941),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1065),
.B(n_1107),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_982),
.B(n_855),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1003),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1033),
.A2(n_1048),
.B(n_955),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1026),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1011),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_959),
.A2(n_924),
.B1(n_928),
.B2(n_857),
.Y(n_1152)
);

AOI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1131),
.A2(n_943),
.B(n_908),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_985),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1000),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_L g1156 ( 
.A(n_1057),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1048),
.A2(n_816),
.B(n_945),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1018),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1010),
.B(n_933),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_962),
.B(n_880),
.Y(n_1160)
);

NOR2xp67_ASAP7_75t_L g1161 ( 
.A(n_1106),
.B(n_945),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_L g1162 ( 
.A(n_998),
.B(n_407),
.C(n_385),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1043),
.A2(n_899),
.B(n_880),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_978),
.A2(n_870),
.B1(n_816),
.B2(n_351),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1024),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_994),
.A2(n_951),
.B(n_946),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1120),
.A2(n_1039),
.B(n_1013),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1005),
.B(n_411),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1075),
.B(n_899),
.Y(n_1169)
);

AND2x6_ASAP7_75t_L g1170 ( 
.A(n_1026),
.B(n_901),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1034),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1058),
.B(n_901),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1060),
.B(n_902),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1030),
.B(n_902),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1141),
.Y(n_1175)
);

NOR2x1_ASAP7_75t_R g1176 ( 
.A(n_1134),
.B(n_245),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1049),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_980),
.A2(n_951),
.B(n_946),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1026),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_R g1180 ( 
.A(n_969),
.B(n_996),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_975),
.B(n_412),
.C(n_413),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_957),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_SL g1183 ( 
.A(n_1052),
.B(n_256),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_953),
.A2(n_910),
.B1(n_923),
.B2(n_906),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1053),
.A2(n_923),
.B(n_906),
.C(n_905),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1094),
.B(n_903),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1044),
.A2(n_905),
.B(n_904),
.C(n_903),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1141),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_987),
.B(n_245),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1122),
.A2(n_904),
.B(n_569),
.C(n_555),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_961),
.A2(n_426),
.B1(n_359),
.B2(n_358),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1036),
.B(n_988),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1087),
.B(n_258),
.Y(n_1193)
);

NAND2xp33_ASAP7_75t_R g1194 ( 
.A(n_970),
.B(n_1016),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1069),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_L g1196 ( 
.A(n_984),
.B(n_364),
.C(n_426),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_974),
.B(n_258),
.Y(n_1197)
);

O2A1O1Ixp5_ASAP7_75t_L g1198 ( 
.A1(n_966),
.A2(n_555),
.B(n_418),
.C(n_383),
.Y(n_1198)
);

BUFx4f_ASAP7_75t_L g1199 ( 
.A(n_1130),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_965),
.A2(n_362),
.B(n_372),
.C(n_361),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_952),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_977),
.B(n_259),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_995),
.A2(n_1081),
.B(n_976),
.C(n_990),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_972),
.A2(n_571),
.B(n_345),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_SL g1205 ( 
.A(n_1003),
.B(n_259),
.Y(n_1205)
);

BUFx2_ASAP7_75t_SL g1206 ( 
.A(n_1003),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1069),
.Y(n_1207)
);

CKINVDCx11_ASAP7_75t_R g1208 ( 
.A(n_1076),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_960),
.A2(n_262),
.B1(n_261),
.B2(n_265),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_989),
.A2(n_571),
.B(n_354),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_958),
.A2(n_555),
.B(n_390),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1020),
.B(n_246),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_970),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_964),
.A2(n_378),
.B1(n_392),
.B2(n_393),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_999),
.B(n_261),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1003),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1102),
.A2(n_257),
.B(n_248),
.C(n_247),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1045),
.B(n_260),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_997),
.B(n_260),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1082),
.A2(n_399),
.B(n_357),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1075),
.B(n_992),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1075),
.B(n_262),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1085),
.A2(n_405),
.B(n_386),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1128),
.A2(n_263),
.B(n_358),
.C(n_359),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1127),
.A2(n_263),
.B(n_364),
.C(n_367),
.Y(n_1225)
);

OAI22x1_ASAP7_75t_L g1226 ( 
.A1(n_1112),
.A2(n_423),
.B1(n_422),
.B2(n_417),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_1137),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1027),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_954),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1007),
.B(n_367),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_973),
.B(n_265),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1027),
.B(n_360),
.Y(n_1232)
);

INVxp67_ASAP7_75t_L g1233 ( 
.A(n_1137),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1027),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1130),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1031),
.A2(n_360),
.B1(n_362),
.B2(n_375),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1040),
.B(n_361),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_986),
.B(n_417),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1040),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1130),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1019),
.B(n_422),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_968),
.A2(n_423),
.B1(n_406),
.B2(n_408),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1097),
.A2(n_398),
.B1(n_578),
.B2(n_580),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1072),
.B(n_578),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1096),
.B(n_578),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1086),
.A2(n_578),
.B(n_584),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1079),
.B(n_578),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_979),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1031),
.B(n_578),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1002),
.A2(n_1014),
.B(n_1119),
.C(n_1115),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1126),
.A2(n_418),
.B1(n_584),
.B2(n_583),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1040),
.B(n_418),
.Y(n_1252)
);

OR2x4_ASAP7_75t_L g1253 ( 
.A(n_1056),
.B(n_578),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_983),
.A2(n_578),
.B(n_580),
.C(n_583),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1032),
.B(n_14),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1006),
.A2(n_580),
.B(n_584),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1032),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_1008),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_967),
.A2(n_580),
.B1(n_583),
.B2(n_584),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_993),
.B(n_1021),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1099),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1120),
.A2(n_618),
.B(n_606),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_991),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1001),
.B(n_79),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_971),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1090),
.A2(n_580),
.B1(n_583),
.B2(n_584),
.Y(n_1266)
);

AO32x1_ASAP7_75t_L g1267 ( 
.A1(n_1037),
.A2(n_16),
.A3(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1017),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1093),
.A2(n_1124),
.B1(n_1074),
.B2(n_1139),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1015),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1015),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1083),
.A2(n_1004),
.B(n_1046),
.C(n_1061),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_993),
.B(n_580),
.Y(n_1273)
);

AND2x2_ASAP7_75t_SL g1274 ( 
.A(n_1098),
.B(n_19),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1062),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1089),
.A2(n_580),
.B(n_584),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1015),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_993),
.B(n_580),
.Y(n_1278)
);

O2A1O1Ixp5_ASAP7_75t_L g1279 ( 
.A1(n_1054),
.A2(n_103),
.B(n_116),
.C(n_96),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_993),
.A2(n_584),
.B1(n_583),
.B2(n_618),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1042),
.A2(n_583),
.B1(n_584),
.B2(n_25),
.Y(n_1281)
);

CKINVDCx6p67_ASAP7_75t_R g1282 ( 
.A(n_1015),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1025),
.A2(n_583),
.B(n_93),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1063),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1114),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_993),
.B(n_583),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_993),
.B(n_22),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1132),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1035),
.B(n_83),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1067),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_963),
.A2(n_127),
.B(n_213),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1136),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1050),
.B(n_22),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_963),
.A2(n_956),
.B(n_1004),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1138),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1015),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1104),
.B(n_23),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1140),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1077),
.B(n_131),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1077),
.B(n_210),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1041),
.A2(n_618),
.B1(n_606),
.B2(n_30),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1108),
.B(n_208),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1012),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1068),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1109),
.B(n_29),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_981),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1129),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1066),
.B(n_32),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1163),
.A2(n_1055),
.B(n_1039),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1227),
.B(n_1059),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1182),
.B(n_1111),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1235),
.Y(n_1312)
);

BUFx4f_ASAP7_75t_L g1313 ( 
.A(n_1240),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1182),
.B(n_1113),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_SL g1315 ( 
.A1(n_1203),
.A2(n_1121),
.B(n_1028),
.C(n_1105),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1154),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1150),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1149),
.A2(n_956),
.B(n_1091),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1146),
.B(n_1047),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1218),
.B(n_1172),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1150),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1160),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1183),
.A2(n_1095),
.B1(n_1080),
.B2(n_1078),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_SL g1324 ( 
.A(n_1183),
.B(n_1080),
.C(n_1070),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1294),
.A2(n_1055),
.B(n_1029),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1173),
.B(n_1071),
.Y(n_1326)
);

O2A1O1Ixp5_ASAP7_75t_SL g1327 ( 
.A1(n_1259),
.A2(n_1038),
.B(n_1051),
.C(n_1142),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1178),
.A2(n_1029),
.B(n_1064),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1166),
.A2(n_1157),
.B(n_1167),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1155),
.Y(n_1330)
);

AO22x1_ASAP7_75t_L g1331 ( 
.A1(n_1212),
.A2(n_618),
.B1(n_606),
.B2(n_38),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1158),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1168),
.B(n_1135),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1143),
.A2(n_1066),
.B(n_1078),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1174),
.B(n_1073),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1165),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1189),
.B(n_1135),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1171),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1147),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1199),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1159),
.A2(n_1071),
.B1(n_1073),
.B2(n_1070),
.Y(n_1341)
);

NAND2x1p5_ASAP7_75t_L g1342 ( 
.A(n_1199),
.B(n_1148),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1177),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1144),
.A2(n_1009),
.B(n_1022),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1151),
.Y(n_1345)
);

AOI21xp33_ASAP7_75t_L g1346 ( 
.A1(n_1192),
.A2(n_1009),
.B(n_1022),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1224),
.A2(n_1133),
.B(n_1125),
.C(n_1118),
.Y(n_1347)
);

AOI221x1_ASAP7_75t_L g1348 ( 
.A1(n_1200),
.A2(n_1133),
.B1(n_1023),
.B2(n_1117),
.C(n_1118),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1167),
.A2(n_1023),
.B(n_1117),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1201),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1257),
.Y(n_1351)
);

A2O1A1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1219),
.A2(n_1230),
.B(n_1241),
.C(n_1153),
.Y(n_1352)
);

CKINVDCx9p33_ASAP7_75t_R g1353 ( 
.A(n_1253),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1254),
.A2(n_1101),
.A3(n_1092),
.B(n_1088),
.Y(n_1354)
);

AOI21x1_ASAP7_75t_SL g1355 ( 
.A1(n_1308),
.A2(n_1084),
.B(n_1110),
.Y(n_1355)
);

BUFx12f_ASAP7_75t_L g1356 ( 
.A(n_1208),
.Y(n_1356)
);

O2A1O1Ixp5_ASAP7_75t_SL g1357 ( 
.A1(n_1259),
.A2(n_1116),
.B(n_1103),
.C(n_38),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1207),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1246),
.A2(n_142),
.B(n_207),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1162),
.A2(n_35),
.B(n_36),
.C(n_39),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1196),
.A2(n_36),
.B(n_47),
.C(n_49),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1275),
.B(n_1268),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1150),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1269),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1165),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1145),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_1366)
);

A2O1A1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1145),
.A2(n_1152),
.B(n_1164),
.C(n_1181),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1233),
.B(n_155),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1217),
.B(n_53),
.C(n_56),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1260),
.A2(n_159),
.B(n_202),
.Y(n_1370)
);

BUFx2_ASAP7_75t_R g1371 ( 
.A(n_1206),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1258),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1269),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1225),
.A2(n_59),
.B(n_60),
.C(n_62),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1148),
.B(n_160),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_SL g1376 ( 
.A1(n_1304),
.A2(n_164),
.B(n_200),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1232),
.A2(n_618),
.B1(n_606),
.B2(n_70),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1152),
.B(n_64),
.C(n_69),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1272),
.A2(n_170),
.B(n_197),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1237),
.A2(n_618),
.B1(n_606),
.B2(n_73),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1238),
.B(n_73),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1250),
.A2(n_1245),
.B(n_1278),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_SL g1383 ( 
.A1(n_1302),
.A2(n_175),
.B(n_138),
.C(n_151),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_1176),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1273),
.A2(n_154),
.B(n_157),
.Y(n_1385)
);

AO31x2_ASAP7_75t_L g1386 ( 
.A1(n_1243),
.A2(n_618),
.A3(n_606),
.B(n_74),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1286),
.A2(n_181),
.B(n_184),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1256),
.A2(n_618),
.B(n_606),
.Y(n_1388)
);

O2A1O1Ixp5_ASAP7_75t_SL g1389 ( 
.A1(n_1243),
.A2(n_606),
.B(n_618),
.C(n_1281),
.Y(n_1389)
);

AOI221xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1191),
.A2(n_606),
.B1(n_618),
.B2(n_1242),
.C(n_1209),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1229),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1271),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1274),
.A2(n_606),
.B1(n_1186),
.B2(n_1242),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1161),
.A2(n_606),
.B(n_1293),
.C(n_1305),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1179),
.Y(n_1395)
);

AO21x1_ASAP7_75t_L g1396 ( 
.A1(n_1287),
.A2(n_1297),
.B(n_1255),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1303),
.A2(n_1202),
.B(n_1279),
.C(n_1261),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1306),
.A2(n_1276),
.B(n_1249),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1205),
.A2(n_1184),
.B(n_1283),
.Y(n_1399)
);

AO32x2_ASAP7_75t_L g1400 ( 
.A1(n_1281),
.A2(n_1191),
.A3(n_1184),
.B1(n_1266),
.B2(n_1267),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1193),
.B(n_1222),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1248),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1156),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1186),
.A2(n_1180),
.B1(n_1264),
.B2(n_1231),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1190),
.A2(n_1290),
.B(n_1185),
.C(n_1198),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1263),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1187),
.A2(n_1307),
.B(n_1262),
.Y(n_1407)
);

AO32x2_ASAP7_75t_L g1408 ( 
.A1(n_1266),
.A2(n_1267),
.A3(n_1236),
.B1(n_1296),
.B2(n_1284),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1307),
.A2(n_1262),
.B(n_1210),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1197),
.A2(n_1215),
.B(n_1204),
.Y(n_1410)
);

AOI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1226),
.A2(n_1265),
.B1(n_1301),
.B2(n_1195),
.C(n_1291),
.Y(n_1411)
);

AOI221xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1275),
.A2(n_1223),
.B1(n_1220),
.B2(n_1285),
.C(n_1288),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1239),
.Y(n_1413)
);

AO31x2_ASAP7_75t_L g1414 ( 
.A1(n_1292),
.A2(n_1298),
.A3(n_1295),
.B(n_1211),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1289),
.A2(n_1252),
.B(n_1169),
.Y(n_1415)
);

NOR2xp67_ASAP7_75t_R g1416 ( 
.A(n_1270),
.B(n_1277),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1211),
.A2(n_1216),
.B(n_1221),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1234),
.B(n_1228),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1282),
.A2(n_1253),
.B1(n_1277),
.B2(n_1264),
.Y(n_1419)
);

AO32x2_ASAP7_75t_L g1420 ( 
.A1(n_1267),
.A2(n_1194),
.A3(n_1205),
.B1(n_1170),
.B2(n_1299),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1214),
.B(n_1228),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1277),
.A2(n_1213),
.B1(n_1188),
.B2(n_1175),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1244),
.A2(n_1247),
.B(n_1251),
.C(n_1234),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1228),
.Y(n_1424)
);

AO31x2_ASAP7_75t_L g1425 ( 
.A1(n_1280),
.A2(n_1170),
.A3(n_1299),
.B(n_1300),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1179),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1156),
.Y(n_1427)
);

AOI22x1_ASAP7_75t_SL g1428 ( 
.A1(n_1216),
.A2(n_1299),
.B1(n_1300),
.B2(n_1170),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1170),
.A2(n_1300),
.B(n_1179),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1154),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1151),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1146),
.B(n_814),
.Y(n_1433)
);

OAI21xp33_ASAP7_75t_L g1434 ( 
.A1(n_1218),
.A2(n_814),
.B(n_788),
.Y(n_1434)
);

O2A1O1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1218),
.A2(n_814),
.B(n_788),
.C(n_652),
.Y(n_1435)
);

AO21x1_ASAP7_75t_L g1436 ( 
.A1(n_1152),
.A2(n_814),
.B(n_788),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1437)
);

AO32x2_ASAP7_75t_L g1438 ( 
.A1(n_1152),
.A2(n_1281),
.A3(n_1243),
.B1(n_1145),
.B2(n_1259),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1440)
);

AO31x2_ASAP7_75t_L g1441 ( 
.A1(n_1254),
.A2(n_1054),
.A3(n_1294),
.B(n_966),
.Y(n_1441)
);

NAND2x1p5_ASAP7_75t_L g1442 ( 
.A(n_1199),
.B(n_1003),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1154),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1150),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1146),
.B(n_1024),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1218),
.A2(n_814),
.B(n_788),
.C(n_1065),
.Y(n_1447)
);

BUFx12f_ASAP7_75t_L g1448 ( 
.A(n_1235),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1150),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1154),
.Y(n_1450)
);

OAI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1183),
.A2(n_814),
.B1(n_788),
.B2(n_660),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1163),
.A2(n_1294),
.B(n_1178),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1453)
);

AO31x2_ASAP7_75t_L g1454 ( 
.A1(n_1254),
.A2(n_1054),
.A3(n_1294),
.B(n_966),
.Y(n_1454)
);

AO22x2_ASAP7_75t_L g1455 ( 
.A1(n_1145),
.A2(n_1065),
.B1(n_1152),
.B2(n_1191),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1154),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1146),
.B(n_814),
.Y(n_1457)
);

AOI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1218),
.A2(n_814),
.B1(n_788),
.B2(n_652),
.C(n_834),
.Y(n_1458)
);

NAND2x1_ASAP7_75t_L g1459 ( 
.A(n_1170),
.B(n_1148),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1146),
.B(n_814),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1461)
);

CKINVDCx6p67_ASAP7_75t_R g1462 ( 
.A(n_1151),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1463)
);

NAND4xp25_ASAP7_75t_L g1464 ( 
.A(n_1147),
.B(n_660),
.C(n_834),
.D(n_885),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1146),
.B(n_942),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1189),
.A2(n_814),
.B(n_802),
.Y(n_1467)
);

NOR2xp67_ASAP7_75t_SL g1468 ( 
.A(n_1206),
.B(n_1011),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1218),
.A2(n_814),
.B(n_788),
.C(n_652),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1160),
.Y(n_1470)
);

AO31x2_ASAP7_75t_L g1471 ( 
.A1(n_1254),
.A2(n_1054),
.A3(n_1294),
.B(n_966),
.Y(n_1471)
);

AO31x2_ASAP7_75t_L g1472 ( 
.A1(n_1254),
.A2(n_1054),
.A3(n_1294),
.B(n_966),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1151),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1183),
.A2(n_814),
.B1(n_788),
.B2(n_660),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1254),
.A2(n_1054),
.A3(n_1294),
.B(n_966),
.Y(n_1475)
);

BUFx2_ASAP7_75t_R g1476 ( 
.A(n_1207),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1146),
.B(n_814),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1167),
.A2(n_1149),
.B(n_1294),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1154),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1227),
.B(n_1024),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1144),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1458),
.A2(n_1464),
.B1(n_1451),
.B2(n_1474),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1330),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1330),
.Y(n_1486)
);

BUFx12f_ASAP7_75t_L g1487 ( 
.A(n_1392),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1362),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1320),
.A2(n_1433),
.B1(n_1447),
.B2(n_1434),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1343),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1446),
.B(n_1457),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1316),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1436),
.A2(n_1455),
.B1(n_1378),
.B2(n_1401),
.Y(n_1493)
);

CKINVDCx11_ASAP7_75t_R g1494 ( 
.A(n_1356),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1455),
.A2(n_1411),
.B1(n_1460),
.B2(n_1477),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1319),
.B(n_1435),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1428),
.A2(n_1372),
.B1(n_1381),
.B2(n_1322),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1343),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1431),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1332),
.Y(n_1500)
);

INVx6_ASAP7_75t_L g1501 ( 
.A(n_1448),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1467),
.A2(n_1352),
.B1(n_1339),
.B2(n_1404),
.Y(n_1502)
);

CKINVDCx11_ASAP7_75t_R g1503 ( 
.A(n_1462),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1338),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1363),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1337),
.A2(n_1369),
.B1(n_1333),
.B2(n_1396),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1431),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1336),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1473),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1345),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1470),
.B(n_1466),
.Y(n_1511)
);

INVx8_ASAP7_75t_L g1512 ( 
.A(n_1317),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1310),
.A2(n_1393),
.B1(n_1421),
.B2(n_1399),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1310),
.A2(n_1482),
.B1(n_1368),
.B2(n_1376),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1413),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_L g1516 ( 
.A(n_1427),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1432),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1313),
.Y(n_1518)
);

BUFx8_ASAP7_75t_L g1519 ( 
.A(n_1403),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1482),
.B(n_1365),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1368),
.A2(n_1324),
.B1(n_1384),
.B2(n_1312),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1350),
.Y(n_1522)
);

INVx6_ASAP7_75t_L g1523 ( 
.A(n_1321),
.Y(n_1523)
);

BUFx12f_ASAP7_75t_L g1524 ( 
.A(n_1358),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1313),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1469),
.A2(n_1366),
.B1(n_1367),
.B2(n_1456),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1456),
.A2(n_1481),
.B1(n_1444),
.B2(n_1450),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1410),
.A2(n_1311),
.B1(n_1314),
.B2(n_1379),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1379),
.A2(n_1402),
.B1(n_1373),
.B2(n_1364),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1364),
.A2(n_1373),
.B1(n_1346),
.B2(n_1391),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1424),
.Y(n_1531)
);

INVx6_ASAP7_75t_L g1532 ( 
.A(n_1395),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1481),
.A2(n_1326),
.B1(n_1429),
.B2(n_1406),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1419),
.A2(n_1351),
.B1(n_1340),
.B2(n_1375),
.Y(n_1534)
);

BUFx2_ASAP7_75t_SL g1535 ( 
.A(n_1418),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_1353),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1406),
.A2(n_1335),
.B1(n_1468),
.B2(n_1422),
.Y(n_1537)
);

INVx4_ASAP7_75t_L g1538 ( 
.A(n_1442),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1414),
.Y(n_1539)
);

CKINVDCx11_ASAP7_75t_R g1540 ( 
.A(n_1476),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1414),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1371),
.A2(n_1397),
.B1(n_1394),
.B2(n_1374),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1414),
.Y(n_1543)
);

CKINVDCx11_ASAP7_75t_R g1544 ( 
.A(n_1395),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_1395),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1382),
.B(n_1341),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1370),
.A2(n_1377),
.B1(n_1380),
.B2(n_1415),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1361),
.A2(n_1360),
.B(n_1387),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1423),
.A2(n_1342),
.B1(n_1405),
.B2(n_1438),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1323),
.A2(n_1385),
.B1(n_1426),
.B2(n_1459),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1418),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1445),
.Y(n_1552)
);

CKINVDCx11_ASAP7_75t_R g1553 ( 
.A(n_1445),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1438),
.A2(n_1420),
.B1(n_1400),
.B2(n_1449),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1438),
.A2(n_1420),
.B1(n_1400),
.B2(n_1449),
.Y(n_1555)
);

CKINVDCx11_ASAP7_75t_R g1556 ( 
.A(n_1445),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1416),
.Y(n_1557)
);

INVx4_ASAP7_75t_L g1558 ( 
.A(n_1478),
.Y(n_1558)
);

BUFx12f_ASAP7_75t_L g1559 ( 
.A(n_1412),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1478),
.A2(n_1409),
.B1(n_1407),
.B2(n_1344),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1318),
.A2(n_1483),
.B1(n_1480),
.B2(n_1443),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1425),
.B(n_1386),
.Y(n_1562)
);

CKINVDCx11_ASAP7_75t_R g1563 ( 
.A(n_1331),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1398),
.Y(n_1564)
);

BUFx10_ASAP7_75t_L g1565 ( 
.A(n_1383),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1425),
.Y(n_1566)
);

INVx6_ASAP7_75t_L g1567 ( 
.A(n_1355),
.Y(n_1567)
);

INVx6_ASAP7_75t_L g1568 ( 
.A(n_1417),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1441),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1441),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1359),
.A2(n_1420),
.B1(n_1465),
.B2(n_1463),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1347),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1349),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1329),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1441),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1454),
.Y(n_1576)
);

INVx5_ASAP7_75t_L g1577 ( 
.A(n_1390),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1430),
.A2(n_1479),
.B1(n_1461),
.B2(n_1453),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1437),
.A2(n_1439),
.B1(n_1440),
.B2(n_1400),
.Y(n_1579)
);

BUFx12f_ASAP7_75t_L g1580 ( 
.A(n_1357),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1386),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1315),
.A2(n_1334),
.B1(n_1325),
.B2(n_1328),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1452),
.A2(n_1388),
.B1(n_1309),
.B2(n_1348),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1327),
.B(n_1475),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1386),
.B(n_1408),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1454),
.B(n_1471),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1454),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1408),
.A2(n_1389),
.B1(n_1471),
.B2(n_1472),
.Y(n_1588)
);

INVx6_ASAP7_75t_L g1589 ( 
.A(n_1354),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1408),
.A2(n_1472),
.B1(n_1475),
.B2(n_1354),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1475),
.A2(n_814),
.B1(n_1458),
.B2(n_788),
.Y(n_1591)
);

CKINVDCx11_ASAP7_75t_R g1592 ( 
.A(n_1354),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_SL g1593 ( 
.A1(n_1433),
.A2(n_1183),
.B1(n_814),
.B2(n_1052),
.Y(n_1593)
);

CKINVDCx14_ASAP7_75t_R g1594 ( 
.A(n_1462),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1433),
.A2(n_1183),
.B1(n_814),
.B2(n_1052),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1451),
.A2(n_1183),
.B1(n_1474),
.B2(n_1464),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1451),
.A2(n_1474),
.B1(n_1458),
.B2(n_1320),
.Y(n_1597)
);

INVx6_ASAP7_75t_L g1598 ( 
.A(n_1363),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1436),
.B(n_1447),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1330),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1602)
);

AOI21xp33_ASAP7_75t_L g1603 ( 
.A1(n_1435),
.A2(n_1469),
.B(n_814),
.Y(n_1603)
);

OAI22x1_ASAP7_75t_L g1604 ( 
.A1(n_1433),
.A2(n_1378),
.B1(n_814),
.B2(n_1322),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_SL g1605 ( 
.A1(n_1433),
.A2(n_1183),
.B1(n_814),
.B2(n_1052),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1330),
.Y(n_1606)
);

INVx6_ASAP7_75t_SL g1607 ( 
.A(n_1482),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1458),
.A2(n_814),
.B(n_1467),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1609)
);

INVx8_ASAP7_75t_L g1610 ( 
.A(n_1363),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1433),
.A2(n_1183),
.B1(n_814),
.B2(n_1052),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1451),
.A2(n_1474),
.B1(n_1458),
.B2(n_1320),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1451),
.A2(n_1474),
.B1(n_1458),
.B2(n_1320),
.Y(n_1615)
);

BUFx8_ASAP7_75t_L g1616 ( 
.A(n_1356),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1451),
.A2(n_1474),
.B1(n_1458),
.B2(n_1320),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1436),
.B(n_1447),
.Y(n_1618)
);

INVx5_ASAP7_75t_L g1619 ( 
.A(n_1363),
.Y(n_1619)
);

INVx6_ASAP7_75t_L g1620 ( 
.A(n_1363),
.Y(n_1620)
);

OAI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1451),
.A2(n_1183),
.B1(n_1474),
.B2(n_1464),
.Y(n_1621)
);

INVx5_ASAP7_75t_L g1622 ( 
.A(n_1363),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1448),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1316),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1626)
);

BUFx8_ASAP7_75t_L g1627 ( 
.A(n_1356),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1436),
.B(n_1447),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1448),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1436),
.B(n_1447),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1631)
);

BUFx8_ASAP7_75t_SL g1632 ( 
.A(n_1356),
.Y(n_1632)
);

NAND2x1p5_ASAP7_75t_L g1633 ( 
.A(n_1468),
.B(n_1003),
.Y(n_1633)
);

BUFx8_ASAP7_75t_L g1634 ( 
.A(n_1356),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1363),
.Y(n_1635)
);

CKINVDCx11_ASAP7_75t_R g1636 ( 
.A(n_1356),
.Y(n_1636)
);

INVx6_ASAP7_75t_L g1637 ( 
.A(n_1363),
.Y(n_1637)
);

OAI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1451),
.A2(n_1183),
.B1(n_1474),
.B2(n_1464),
.Y(n_1638)
);

INVx6_ASAP7_75t_L g1639 ( 
.A(n_1363),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1330),
.Y(n_1641)
);

INVx6_ASAP7_75t_L g1642 ( 
.A(n_1448),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1436),
.B(n_1447),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1644)
);

BUFx4f_ASAP7_75t_SL g1645 ( 
.A(n_1363),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1316),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1448),
.Y(n_1647)
);

BUFx2_ASAP7_75t_SL g1648 ( 
.A(n_1403),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1458),
.A2(n_814),
.B1(n_788),
.B2(n_1464),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1451),
.A2(n_1474),
.B1(n_1458),
.B2(n_1320),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1363),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1541),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1560),
.A2(n_1583),
.B(n_1561),
.Y(n_1653)
);

BUFx4f_ASAP7_75t_SL g1654 ( 
.A(n_1487),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1543),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1485),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1486),
.Y(n_1657)
);

OAI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1608),
.A2(n_1597),
.B1(n_1615),
.B2(n_1614),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1567),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1490),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1584),
.A2(n_1581),
.B(n_1590),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1498),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1539),
.Y(n_1663)
);

OR2x6_ASAP7_75t_L g1664 ( 
.A(n_1566),
.B(n_1546),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1633),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1488),
.B(n_1489),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1545),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1569),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1511),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1570),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1499),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1489),
.B(n_1600),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1508),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1575),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1507),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1562),
.B(n_1585),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1602),
.B(n_1609),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1601),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1582),
.A2(n_1564),
.B(n_1546),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1597),
.A2(n_1615),
.B(n_1614),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1606),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1593),
.A2(n_1611),
.B1(n_1595),
.B2(n_1605),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1574),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1586),
.Y(n_1684)
);

BUFx8_ASAP7_75t_SL g1685 ( 
.A(n_1632),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1617),
.A2(n_1650),
.B(n_1578),
.Y(n_1686)
);

INVxp33_ASAP7_75t_L g1687 ( 
.A(n_1491),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1515),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1608),
.B(n_1502),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1586),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1612),
.B(n_1613),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1641),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1572),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1599),
.B(n_1618),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1566),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1512),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1512),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1628),
.B(n_1630),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1576),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1573),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1496),
.B(n_1628),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1554),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1589),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1540),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1568),
.Y(n_1705)
);

AOI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1584),
.A2(n_1643),
.B(n_1630),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1625),
.B(n_1626),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1520),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1529),
.A2(n_1643),
.B(n_1549),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1496),
.B(n_1555),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1559),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1493),
.B(n_1484),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1587),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1558),
.B(n_1577),
.Y(n_1714)
);

OA21x2_ASAP7_75t_L g1715 ( 
.A1(n_1530),
.A2(n_1528),
.B(n_1603),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1527),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1631),
.B(n_1640),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1527),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1617),
.A2(n_1650),
.B(n_1644),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1568),
.Y(n_1720)
);

INVx4_ASAP7_75t_L g1721 ( 
.A(n_1633),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1592),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1596),
.A2(n_1621),
.B1(n_1638),
.B2(n_1649),
.Y(n_1723)
);

AO21x1_ASAP7_75t_SL g1724 ( 
.A1(n_1513),
.A2(n_1506),
.B(n_1603),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1495),
.B(n_1588),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1492),
.B(n_1500),
.Y(n_1726)
);

OAI21x1_ASAP7_75t_L g1727 ( 
.A1(n_1549),
.A2(n_1526),
.B(n_1533),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1504),
.Y(n_1728)
);

CKINVDCx11_ASAP7_75t_R g1729 ( 
.A(n_1494),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1533),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1557),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1577),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1512),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1579),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1591),
.A2(n_1548),
.B(n_1526),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1577),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1624),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1646),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1577),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1522),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1580),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1604),
.B(n_1537),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1563),
.A2(n_1497),
.B1(n_1521),
.B2(n_1542),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1551),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1542),
.B(n_1548),
.Y(n_1745)
);

BUFx2_ASAP7_75t_SL g1746 ( 
.A(n_1619),
.Y(n_1746)
);

OA21x2_ASAP7_75t_L g1747 ( 
.A1(n_1547),
.A2(n_1571),
.B(n_1514),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1648),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1565),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1552),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1534),
.A2(n_1536),
.B1(n_1623),
.B2(n_1629),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1550),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1565),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1535),
.Y(n_1754)
);

OAI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1619),
.A2(n_1622),
.B1(n_1607),
.B2(n_1501),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1523),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1523),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1531),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_1503),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1532),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1532),
.B(n_1538),
.Y(n_1761)
);

OAI21x1_ASAP7_75t_L g1762 ( 
.A1(n_1607),
.A2(n_1619),
.B(n_1622),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1532),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1619),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1622),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1509),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1622),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1518),
.B(n_1647),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1598),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1598),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1544),
.B(n_1556),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1553),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1594),
.B(n_1651),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1598),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1620),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1501),
.A2(n_1642),
.B1(n_1516),
.B2(n_1510),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1517),
.B(n_1525),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1620),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1620),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1637),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1642),
.A2(n_1524),
.B1(n_1519),
.B2(n_1639),
.Y(n_1781)
);

A2O1A1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1689),
.A2(n_1610),
.B(n_1635),
.C(n_1505),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1743),
.A2(n_1639),
.B1(n_1637),
.B2(n_1645),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1686),
.A2(n_1610),
.B(n_1651),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1666),
.B(n_1610),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1669),
.B(n_1505),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1735),
.A2(n_1505),
.B(n_1635),
.C(n_1651),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1658),
.A2(n_1719),
.B1(n_1680),
.B2(n_1682),
.C(n_1672),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1676),
.B(n_1635),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_SL g1790 ( 
.A1(n_1711),
.A2(n_1616),
.B(n_1627),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1687),
.B(n_1636),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1720),
.B(n_1519),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1676),
.B(n_1616),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1677),
.A2(n_1627),
.B1(n_1634),
.B2(n_1707),
.C(n_1691),
.Y(n_1794)
);

AND2x2_ASAP7_75t_SL g1795 ( 
.A(n_1745),
.B(n_1634),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1722),
.B(n_1708),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1701),
.B(n_1742),
.Y(n_1797)
);

BUFx12f_ASAP7_75t_L g1798 ( 
.A(n_1729),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1723),
.A2(n_1717),
.B1(n_1745),
.B2(n_1751),
.Y(n_1799)
);

AOI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1742),
.A2(n_1712),
.B(n_1741),
.C(n_1755),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1712),
.A2(n_1752),
.B1(n_1725),
.B2(n_1730),
.C(n_1741),
.Y(n_1801)
);

AO32x2_ASAP7_75t_L g1802 ( 
.A1(n_1660),
.A2(n_1692),
.A3(n_1675),
.B1(n_1711),
.B2(n_1702),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1710),
.B(n_1694),
.Y(n_1803)
);

OA21x2_ASAP7_75t_L g1804 ( 
.A1(n_1727),
.A2(n_1679),
.B(n_1709),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1656),
.B(n_1657),
.Y(n_1805)
);

A2O1A1Ixp33_ASAP7_75t_L g1806 ( 
.A1(n_1727),
.A2(n_1709),
.B(n_1752),
.C(n_1725),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1662),
.B(n_1671),
.Y(n_1807)
);

OAI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1715),
.A2(n_1747),
.B1(n_1781),
.B2(n_1776),
.C(n_1734),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1711),
.A2(n_1748),
.B1(n_1753),
.B2(n_1749),
.Y(n_1809)
);

OA21x2_ASAP7_75t_L g1810 ( 
.A1(n_1653),
.A2(n_1734),
.B(n_1730),
.Y(n_1810)
);

AO32x2_ASAP7_75t_L g1811 ( 
.A1(n_1660),
.A2(n_1675),
.A3(n_1692),
.B1(n_1711),
.B2(n_1702),
.Y(n_1811)
);

NOR2x1_ASAP7_75t_L g1812 ( 
.A(n_1753),
.B(n_1749),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1698),
.B(n_1688),
.Y(n_1813)
);

A2O1A1Ixp33_ASAP7_75t_L g1814 ( 
.A1(n_1724),
.A2(n_1739),
.B(n_1732),
.C(n_1736),
.Y(n_1814)
);

AO21x1_ASAP7_75t_L g1815 ( 
.A1(n_1699),
.A2(n_1693),
.B(n_1764),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1731),
.B(n_1659),
.Y(n_1816)
);

NOR2x1_ASAP7_75t_SL g1817 ( 
.A(n_1664),
.B(n_1746),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1724),
.A2(n_1739),
.B(n_1732),
.C(n_1736),
.Y(n_1818)
);

A2O1A1Ixp33_ASAP7_75t_L g1819 ( 
.A1(n_1732),
.A2(n_1736),
.B(n_1739),
.C(n_1718),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1705),
.B(n_1731),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1673),
.B(n_1726),
.Y(n_1821)
);

OR2x2_ASAP7_75t_SL g1822 ( 
.A(n_1772),
.B(n_1774),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1667),
.B(n_1744),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1678),
.B(n_1681),
.Y(n_1824)
);

A2O1A1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1716),
.A2(n_1718),
.B(n_1693),
.C(n_1695),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1769),
.A2(n_1775),
.B1(n_1779),
.B2(n_1778),
.Y(n_1826)
);

AND2x2_ASAP7_75t_SL g1827 ( 
.A(n_1747),
.B(n_1715),
.Y(n_1827)
);

INVxp33_ASAP7_75t_L g1828 ( 
.A(n_1750),
.Y(n_1828)
);

CKINVDCx6p67_ASAP7_75t_R g1829 ( 
.A(n_1759),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1772),
.A2(n_1704),
.B1(n_1654),
.B2(n_1766),
.Y(n_1830)
);

OR2x6_ASAP7_75t_L g1831 ( 
.A(n_1664),
.B(n_1683),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1652),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1769),
.A2(n_1775),
.B1(n_1779),
.B2(n_1778),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1685),
.Y(n_1834)
);

O2A1O1Ixp33_ASAP7_75t_SL g1835 ( 
.A1(n_1770),
.A2(n_1780),
.B(n_1767),
.C(n_1765),
.Y(n_1835)
);

OAI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1715),
.A2(n_1762),
.B(n_1754),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1655),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1714),
.A2(n_1715),
.B(n_1690),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1762),
.A2(n_1767),
.B(n_1765),
.Y(n_1839)
);

OAI211xp5_ASAP7_75t_L g1840 ( 
.A1(n_1706),
.A2(n_1771),
.B(n_1704),
.C(n_1740),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1766),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1770),
.A2(n_1768),
.B1(n_1758),
.B2(n_1665),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1788),
.A2(n_1758),
.B1(n_1771),
.B2(n_1773),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1827),
.B(n_1661),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1788),
.A2(n_1773),
.B1(n_1721),
.B2(n_1761),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1802),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1832),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1827),
.B(n_1661),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1797),
.B(n_1690),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1810),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1799),
.A2(n_1728),
.B1(n_1737),
.B2(n_1738),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1837),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1802),
.B(n_1684),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1810),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1797),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1802),
.B(n_1684),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1794),
.A2(n_1738),
.B1(n_1728),
.B2(n_1737),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1822),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1801),
.A2(n_1721),
.B1(n_1761),
.B2(n_1764),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1811),
.B(n_1700),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1811),
.B(n_1700),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1803),
.B(n_1706),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1838),
.B(n_1674),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1811),
.B(n_1713),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1811),
.B(n_1713),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1812),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1804),
.B(n_1663),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1823),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1836),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1804),
.B(n_1838),
.Y(n_1870)
);

INVx5_ASAP7_75t_L g1871 ( 
.A(n_1831),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1815),
.Y(n_1872)
);

AND2x4_ASAP7_75t_L g1873 ( 
.A(n_1817),
.B(n_1703),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1794),
.A2(n_1777),
.B1(n_1668),
.B2(n_1670),
.Y(n_1874)
);

NAND3xp33_ASAP7_75t_L g1875 ( 
.A(n_1801),
.B(n_1763),
.C(n_1760),
.Y(n_1875)
);

BUFx2_ASAP7_75t_L g1876 ( 
.A(n_1839),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1824),
.Y(n_1877)
);

BUFx12f_ASAP7_75t_L g1878 ( 
.A(n_1798),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1840),
.B(n_1683),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1831),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1805),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1852),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1852),
.Y(n_1883)
);

OAI33xp33_ASAP7_75t_L g1884 ( 
.A1(n_1879),
.A2(n_1809),
.A3(n_1785),
.B1(n_1833),
.B2(n_1826),
.B3(n_1842),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1843),
.A2(n_1808),
.B1(n_1795),
.B2(n_1783),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1852),
.Y(n_1886)
);

OAI31xp33_ASAP7_75t_SL g1887 ( 
.A1(n_1875),
.A2(n_1840),
.A3(n_1808),
.B(n_1816),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1860),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1843),
.A2(n_1845),
.B1(n_1874),
.B2(n_1875),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1855),
.B(n_1813),
.Y(n_1890)
);

NOR3xp33_ASAP7_75t_L g1891 ( 
.A(n_1879),
.B(n_1869),
.C(n_1784),
.Y(n_1891)
);

INVx5_ASAP7_75t_SL g1892 ( 
.A(n_1873),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_SL g1893 ( 
.A1(n_1872),
.A2(n_1795),
.B1(n_1793),
.B2(n_1784),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1876),
.A2(n_1791),
.B1(n_1786),
.B2(n_1790),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1860),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1878),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1868),
.B(n_1796),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1845),
.A2(n_1806),
.B(n_1800),
.Y(n_1898)
);

INVx4_ASAP7_75t_L g1899 ( 
.A(n_1878),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1862),
.B(n_1825),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1860),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1861),
.Y(n_1902)
);

AO21x2_ASAP7_75t_L g1903 ( 
.A1(n_1870),
.A2(n_1872),
.B(n_1854),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1862),
.B(n_1849),
.Y(n_1904)
);

OAI221xp5_ASAP7_75t_L g1905 ( 
.A1(n_1874),
.A2(n_1787),
.B1(n_1814),
.B2(n_1818),
.C(n_1782),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1849),
.B(n_1881),
.Y(n_1906)
);

BUFx2_ASAP7_75t_L g1907 ( 
.A(n_1858),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1869),
.B(n_1807),
.Y(n_1908)
);

AND2x2_ASAP7_75t_SL g1909 ( 
.A(n_1846),
.B(n_1820),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1861),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1844),
.B(n_1821),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1861),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1871),
.B(n_1819),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1881),
.B(n_1825),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1878),
.B(n_1828),
.Y(n_1915)
);

INVx3_ASAP7_75t_L g1916 ( 
.A(n_1873),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1844),
.B(n_1848),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1867),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1848),
.B(n_1880),
.Y(n_1919)
);

NAND3xp33_ASAP7_75t_L g1920 ( 
.A(n_1851),
.B(n_1787),
.C(n_1818),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1867),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1880),
.B(n_1828),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1859),
.A2(n_1857),
.B1(n_1851),
.B2(n_1846),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1847),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_1907),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1888),
.B(n_1846),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1888),
.B(n_1869),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1888),
.B(n_1876),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1882),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1895),
.B(n_1876),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1903),
.B(n_1863),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1882),
.Y(n_1932)
);

INVxp67_ASAP7_75t_L g1933 ( 
.A(n_1884),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1900),
.B(n_1853),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1901),
.B(n_1853),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1901),
.B(n_1853),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1918),
.Y(n_1937)
);

CKINVDCx16_ASAP7_75t_R g1938 ( 
.A(n_1898),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1902),
.B(n_1856),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1902),
.B(n_1856),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1918),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1903),
.B(n_1863),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1902),
.B(n_1856),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1903),
.Y(n_1944)
);

NOR2xp67_ASAP7_75t_L g1945 ( 
.A(n_1913),
.B(n_1871),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1900),
.B(n_1877),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1889),
.A2(n_1898),
.B1(n_1884),
.B2(n_1885),
.Y(n_1947)
);

CKINVDCx16_ASAP7_75t_R g1948 ( 
.A(n_1889),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1910),
.B(n_1858),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1896),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1910),
.B(n_1858),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1903),
.B(n_1863),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1912),
.B(n_1858),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1912),
.B(n_1850),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1883),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1924),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1918),
.B(n_1850),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1917),
.B(n_1864),
.Y(n_1958)
);

BUFx2_ASAP7_75t_L g1959 ( 
.A(n_1909),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1917),
.B(n_1864),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1883),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1921),
.B(n_1854),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1886),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1909),
.B(n_1864),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1921),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1907),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1909),
.B(n_1865),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1919),
.B(n_1865),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1904),
.B(n_1877),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1934),
.B(n_1946),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1956),
.Y(n_1971)
);

AOI21xp33_ASAP7_75t_SL g1972 ( 
.A1(n_1938),
.A2(n_1891),
.B(n_1887),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1956),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1948),
.B(n_1890),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1959),
.B(n_1919),
.Y(n_1975)
);

INVx1_ASAP7_75t_SL g1976 ( 
.A(n_1950),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1933),
.B(n_1899),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1925),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1929),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1948),
.B(n_1890),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1938),
.B(n_1948),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1934),
.B(n_1904),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1959),
.B(n_1892),
.Y(n_1983)
);

INVxp67_ASAP7_75t_L g1984 ( 
.A(n_1950),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1929),
.Y(n_1985)
);

NOR2x1_ASAP7_75t_L g1986 ( 
.A(n_1950),
.B(n_1896),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1929),
.Y(n_1987)
);

AOI21xp33_ASAP7_75t_SL g1988 ( 
.A1(n_1938),
.A2(n_1887),
.B(n_1830),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1959),
.B(n_1892),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1932),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1950),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1947),
.B(n_1911),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1947),
.B(n_1911),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1964),
.B(n_1892),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1932),
.Y(n_1995)
);

AOI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1933),
.A2(n_1923),
.B1(n_1893),
.B2(n_1920),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1946),
.B(n_1922),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1925),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1932),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1955),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1969),
.B(n_1899),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1969),
.B(n_1914),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1945),
.B(n_1893),
.Y(n_2003)
);

OAI32xp33_ASAP7_75t_L g2004 ( 
.A1(n_1931),
.A2(n_1923),
.A3(n_1920),
.B1(n_1914),
.B2(n_1905),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1964),
.B(n_1892),
.Y(n_2005)
);

INVx1_ASAP7_75t_SL g2006 ( 
.A(n_1966),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1964),
.B(n_1892),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1955),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1966),
.B(n_1922),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1955),
.Y(n_2010)
);

BUFx2_ASAP7_75t_L g2011 ( 
.A(n_1967),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1961),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1954),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1928),
.B(n_1897),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1928),
.B(n_1897),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1931),
.B(n_1908),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_2011),
.B(n_1967),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1971),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_2002),
.B(n_1931),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1971),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_2011),
.B(n_1967),
.Y(n_2021)
);

INVxp67_ASAP7_75t_SL g2022 ( 
.A(n_2003),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1985),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1994),
.B(n_1968),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1994),
.B(n_1968),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2005),
.B(n_1968),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_2005),
.B(n_1958),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_2007),
.B(n_1958),
.Y(n_2028)
);

NAND2x1p5_ASAP7_75t_L g2029 ( 
.A(n_1986),
.B(n_1899),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_2002),
.B(n_1942),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1996),
.B(n_1894),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1985),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1977),
.B(n_1958),
.Y(n_2033)
);

OAI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1972),
.A2(n_1905),
.B(n_1915),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1992),
.B(n_1949),
.Y(n_2035)
);

NOR3xp33_ASAP7_75t_SL g2036 ( 
.A(n_1981),
.B(n_1834),
.C(n_1841),
.Y(n_2036)
);

NOR2x1_ASAP7_75t_L g2037 ( 
.A(n_1981),
.B(n_1899),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2007),
.B(n_1975),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1975),
.B(n_1960),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1978),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1982),
.B(n_1942),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1988),
.B(n_1896),
.Y(n_2042)
);

AO21x2_ASAP7_75t_L g2043 ( 
.A1(n_2003),
.A2(n_1944),
.B(n_1942),
.Y(n_2043)
);

INVxp67_ASAP7_75t_L g2044 ( 
.A(n_1974),
.Y(n_2044)
);

INVx1_ASAP7_75t_SL g2045 ( 
.A(n_1998),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1983),
.B(n_1960),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1979),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1983),
.B(n_1945),
.Y(n_2048)
);

INVx1_ASAP7_75t_SL g2049 ( 
.A(n_2006),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1993),
.B(n_1960),
.Y(n_2050)
);

INVxp67_ASAP7_75t_L g2051 ( 
.A(n_1980),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1984),
.B(n_1949),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_1982),
.B(n_1970),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1989),
.B(n_1949),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1976),
.B(n_1951),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_2045),
.B(n_2014),
.Y(n_2056)
);

OAI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_2034),
.A2(n_2004),
.B(n_2001),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2045),
.B(n_2004),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2049),
.B(n_1991),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_2022),
.A2(n_2009),
.B1(n_1989),
.B2(n_1991),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_2033),
.B(n_1970),
.Y(n_2061)
);

INVxp67_ASAP7_75t_L g2062 ( 
.A(n_2040),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2017),
.Y(n_2063)
);

AOI322xp5_ASAP7_75t_L g2064 ( 
.A1(n_2031),
.A2(n_2049),
.A3(n_2050),
.B1(n_2037),
.B2(n_2042),
.C1(n_2051),
.C2(n_2044),
.Y(n_2064)
);

OAI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_2034),
.A2(n_1991),
.B(n_1952),
.Y(n_2065)
);

AOI21xp33_ASAP7_75t_L g2066 ( 
.A1(n_2037),
.A2(n_2043),
.B(n_2035),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2038),
.B(n_1997),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2023),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2023),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2038),
.B(n_2015),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2017),
.B(n_1951),
.Y(n_2071)
);

OAI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_2050),
.A2(n_1944),
.B(n_1952),
.C(n_1859),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2021),
.A2(n_1913),
.B1(n_1951),
.B2(n_1953),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2021),
.B(n_1973),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2033),
.B(n_1953),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2032),
.Y(n_2076)
);

OAI211xp5_ASAP7_75t_L g2077 ( 
.A1(n_2052),
.A2(n_1952),
.B(n_2016),
.C(n_2013),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2039),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2032),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2024),
.B(n_1953),
.Y(n_2080)
);

NAND2x1_ASAP7_75t_L g2081 ( 
.A(n_2048),
.B(n_2013),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2047),
.Y(n_2082)
);

OAI211xp5_ASAP7_75t_L g2083 ( 
.A1(n_2055),
.A2(n_2018),
.B(n_2020),
.C(n_2036),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2047),
.Y(n_2084)
);

INVx3_ASAP7_75t_L g2085 ( 
.A(n_2029),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2063),
.B(n_2054),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2063),
.Y(n_2087)
);

OAI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_2057),
.A2(n_2029),
.B(n_2048),
.Y(n_2088)
);

INVxp67_ASAP7_75t_L g2089 ( 
.A(n_2058),
.Y(n_2089)
);

AOI221xp5_ASAP7_75t_SL g2090 ( 
.A1(n_2065),
.A2(n_2054),
.B1(n_2024),
.B2(n_2025),
.C(n_2026),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2060),
.A2(n_2043),
.B1(n_2048),
.B2(n_2026),
.Y(n_2091)
);

AOI21xp33_ASAP7_75t_L g2092 ( 
.A1(n_2062),
.A2(n_2043),
.B(n_2029),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_2062),
.A2(n_2056),
.B1(n_2083),
.B2(n_2070),
.Y(n_2093)
);

NAND2x1p5_ASAP7_75t_L g2094 ( 
.A(n_2085),
.B(n_2048),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2068),
.Y(n_2095)
);

BUFx2_ASAP7_75t_SL g2096 ( 
.A(n_2085),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_2059),
.B(n_1878),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2069),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2076),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2064),
.B(n_2025),
.Y(n_2100)
);

AOI211xp5_ASAP7_75t_SL g2101 ( 
.A1(n_2066),
.A2(n_2085),
.B(n_2077),
.C(n_2072),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2079),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2074),
.Y(n_2103)
);

AOI32xp33_ASAP7_75t_L g2104 ( 
.A1(n_2074),
.A2(n_2027),
.A3(n_2028),
.B1(n_2046),
.B2(n_2039),
.Y(n_2104)
);

NOR3xp33_ASAP7_75t_L g2105 ( 
.A(n_2082),
.B(n_2020),
.C(n_2018),
.Y(n_2105)
);

INVx1_ASAP7_75t_SL g2106 ( 
.A(n_2081),
.Y(n_2106)
);

A2O1A1Ixp33_ASAP7_75t_L g2107 ( 
.A1(n_2073),
.A2(n_2053),
.B(n_2019),
.C(n_2030),
.Y(n_2107)
);

OAI221xp5_ASAP7_75t_L g2108 ( 
.A1(n_2067),
.A2(n_2053),
.B1(n_2027),
.B2(n_2028),
.C(n_2046),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2084),
.Y(n_2109)
);

OAI211xp5_ASAP7_75t_L g2110 ( 
.A1(n_2101),
.A2(n_2100),
.B(n_2091),
.C(n_2088),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2087),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_2093),
.B(n_2061),
.Y(n_2112)
);

NOR2x1_ASAP7_75t_L g2113 ( 
.A(n_2096),
.B(n_2078),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2103),
.Y(n_2114)
);

NOR3xp33_ASAP7_75t_L g2115 ( 
.A(n_2097),
.B(n_2089),
.C(n_2092),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2094),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_2089),
.B(n_2078),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2086),
.B(n_2071),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2095),
.Y(n_2119)
);

OAI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_2106),
.A2(n_2061),
.B1(n_2075),
.B2(n_2080),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2098),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_2094),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2099),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2102),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2109),
.Y(n_2125)
);

OAI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_2107),
.A2(n_2030),
.B(n_2019),
.Y(n_2126)
);

NOR3xp33_ASAP7_75t_L g2127 ( 
.A(n_2110),
.B(n_2108),
.C(n_2105),
.Y(n_2127)
);

NOR2xp67_ASAP7_75t_L g2128 ( 
.A(n_2116),
.B(n_2041),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_SL g2129 ( 
.A1(n_2126),
.A2(n_2112),
.B1(n_2122),
.B2(n_2120),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2111),
.Y(n_2130)
);

OAI211xp5_ASAP7_75t_L g2131 ( 
.A1(n_2113),
.A2(n_2115),
.B(n_2117),
.C(n_2116),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2117),
.B(n_2118),
.Y(n_2132)
);

AOI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_2114),
.A2(n_2090),
.B1(n_2105),
.B2(n_1913),
.Y(n_2133)
);

NOR2x1_ASAP7_75t_L g2134 ( 
.A(n_2123),
.B(n_2041),
.Y(n_2134)
);

OAI21xp33_ASAP7_75t_L g2135 ( 
.A1(n_2119),
.A2(n_2104),
.B(n_2016),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_2121),
.B(n_1829),
.Y(n_2136)
);

AOI21xp33_ASAP7_75t_L g2137 ( 
.A1(n_2111),
.A2(n_2012),
.B(n_1990),
.Y(n_2137)
);

NOR4xp25_ASAP7_75t_L g2138 ( 
.A(n_2124),
.B(n_2010),
.C(n_2008),
.D(n_2000),
.Y(n_2138)
);

NOR3xp33_ASAP7_75t_L g2139 ( 
.A(n_2125),
.B(n_1782),
.C(n_1792),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2123),
.B(n_1928),
.Y(n_2140)
);

A2O1A1Ixp33_ASAP7_75t_L g2141 ( 
.A1(n_2110),
.A2(n_1930),
.B(n_1866),
.C(n_1927),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2134),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2130),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2128),
.Y(n_2144)
);

OAI221xp5_ASAP7_75t_L g2145 ( 
.A1(n_2129),
.A2(n_1857),
.B1(n_1995),
.B2(n_1987),
.C(n_1999),
.Y(n_2145)
);

INVx8_ASAP7_75t_L g2146 ( 
.A(n_2132),
.Y(n_2146)
);

AND4x1_ASAP7_75t_L g2147 ( 
.A(n_2127),
.B(n_1814),
.C(n_1927),
.D(n_1930),
.Y(n_2147)
);

OAI211xp5_ASAP7_75t_SL g2148 ( 
.A1(n_2141),
.A2(n_1906),
.B(n_1954),
.C(n_1789),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_2131),
.A2(n_1792),
.B(n_1927),
.Y(n_2149)
);

AOI221xp5_ASAP7_75t_L g2150 ( 
.A1(n_2142),
.A2(n_2135),
.B1(n_2138),
.B2(n_2137),
.C(n_2133),
.Y(n_2150)
);

AOI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_2145),
.A2(n_2144),
.B1(n_2149),
.B2(n_2143),
.C(n_2146),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2147),
.Y(n_2152)
);

OAI21xp5_ASAP7_75t_SL g2153 ( 
.A1(n_2148),
.A2(n_2136),
.B(n_2139),
.Y(n_2153)
);

AOI221xp5_ASAP7_75t_L g2154 ( 
.A1(n_2142),
.A2(n_2140),
.B1(n_1930),
.B2(n_1866),
.C(n_1870),
.Y(n_2154)
);

AOI211x1_ASAP7_75t_SL g2155 ( 
.A1(n_2149),
.A2(n_1965),
.B(n_1941),
.C(n_1937),
.Y(n_2155)
);

NAND3xp33_ASAP7_75t_L g2156 ( 
.A(n_2142),
.B(n_1757),
.C(n_1756),
.Y(n_2156)
);

NAND3xp33_ASAP7_75t_L g2157 ( 
.A(n_2142),
.B(n_1757),
.C(n_1756),
.Y(n_2157)
);

INVxp67_ASAP7_75t_L g2158 ( 
.A(n_2152),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2156),
.Y(n_2159)
);

NAND4xp75_ASAP7_75t_L g2160 ( 
.A(n_2151),
.B(n_1926),
.C(n_1733),
.D(n_1696),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2157),
.Y(n_2161)
);

NOR2x1_ASAP7_75t_L g2162 ( 
.A(n_2153),
.B(n_1954),
.Y(n_2162)
);

AND2x4_ASAP7_75t_SL g2163 ( 
.A(n_2150),
.B(n_2155),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2154),
.B(n_1926),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_2162),
.A2(n_1941),
.B(n_1937),
.Y(n_2165)
);

AOI211xp5_ASAP7_75t_SL g2166 ( 
.A1(n_2158),
.A2(n_1835),
.B(n_1913),
.C(n_1962),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2160),
.A2(n_2163),
.B1(n_2161),
.B2(n_2159),
.Y(n_2167)
);

BUFx2_ASAP7_75t_L g2168 ( 
.A(n_2167),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2168),
.Y(n_2169)
);

XOR2x1_ASAP7_75t_L g2170 ( 
.A(n_2169),
.B(n_2159),
.Y(n_2170)
);

XNOR2x1_ASAP7_75t_L g2171 ( 
.A(n_2169),
.B(n_2164),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_2171),
.A2(n_2165),
.B1(n_2166),
.B2(n_1916),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_L g2173 ( 
.A(n_2170),
.B(n_1957),
.Y(n_2173)
);

AO21x2_ASAP7_75t_L g2174 ( 
.A1(n_2173),
.A2(n_1941),
.B(n_1937),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2172),
.Y(n_2175)
);

AOI322xp5_ASAP7_75t_SL g2176 ( 
.A1(n_2174),
.A2(n_1926),
.A3(n_1939),
.B1(n_1936),
.B2(n_1943),
.C1(n_1935),
.C2(n_1940),
.Y(n_2176)
);

AOI22x1_ASAP7_75t_L g2177 ( 
.A1(n_2176),
.A2(n_2175),
.B1(n_2174),
.B2(n_1696),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2177),
.Y(n_2178)
);

AOI221xp5_ASAP7_75t_L g2179 ( 
.A1(n_2178),
.A2(n_1961),
.B1(n_1963),
.B2(n_1941),
.C(n_1965),
.Y(n_2179)
);

AOI211xp5_ASAP7_75t_L g2180 ( 
.A1(n_2179),
.A2(n_1697),
.B(n_1733),
.C(n_1835),
.Y(n_2180)
);


endmodule