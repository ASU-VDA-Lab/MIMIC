module real_jpeg_25175_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g11 ( 
.A1(n_1),
.A2(n_12),
.B(n_21),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_4),
.Y(n_10)
);

AO21x1_ASAP7_75t_SL g16 ( 
.A1(n_2),
.A2(n_17),
.B(n_19),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_18),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_11),
.B1(n_24),
.B2(n_25),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_9),
.B(n_10),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_8),
.B(n_15),
.Y(n_14)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_13),
.A2(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_20),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);


endmodule