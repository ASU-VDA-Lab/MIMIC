module fake_jpeg_12992_n_261 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_44),
.B(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_3),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_47),
.B(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_3),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_4),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_25),
.B(n_5),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_69),
.Y(n_100)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_54),
.B(n_70),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_68),
.Y(n_109)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_9),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_27),
.B(n_6),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_28),
.B(n_6),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_36),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_31),
.B1(n_23),
.B2(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_93),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_23),
.B1(n_37),
.B2(n_34),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_37),
.B1(n_34),
.B2(n_31),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_30),
.B1(n_39),
.B2(n_28),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_73),
.B1(n_64),
.B2(n_61),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_51),
.B(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_92),
.Y(n_121)
);

AO22x1_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_21),
.B1(n_29),
.B2(n_22),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_42),
.B(n_35),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_35),
.B1(n_21),
.B2(n_29),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_22),
.B1(n_30),
.B2(n_36),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_95),
.A2(n_102),
.B1(n_114),
.B2(n_76),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_106),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_56),
.B(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_107),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_8),
.B(n_9),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_108),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_36),
.B1(n_40),
.B2(n_11),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_114),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_10),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_46),
.A2(n_40),
.B(n_13),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_67),
.A2(n_40),
.B1(n_13),
.B2(n_14),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_102),
.B1(n_100),
.B2(n_87),
.Y(n_137)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_143),
.Y(n_162)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_119),
.Y(n_167)
);

AO21x2_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_124),
.B(n_149),
.Y(n_164)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_60),
.B1(n_71),
.B2(n_53),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_59),
.C(n_40),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_11),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_132),
.B(n_136),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_14),
.B1(n_77),
.B2(n_78),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_148),
.B(n_126),
.Y(n_172)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_144),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_86),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_141),
.B1(n_142),
.B2(n_80),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_145),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_110),
.B1(n_82),
.B2(n_90),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_106),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_82),
.A2(n_85),
.B1(n_90),
.B2(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_83),
.B(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_149),
.Y(n_174)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_106),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_153),
.B(n_154),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_158),
.A2(n_171),
.B1(n_117),
.B2(n_127),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_80),
.B1(n_138),
.B2(n_116),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_181),
.B1(n_175),
.B2(n_174),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_119),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_145),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_137),
.B1(n_151),
.B2(n_139),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_178),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_129),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_121),
.B(n_130),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_180),
.B(n_148),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_132),
.A2(n_128),
.B1(n_149),
.B2(n_152),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_165),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_184),
.Y(n_210)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_188),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_197),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_123),
.C(n_125),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_194),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_132),
.B(n_149),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_162),
.B(n_176),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_164),
.B1(n_173),
.B2(n_159),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_134),
.Y(n_194)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_156),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_176),
.A3(n_164),
.B1(n_182),
.B2(n_179),
.C1(n_157),
.C2(n_155),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_163),
.C(n_156),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_198),
.A2(n_164),
.B1(n_172),
.B2(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_161),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_159),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_168),
.B1(n_158),
.B2(n_163),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_164),
.B1(n_157),
.B2(n_179),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_214),
.B1(n_218),
.B2(n_167),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_196),
.B(n_197),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_216),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_195),
.A3(n_191),
.B1(n_193),
.B2(n_187),
.C1(n_202),
.C2(n_198),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_201),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_155),
.B1(n_167),
.B2(n_182),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_227),
.B1(n_229),
.B2(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_194),
.C(n_190),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_200),
.C(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_185),
.C(n_167),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_228),
.A2(n_212),
.B(n_207),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_164),
.B1(n_203),
.B2(n_216),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_210),
.C(n_209),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_240),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_229),
.B1(n_227),
.B2(n_222),
.Y(n_247)
);

NOR4xp25_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_210),
.C(n_211),
.D(n_207),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_236),
.B(n_239),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_221),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_215),
.B(n_219),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_218),
.B(n_205),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_223),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_244),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_215),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_247),
.B(n_244),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_245),
.A2(n_240),
.B1(n_205),
.B2(n_208),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_250),
.B1(n_164),
.B2(n_252),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_237),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_243),
.B1(n_225),
.B2(n_213),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_248),
.A2(n_228),
.B1(n_241),
.B2(n_217),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_237),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_255),
.A2(n_256),
.B(n_252),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_257),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_250),
.B(n_253),
.C(n_254),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_260),
.B(n_258),
.Y(n_261)
);


endmodule