module fake_netlist_6_3435_n_1655 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1655);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1655;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1605;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_16),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_11),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_60),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_44),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_19),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_77),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_33),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_44),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_122),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_121),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_36),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_94),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_57),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_9),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_20),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_147),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_6),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_18),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_126),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_52),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_48),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_38),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_55),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_79),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_42),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_110),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_21),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_45),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_61),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_71),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_96),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_12),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_114),
.Y(n_196)
);

BUFx2_ASAP7_75t_SL g197 ( 
.A(n_40),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_58),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_64),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_63),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_134),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_8),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_36),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_81),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_19),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_34),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_4),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_106),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_70),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_35),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_85),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_101),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_124),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_32),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_14),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_86),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_59),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_5),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_103),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_38),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_74),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_123),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_30),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_136),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_17),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_128),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_144),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_1),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_50),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_67),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_75),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_1),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_73),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_48),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_76),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_88),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_7),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_3),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_99),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_102),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_84),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_90),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_91),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_25),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_27),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_4),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_3),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_10),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_135),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_120),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_8),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_18),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_127),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_9),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_47),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_56),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_145),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_65),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_0),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_125),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_118),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_30),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_53),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_51),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_83),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_21),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_47),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_92),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_130),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_111),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_23),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_5),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_31),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_97),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_152),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_27),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_119),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_69),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_133),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_15),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_46),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_33),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_95),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_131),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_22),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_26),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_17),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_113),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_149),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_132),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_62),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_107),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_109),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_54),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_72),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_40),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_163),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_186),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_166),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_190),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_191),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_235),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_220),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_153),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_153),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_257),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_153),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_179),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_205),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_153),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_238),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_153),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_211),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_212),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_241),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_192),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_273),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_245),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_175),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_187),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_211),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_187),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_212),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_193),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_196),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_249),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_249),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_157),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_208),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_156),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_228),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_230),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_154),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_252),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_198),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_258),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_200),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_201),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_202),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_261),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_209),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_269),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_213),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_280),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_288),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_215),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_290),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_293),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_294),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_181),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_216),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_217),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_218),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_154),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_181),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_243),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_155),
.Y(n_378)
);

NOR2x1_ASAP7_75t_L g379 ( 
.A(n_321),
.B(n_160),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_356),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_330),
.B(n_212),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_323),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g384 ( 
.A(n_327),
.B(n_160),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_305),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_310),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_305),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_306),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_320),
.B(n_155),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_306),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_308),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_320),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_311),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_329),
.B(n_210),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_311),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_320),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_312),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_316),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_316),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_372),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_313),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_352),
.B(n_161),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_317),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_324),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_333),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_340),
.B(n_210),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_314),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_348),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_325),
.A2(n_304),
.B1(n_164),
.B2(n_167),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_333),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_337),
.A2(n_262),
.B1(n_266),
.B2(n_171),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_355),
.A2(n_278),
.B(n_248),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_339),
.B(n_162),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_331),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_373),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_335),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_359),
.B(n_248),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_339),
.B(n_278),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_315),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_347),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_330),
.B(n_327),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_338),
.A2(n_296),
.B(n_287),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_387),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_387),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

AOI21x1_ASAP7_75t_L g445 ( 
.A1(n_407),
.A2(n_296),
.B(n_287),
.Y(n_445)
);

NOR2x1p5_ASAP7_75t_L g446 ( 
.A(n_389),
.B(n_342),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_387),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_396),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_407),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_396),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_420),
.Y(n_454)
);

OR2x6_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_197),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_411),
.B(n_332),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_378),
.B(n_343),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_396),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_390),
.Y(n_463)
);

INVx6_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_414),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_398),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_398),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_384),
.B(n_344),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_398),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_414),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_400),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_384),
.A2(n_322),
.B1(n_318),
.B2(n_214),
.Y(n_474)
);

AOI21x1_ASAP7_75t_L g475 ( 
.A1(n_441),
.A2(n_177),
.B(n_159),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_400),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_402),
.B(n_341),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_384),
.B(n_354),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_378),
.B(n_358),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_400),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_418),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_427),
.B(n_307),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_384),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_401),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_L g487 ( 
.A(n_378),
.B(n_360),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_402),
.A2(n_417),
.B1(n_432),
.B2(n_433),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_401),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_403),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_417),
.Y(n_493)
);

INVxp33_ASAP7_75t_L g494 ( 
.A(n_422),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_435),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_417),
.B(n_363),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_382),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_390),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_420),
.B(n_319),
.Y(n_499)
);

AOI21x1_ASAP7_75t_L g500 ( 
.A1(n_441),
.A2(n_184),
.B(n_183),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_403),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_390),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_392),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_404),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_404),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_435),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_412),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_432),
.A2(n_243),
.B1(n_374),
.B2(n_229),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_382),
.B(n_366),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_438),
.B(n_371),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_390),
.Y(n_516)
);

AO21x2_ASAP7_75t_L g517 ( 
.A1(n_425),
.A2(n_194),
.B(n_189),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_381),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_412),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_438),
.B(n_342),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_412),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_431),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_390),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_433),
.B(n_341),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_391),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_380),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_437),
.B(n_345),
.Y(n_527)
);

INVx8_ASAP7_75t_L g528 ( 
.A(n_392),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_392),
.B(n_433),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_392),
.B(n_169),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_437),
.B(n_345),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_422),
.B(n_297),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_380),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_397),
.B(n_182),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_383),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_439),
.B(n_346),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_432),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_439),
.B(n_346),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_377),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_397),
.B(n_271),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_391),
.Y(n_541)
);

INVx8_ASAP7_75t_L g542 ( 
.A(n_391),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_391),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_377),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_410),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_377),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_410),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_397),
.B(n_227),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_432),
.A2(n_229),
.B1(n_369),
.B2(n_368),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_381),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_391),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_383),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_386),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_377),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_377),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_397),
.B(n_232),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_432),
.B(n_297),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_395),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_395),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_391),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_385),
.B(n_297),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_385),
.B(n_162),
.Y(n_562)
);

BUFx6f_ASAP7_75t_SL g563 ( 
.A(n_440),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_391),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_440),
.B(n_388),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_397),
.B(n_234),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_415),
.B(n_338),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_395),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_395),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_441),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_388),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_409),
.B(n_165),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_399),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_399),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_409),
.B(n_165),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_430),
.Y(n_576)
);

OAI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_425),
.A2(n_376),
.B(n_375),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_415),
.B(n_370),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_391),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_395),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_441),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_425),
.A2(n_272),
.B(n_285),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_393),
.Y(n_583)
);

NOR3xp33_ASAP7_75t_L g584 ( 
.A(n_430),
.B(n_239),
.C(n_203),
.Y(n_584)
);

NOR2x1p5_ASAP7_75t_L g585 ( 
.A(n_419),
.B(n_158),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_441),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_441),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_419),
.B(n_370),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_529),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_493),
.B(n_393),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_442),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_496),
.B(n_168),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_442),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_442),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_529),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_457),
.B(n_168),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_484),
.B(n_393),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_528),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_443),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_493),
.B(n_393),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_529),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_443),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_529),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_488),
.B(n_393),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_511),
.B(n_375),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_484),
.B(n_393),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_524),
.B(n_350),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_505),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_451),
.B(n_458),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_L g610 ( 
.A(n_469),
.B(n_222),
.C(n_199),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_531),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_531),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_479),
.B(n_393),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_538),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_538),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_490),
.B(n_393),
.Y(n_616)
);

BUFx8_ASAP7_75t_L g617 ( 
.A(n_563),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_451),
.B(n_394),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_458),
.B(n_394),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_497),
.A2(n_231),
.B1(n_224),
.B2(n_226),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_478),
.B(n_303),
.C(n_236),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_460),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_490),
.B(n_394),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_483),
.B(n_172),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_465),
.B(n_394),
.Y(n_626)
);

BUFx6f_ASAP7_75t_SL g627 ( 
.A(n_518),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_477),
.B(n_351),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_460),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_464),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_577),
.A2(n_379),
.B(n_300),
.C(n_292),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_465),
.B(n_394),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_528),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_528),
.B(n_240),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_471),
.B(n_394),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_537),
.B(n_394),
.Y(n_636)
);

BUFx8_ASAP7_75t_L g637 ( 
.A(n_563),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_514),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_585),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_471),
.B(n_394),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_462),
.B(n_406),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_537),
.B(n_406),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_462),
.B(n_570),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_526),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_483),
.B(n_172),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_474),
.B(n_487),
.C(n_513),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_526),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_552),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_462),
.B(n_406),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_524),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_577),
.B(n_406),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_581),
.B(n_406),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_581),
.B(n_406),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_528),
.B(n_256),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_586),
.B(n_406),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_586),
.B(n_406),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_552),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_587),
.A2(n_405),
.B(n_434),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_466),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_587),
.B(n_423),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_534),
.B(n_423),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_455),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_464),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_553),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_456),
.B(n_173),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_455),
.B(n_173),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_468),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_448),
.B(n_174),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_455),
.B(n_174),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_L g670 ( 
.A1(n_494),
.A2(n_158),
.B1(n_274),
.B2(n_275),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_448),
.B(n_351),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_522),
.B(n_353),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_540),
.B(n_229),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_547),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_468),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_455),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_455),
.B(n_178),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_464),
.A2(n_221),
.B1(n_178),
.B2(n_263),
.Y(n_678)
);

BUFx5_ASAP7_75t_L g679 ( 
.A(n_502),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_448),
.B(n_229),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_SL g681 ( 
.A1(n_532),
.A2(n_170),
.B1(n_275),
.B2(n_284),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_464),
.A2(n_563),
.B1(n_530),
.B2(n_515),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_588),
.B(n_361),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_L g684 ( 
.A(n_520),
.B(n_221),
.C(n_263),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_571),
.B(n_423),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_571),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_573),
.B(n_423),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_448),
.B(n_229),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_573),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_574),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_574),
.B(n_423),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_567),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_565),
.B(n_424),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_468),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_533),
.B(n_424),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_SL g696 ( 
.A(n_563),
.B(n_170),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_557),
.B(n_264),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_470),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_470),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_548),
.B(n_260),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_556),
.B(n_291),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_533),
.B(n_424),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_535),
.B(n_424),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_535),
.B(n_424),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_482),
.B(n_264),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_566),
.B(n_416),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_567),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_470),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_472),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_588),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_453),
.B(n_416),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_583),
.B(n_560),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_583),
.B(n_265),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_527),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_517),
.A2(n_176),
.B1(n_284),
.B2(n_180),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_453),
.B(n_416),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_463),
.B(n_416),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_463),
.B(n_416),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_536),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_578),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_517),
.A2(n_582),
.B1(n_549),
.B2(n_473),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_463),
.B(n_416),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_463),
.B(n_421),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_467),
.B(n_421),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_576),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_562),
.B(n_265),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_560),
.Y(n_727)
);

BUFx6f_ASAP7_75t_SL g728 ( 
.A(n_518),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_467),
.B(n_516),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_467),
.B(n_421),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_572),
.B(n_267),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_516),
.B(n_421),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_446),
.B(n_361),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_583),
.B(n_560),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_446),
.B(n_267),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_560),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_516),
.B(n_421),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_580),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_516),
.B(n_421),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_525),
.B(n_421),
.Y(n_740)
);

BUFx6f_ASAP7_75t_SL g741 ( 
.A(n_518),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_525),
.B(n_436),
.Y(n_742)
);

BUFx4f_ASAP7_75t_L g743 ( 
.A(n_605),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_646),
.A2(n_584),
.B1(n_582),
.B2(n_517),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_720),
.B(n_495),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_720),
.B(n_509),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_692),
.B(n_473),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_692),
.B(n_476),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_714),
.B(n_476),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_719),
.B(n_481),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_589),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_725),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_604),
.A2(n_561),
.B1(n_575),
.B2(n_475),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_SL g754 ( 
.A1(n_674),
.A2(n_454),
.B1(n_413),
.B2(n_428),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_595),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_633),
.B(n_502),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_609),
.B(n_481),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_650),
.B(n_545),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_596),
.B(n_413),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_672),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_671),
.B(n_550),
.Y(n_761)
);

AND3x4_ASAP7_75t_L g762 ( 
.A(n_684),
.B(n_454),
.C(n_499),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_627),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_643),
.B(n_485),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_652),
.A2(n_542),
.B(n_582),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_644),
.B(n_485),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_652),
.A2(n_655),
.B(n_653),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_601),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_603),
.A2(n_525),
.B1(n_541),
.B2(n_564),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_647),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_610),
.A2(n_622),
.B1(n_715),
.B2(n_624),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_738),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_648),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_738),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_662),
.Y(n_775)
);

O2A1O1Ixp5_ASAP7_75t_L g776 ( 
.A1(n_631),
.A2(n_445),
.B(n_500),
.C(n_475),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_L g777 ( 
.A(n_633),
.B(n_502),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_592),
.A2(n_525),
.B1(n_564),
.B2(n_541),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_657),
.B(n_486),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_662),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_596),
.B(n_428),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_664),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_607),
.B(n_362),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_591),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_593),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_L g786 ( 
.A(n_665),
.B(n_499),
.C(n_188),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_733),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_676),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_594),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_599),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_592),
.A2(n_543),
.B1(n_541),
.B2(n_551),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_663),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_663),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_665),
.B(n_550),
.Y(n_794)
);

OR2x6_ASAP7_75t_L g795 ( 
.A(n_676),
.B(n_550),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_610),
.A2(n_543),
.B1(n_541),
.B2(n_551),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_633),
.B(n_560),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_607),
.Y(n_798)
);

INVx5_ASAP7_75t_L g799 ( 
.A(n_633),
.Y(n_799)
);

AND2x6_ASAP7_75t_SL g800 ( 
.A(n_726),
.B(n_362),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_683),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_L g802 ( 
.A(n_663),
.B(n_560),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_622),
.A2(n_543),
.B1(n_564),
.B2(n_551),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_625),
.B(n_550),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_686),
.B(n_486),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_602),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_616),
.A2(n_551),
.B1(n_543),
.B2(n_564),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_689),
.B(n_492),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_690),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_693),
.B(n_492),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_628),
.Y(n_811)
);

AND3x1_ASAP7_75t_SL g812 ( 
.A(n_710),
.B(n_367),
.C(n_364),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_611),
.B(n_507),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_612),
.B(n_507),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_645),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_639),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_715),
.A2(n_510),
.B1(n_519),
.B2(n_512),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_614),
.B(n_510),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_615),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_613),
.B(n_512),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_668),
.B(n_498),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_613),
.B(n_519),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_608),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_682),
.B(n_268),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_726),
.B(n_268),
.Y(n_825)
);

AND3x2_ASAP7_75t_SL g826 ( 
.A(n_681),
.B(n_670),
.C(n_669),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_617),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_663),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_707),
.B(n_521),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_590),
.B(n_521),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_600),
.B(n_444),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_616),
.A2(n_624),
.B1(n_731),
.B2(n_669),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_L g833 ( 
.A1(n_638),
.A2(n_299),
.B1(n_302),
.B2(n_270),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_617),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_660),
.B(n_444),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_685),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_687),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_656),
.A2(n_542),
.B(n_498),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_691),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_666),
.A2(n_480),
.B1(n_447),
.B2(n_449),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_731),
.A2(n_523),
.B1(n_498),
.B2(n_579),
.Y(n_841)
);

BUFx12f_ASAP7_75t_L g842 ( 
.A(n_637),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_597),
.B(n_447),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_597),
.B(n_449),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_SL g845 ( 
.A(n_684),
.B(n_697),
.C(n_677),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_666),
.B(n_365),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_637),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_721),
.A2(n_500),
.B1(n_523),
.B2(n_276),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_677),
.B(n_276),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_627),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_700),
.A2(n_523),
.B1(n_579),
.B2(n_498),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_SL g852 ( 
.A1(n_728),
.A2(n_741),
.B1(n_621),
.B2(n_274),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_705),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_700),
.A2(n_579),
.B1(n_480),
.B2(n_450),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_623),
.Y(n_855)
);

BUFx8_ASAP7_75t_L g856 ( 
.A(n_728),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_629),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_678),
.B(n_579),
.Y(n_858)
);

AND2x2_ASAP7_75t_SL g859 ( 
.A(n_735),
.B(n_365),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_721),
.A2(n_277),
.B1(n_282),
.B2(n_283),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_695),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_701),
.A2(n_459),
.B1(n_450),
.B2(n_452),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_696),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_702),
.Y(n_864)
);

INVxp67_ASAP7_75t_SL g865 ( 
.A(n_727),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_630),
.B(n_367),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_598),
.B(n_368),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_606),
.B(n_661),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_703),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_704),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_651),
.A2(n_542),
.B(n_452),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_598),
.B(n_369),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_713),
.B(n_426),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_620),
.B(n_277),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_620),
.B(n_282),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_701),
.A2(n_459),
.B1(n_503),
.B2(n_489),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_606),
.B(n_489),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_727),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_618),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_658),
.B(n_491),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_619),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_741),
.A2(n_204),
.B1(n_185),
.B2(n_195),
.Y(n_882)
);

AND2x6_ASAP7_75t_SL g883 ( 
.A(n_626),
.B(n_426),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_713),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_680),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_680),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_SL g887 ( 
.A1(n_688),
.A2(n_206),
.B1(n_207),
.B2(n_219),
.Y(n_887)
);

BUFx4f_ASAP7_75t_L g888 ( 
.A(n_727),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_679),
.B(n_491),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_736),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_651),
.A2(n_542),
.B(n_491),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_688),
.Y(n_892)
);

AO22x1_ASAP7_75t_L g893 ( 
.A1(n_729),
.A2(n_223),
.B1(n_225),
.B2(n_233),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_641),
.B(n_283),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_649),
.B(n_429),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_679),
.B(n_501),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_736),
.B(n_286),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_632),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_736),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_635),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_673),
.A2(n_503),
.B1(n_504),
.B2(n_506),
.Y(n_901)
);

OAI22xp33_ASAP7_75t_L g902 ( 
.A1(n_640),
.A2(n_706),
.B1(n_742),
.B2(n_673),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_659),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_712),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_667),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_675),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_679),
.B(n_636),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_694),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_698),
.Y(n_909)
);

AND2x6_ASAP7_75t_SL g910 ( 
.A(n_711),
.B(n_429),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_836),
.B(n_679),
.Y(n_911)
);

OAI22x1_ASAP7_75t_L g912 ( 
.A1(n_762),
.A2(n_289),
.B1(n_242),
.B2(n_250),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_888),
.A2(n_542),
.B(n_654),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_815),
.A2(n_634),
.B(n_636),
.C(n_642),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_758),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_804),
.B(n_679),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_784),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_819),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_770),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_832),
.A2(n_740),
.B(n_739),
.C(n_737),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_845),
.A2(n_699),
.B1(n_708),
.B2(n_709),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_797),
.A2(n_734),
.B(n_712),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_745),
.B(n_734),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_890),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_846),
.B(n_811),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_758),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_802),
.A2(n_896),
.B(n_889),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_889),
.A2(n_716),
.B(n_730),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_760),
.B(n_237),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_794),
.A2(n_732),
.B(n_724),
.C(n_723),
.Y(n_930)
);

CKINVDCx8_ASAP7_75t_R g931 ( 
.A(n_752),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_825),
.A2(n_722),
.B(n_718),
.C(n_717),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_746),
.B(n_251),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_842),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_771),
.A2(n_302),
.B(n_298),
.C(n_299),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_775),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_773),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_792),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_892),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_R g940 ( 
.A(n_763),
.B(n_298),
.Y(n_940)
);

CKINVDCx11_ASAP7_75t_R g941 ( 
.A(n_827),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_780),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_786),
.A2(n_301),
.B(n_508),
.C(n_501),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_759),
.B(n_259),
.Y(n_944)
);

NOR2x1_ASAP7_75t_L g945 ( 
.A(n_828),
.B(n_504),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_884),
.A2(n_301),
.B(n_503),
.C(n_504),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_787),
.B(n_506),
.Y(n_947)
);

OAI22x1_ASAP7_75t_L g948 ( 
.A1(n_781),
.A2(n_886),
.B1(n_863),
.B2(n_788),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_816),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_896),
.A2(n_461),
.B(n_506),
.Y(n_950)
);

AOI22x1_ASAP7_75t_L g951 ( 
.A1(n_837),
.A2(n_569),
.B1(n_568),
.B2(n_559),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_850),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_782),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_SL g954 ( 
.A1(n_821),
.A2(n_546),
.B(n_568),
.C(n_559),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_767),
.A2(n_461),
.B(n_559),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_801),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_798),
.B(n_569),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_767),
.A2(n_461),
.B(n_558),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_783),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_799),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_743),
.B(n_569),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_799),
.A2(n_461),
.B(n_555),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_800),
.B(n_2),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_744),
.A2(n_558),
.B(n_555),
.C(n_554),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_785),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_890),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_792),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_783),
.B(n_436),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_890),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_799),
.A2(n_461),
.B(n_554),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_887),
.A2(n_555),
.B(n_554),
.C(n_546),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_789),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_754),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_858),
.A2(n_546),
.B(n_544),
.C(n_539),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_761),
.B(n_2),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_849),
.B(n_6),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_743),
.B(n_544),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_764),
.A2(n_544),
.B(n_539),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_856),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_751),
.A2(n_539),
.B1(n_434),
.B2(n_12),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_SL g981 ( 
.A1(n_894),
.A2(n_151),
.B(n_148),
.C(n_142),
.Y(n_981)
);

BUFx8_ASAP7_75t_SL g982 ( 
.A(n_834),
.Y(n_982)
);

NOR2x1_ASAP7_75t_SL g983 ( 
.A(n_878),
.B(n_139),
.Y(n_983)
);

BUFx4f_ASAP7_75t_L g984 ( 
.A(n_795),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_856),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_755),
.A2(n_10),
.B(n_13),
.C(n_15),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_749),
.A2(n_16),
.B1(n_20),
.B2(n_22),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_768),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_833),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_750),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_790),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_847),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_792),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_750),
.A2(n_29),
.B1(n_34),
.B2(n_37),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_809),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_824),
.A2(n_39),
.B(n_41),
.C(n_42),
.Y(n_996)
);

AO21x1_ASAP7_75t_L g997 ( 
.A1(n_753),
.A2(n_43),
.B(n_45),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_757),
.A2(n_43),
.B1(n_46),
.B2(n_68),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_SL g999 ( 
.A(n_852),
.B(n_78),
.C(n_80),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_839),
.B(n_879),
.Y(n_1000)
);

CKINVDCx11_ASAP7_75t_R g1001 ( 
.A(n_853),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_866),
.B(n_82),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_868),
.A2(n_823),
.B(n_869),
.C(n_861),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_866),
.A2(n_87),
.B1(n_93),
.B2(n_104),
.Y(n_1004)
);

O2A1O1Ixp5_ASAP7_75t_L g1005 ( 
.A1(n_897),
.A2(n_108),
.B(n_112),
.C(n_116),
.Y(n_1005)
);

AOI21xp33_ASAP7_75t_L g1006 ( 
.A1(n_860),
.A2(n_873),
.B(n_859),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_881),
.B(n_898),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_900),
.B(n_868),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_795),
.Y(n_1009)
);

AO32x1_ASAP7_75t_L g1010 ( 
.A1(n_848),
.A2(n_904),
.A3(n_903),
.B1(n_870),
.B2(n_864),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_885),
.A2(n_765),
.B(n_814),
.C(n_829),
.Y(n_1011)
);

INVx6_ASAP7_75t_L g1012 ( 
.A(n_793),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_793),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_757),
.B(n_747),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_883),
.B(n_910),
.Y(n_1015)
);

NAND3xp33_ASAP7_75t_L g1016 ( 
.A(n_852),
.B(n_893),
.C(n_882),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_813),
.A2(n_829),
.B(n_814),
.C(n_818),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_793),
.Y(n_1018)
);

AO21x1_ASAP7_75t_L g1019 ( 
.A1(n_902),
.A2(n_765),
.B(n_810),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_795),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_867),
.B(n_872),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_867),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_776),
.A2(n_891),
.B(n_871),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_747),
.B(n_748),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_810),
.A2(n_907),
.B(n_838),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_838),
.A2(n_830),
.B(n_831),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_830),
.A2(n_831),
.B(n_835),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_806),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_SL g1029 ( 
.A(n_826),
.B(n_875),
.C(n_874),
.Y(n_1029)
);

BUFx12f_ASAP7_75t_L g1030 ( 
.A(n_828),
.Y(n_1030)
);

OA22x2_ASAP7_75t_L g1031 ( 
.A1(n_826),
.A2(n_769),
.B1(n_813),
.B2(n_812),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_899),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_817),
.A2(n_779),
.B1(n_805),
.B2(n_766),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_772),
.B(n_774),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_960),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_919),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_931),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_915),
.B(n_748),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_955),
.A2(n_958),
.B(n_928),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_949),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1033),
.A2(n_841),
.B(n_851),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_950),
.A2(n_776),
.B(n_880),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_SL g1043 ( 
.A1(n_944),
.A2(n_840),
.B(n_791),
.Y(n_1043)
);

INVx6_ASAP7_75t_L g1044 ( 
.A(n_1030),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_959),
.B(n_895),
.Y(n_1045)
);

AOI221xp5_ASAP7_75t_SL g1046 ( 
.A1(n_987),
.A2(n_766),
.B1(n_808),
.B2(n_779),
.C(n_805),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_936),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_927),
.A2(n_880),
.B(n_835),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_1006),
.A2(n_808),
.B(n_778),
.C(n_796),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_925),
.B(n_857),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_937),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_1001),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_953),
.Y(n_1053)
);

AOI221x1_ASAP7_75t_L g1054 ( 
.A1(n_1006),
.A2(n_822),
.B1(n_820),
.B2(n_844),
.C(n_843),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_995),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_976),
.A2(n_909),
.B1(n_908),
.B2(n_906),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_SL g1057 ( 
.A1(n_935),
.A2(n_1003),
.B(n_1008),
.C(n_1014),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_1025),
.A2(n_877),
.B(n_756),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1027),
.A2(n_865),
.B(n_777),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1026),
.A2(n_756),
.B(n_777),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_1019),
.A2(n_877),
.A3(n_844),
.B(n_843),
.Y(n_1061)
);

OAI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_933),
.A2(n_803),
.B(n_862),
.Y(n_1062)
);

OA21x2_ASAP7_75t_L g1063 ( 
.A1(n_1023),
.A2(n_876),
.B(n_854),
.Y(n_1063)
);

AND2x2_ASAP7_75t_SL g1064 ( 
.A(n_984),
.B(n_905),
.Y(n_1064)
);

NOR2x1_ASAP7_75t_L g1065 ( 
.A(n_960),
.B(n_855),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_978),
.A2(n_901),
.B(n_807),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_917),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1007),
.B(n_1008),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_951),
.A2(n_1023),
.B(n_922),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1017),
.A2(n_1033),
.B(n_913),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_SL g1071 ( 
.A(n_1016),
.B(n_1015),
.C(n_963),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_1009),
.B(n_1020),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_926),
.B(n_918),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_989),
.A2(n_1031),
.B1(n_975),
.B2(n_999),
.Y(n_1074)
);

NAND2xp33_ASAP7_75t_L g1075 ( 
.A(n_1029),
.B(n_1007),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1024),
.A2(n_911),
.B(n_930),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_973),
.B(n_942),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_929),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_947),
.B(n_1022),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_997),
.A2(n_920),
.A3(n_964),
.B(n_974),
.Y(n_1080)
);

AOI221xp5_ASAP7_75t_L g1081 ( 
.A1(n_939),
.A2(n_912),
.B1(n_994),
.B2(n_987),
.C(n_990),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_924),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_911),
.A2(n_914),
.B(n_916),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1032),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1021),
.A2(n_932),
.B(n_954),
.Y(n_1085)
);

INVx5_ASAP7_75t_L g1086 ( 
.A(n_924),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_968),
.B(n_1034),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_981),
.A2(n_943),
.B(n_988),
.C(n_986),
.Y(n_1088)
);

O2A1O1Ixp5_ASAP7_75t_L g1089 ( 
.A1(n_1005),
.A2(n_961),
.B(n_977),
.C(n_946),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_992),
.Y(n_1090)
);

CKINVDCx14_ASAP7_75t_R g1091 ( 
.A(n_941),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1034),
.B(n_972),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1002),
.B(n_956),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1010),
.A2(n_971),
.B(n_921),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_1018),
.B(n_924),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_957),
.A2(n_1028),
.B(n_991),
.Y(n_1096)
);

NOR4xp25_ASAP7_75t_L g1097 ( 
.A(n_990),
.B(n_994),
.C(n_996),
.D(n_998),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1010),
.A2(n_970),
.B(n_962),
.Y(n_1098)
);

BUFx10_ASAP7_75t_L g1099 ( 
.A(n_952),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_965),
.B(n_1002),
.Y(n_1100)
);

INVxp67_ASAP7_75t_SL g1101 ( 
.A(n_966),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_SL g1102 ( 
.A1(n_948),
.A2(n_1004),
.B(n_980),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_984),
.A2(n_945),
.B(n_938),
.C(n_993),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_SL g1104 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_969),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_938),
.B(n_967),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_967),
.B(n_993),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1012),
.A2(n_979),
.B1(n_985),
.B2(n_1013),
.Y(n_1107)
);

INVxp67_ASAP7_75t_SL g1108 ( 
.A(n_966),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1012),
.A2(n_1013),
.B(n_966),
.Y(n_1109)
);

AO32x2_ASAP7_75t_L g1110 ( 
.A1(n_969),
.A2(n_1013),
.A3(n_940),
.B1(n_982),
.B2(n_934),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_969),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_919),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1000),
.B(n_815),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1000),
.B(n_815),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_SL g1115 ( 
.A1(n_944),
.A2(n_494),
.B(n_786),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_L g1116 ( 
.A(n_944),
.B(n_794),
.C(n_933),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1011),
.A2(n_832),
.B(n_815),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_944),
.A2(n_794),
.B(n_1006),
.C(n_933),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_960),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_976),
.A2(n_845),
.B1(n_815),
.B2(n_762),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_924),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1033),
.A2(n_620),
.B(n_598),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1000),
.B(n_815),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_960),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_924),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1027),
.A2(n_1026),
.B(n_797),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_955),
.A2(n_958),
.B(n_928),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1009),
.B(n_1020),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_919),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1009),
.B(n_1020),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_955),
.A2(n_958),
.B(n_928),
.Y(n_1131)
);

BUFx12f_ASAP7_75t_L g1132 ( 
.A(n_941),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_919),
.Y(n_1133)
);

INVx6_ASAP7_75t_L g1134 ( 
.A(n_949),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_915),
.B(n_545),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_955),
.A2(n_958),
.B(n_928),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_915),
.B(n_545),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_944),
.B(n_815),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_923),
.A2(n_794),
.B1(n_1000),
.B2(n_832),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_SL g1140 ( 
.A1(n_944),
.A2(n_781),
.B1(n_759),
.B2(n_514),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_955),
.A2(n_958),
.B(n_928),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_919),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1027),
.A2(n_1026),
.B(n_797),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1000),
.B(n_815),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1027),
.A2(n_1025),
.B(n_1026),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1027),
.A2(n_1026),
.B(n_797),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_919),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_1019),
.A2(n_997),
.A3(n_1026),
.B(n_1011),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1027),
.A2(n_1026),
.B(n_797),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1027),
.A2(n_1026),
.B(n_797),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_955),
.A2(n_958),
.B(n_928),
.Y(n_1151)
);

O2A1O1Ixp5_ASAP7_75t_L g1152 ( 
.A1(n_1019),
.A2(n_794),
.B(n_825),
.C(n_997),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1000),
.B(n_815),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1000),
.B(n_815),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_924),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_944),
.A2(n_794),
.B(n_1006),
.C(n_933),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_1019),
.A2(n_997),
.A3(n_1026),
.B(n_1011),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_919),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_955),
.A2(n_958),
.B(n_928),
.Y(n_1159)
);

OA21x2_ASAP7_75t_L g1160 ( 
.A1(n_1070),
.A2(n_1046),
.B(n_1145),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1051),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_1122),
.B(n_1117),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1055),
.Y(n_1163)
);

AO21x2_ASAP7_75t_L g1164 ( 
.A1(n_1041),
.A2(n_1143),
.B(n_1126),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1119),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1134),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1112),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1147),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1158),
.Y(n_1169)
);

AO21x1_ASAP7_75t_L g1170 ( 
.A1(n_1139),
.A2(n_1075),
.B(n_1074),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1136),
.A2(n_1151),
.B(n_1141),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1068),
.B(n_1138),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1036),
.Y(n_1173)
);

NOR2x1_ASAP7_75t_L g1174 ( 
.A(n_1113),
.B(n_1114),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1146),
.A2(n_1150),
.B(n_1149),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1046),
.A2(n_1094),
.B(n_1159),
.Y(n_1176)
);

BUFx2_ASAP7_75t_SL g1177 ( 
.A(n_1040),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1098),
.A2(n_1156),
.A3(n_1118),
.B(n_1083),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1053),
.Y(n_1179)
);

AO21x2_ASAP7_75t_L g1180 ( 
.A1(n_1085),
.A2(n_1069),
.B(n_1076),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1042),
.A2(n_1048),
.B(n_1060),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1093),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1058),
.A2(n_1059),
.B(n_1066),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1129),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1116),
.B(n_1043),
.Y(n_1185)
);

NAND2x1p5_ASAP7_75t_L g1186 ( 
.A(n_1086),
.B(n_1119),
.Y(n_1186)
);

INVxp67_ASAP7_75t_SL g1187 ( 
.A(n_1038),
.Y(n_1187)
);

AO21x2_ASAP7_75t_L g1188 ( 
.A1(n_1049),
.A2(n_1097),
.B(n_1088),
.Y(n_1188)
);

CKINVDCx11_ASAP7_75t_R g1189 ( 
.A(n_1132),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1072),
.B(n_1128),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1120),
.B(n_1045),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_1152),
.A2(n_1054),
.B(n_1062),
.Y(n_1192)
);

CKINVDCx11_ASAP7_75t_R g1193 ( 
.A(n_1099),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1133),
.Y(n_1194)
);

BUFx4f_ASAP7_75t_SL g1195 ( 
.A(n_1099),
.Y(n_1195)
);

INVx3_ASAP7_75t_SL g1196 ( 
.A(n_1037),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1063),
.A2(n_1089),
.B(n_1096),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1063),
.A2(n_1102),
.B(n_1065),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1047),
.Y(n_1199)
);

OAI222xp33_ASAP7_75t_L g1200 ( 
.A1(n_1120),
.A2(n_1077),
.B1(n_1154),
.B2(n_1153),
.C1(n_1123),
.C2(n_1144),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1135),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_1137),
.Y(n_1202)
);

NOR2xp67_ASAP7_75t_SL g1203 ( 
.A(n_1044),
.B(n_1052),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1109),
.A2(n_1062),
.B(n_1104),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1134),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1142),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1056),
.A2(n_1043),
.B(n_1124),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_1091),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1067),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1072),
.B(n_1130),
.Y(n_1210)
);

AOI22x1_ASAP7_75t_L g1211 ( 
.A1(n_1101),
.A2(n_1108),
.B1(n_1078),
.B2(n_1035),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1092),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1050),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1100),
.A2(n_1106),
.B(n_1095),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1071),
.A2(n_1079),
.B1(n_1064),
.B2(n_1130),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1111),
.A2(n_1105),
.B(n_1073),
.Y(n_1216)
);

NOR2xp67_ASAP7_75t_SL g1217 ( 
.A(n_1044),
.B(n_1115),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1148),
.A2(n_1157),
.B(n_1103),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1086),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1107),
.A2(n_1087),
.B(n_1080),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1107),
.A2(n_1080),
.B(n_1157),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1148),
.A2(n_1157),
.A3(n_1080),
.B(n_1097),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1148),
.A2(n_1061),
.A3(n_1057),
.B(n_1035),
.Y(n_1223)
);

INVx6_ASAP7_75t_L g1224 ( 
.A(n_1086),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1084),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1128),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1110),
.A2(n_1090),
.B(n_1082),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1110),
.A2(n_1082),
.B(n_1121),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1110),
.A2(n_1082),
.B(n_1121),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1125),
.A2(n_1159),
.B(n_1127),
.Y(n_1230)
);

INVx6_ASAP7_75t_SL g1231 ( 
.A(n_1125),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1155),
.Y(n_1232)
);

NAND3xp33_ASAP7_75t_L g1233 ( 
.A(n_1140),
.B(n_1116),
.C(n_1118),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1039),
.A2(n_1159),
.B(n_1131),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1116),
.A2(n_1156),
.B(n_1118),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1051),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1120),
.B(n_1045),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1051),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1116),
.B(n_1140),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1086),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1140),
.A2(n_1081),
.B1(n_1116),
.B2(n_845),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1145),
.A2(n_1143),
.B(n_1126),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1119),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1140),
.A2(n_1081),
.B1(n_1116),
.B2(n_845),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1120),
.B(n_1045),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1051),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1051),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1086),
.B(n_799),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1068),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1051),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1145),
.A2(n_1143),
.B(n_1126),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1072),
.B(n_1128),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1140),
.A2(n_1116),
.B1(n_1156),
.B2(n_1118),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1140),
.A2(n_781),
.B1(n_759),
.B2(n_1116),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1140),
.A2(n_1081),
.B1(n_1116),
.B2(n_845),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_SL g1256 ( 
.A1(n_1117),
.A2(n_997),
.B(n_983),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1135),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1116),
.B(n_1140),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1086),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1051),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1093),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1047),
.Y(n_1262)
);

OR2x6_ASAP7_75t_L g1263 ( 
.A(n_1122),
.B(n_1009),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1086),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1140),
.A2(n_1081),
.B1(n_1116),
.B2(n_845),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1051),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1140),
.A2(n_1081),
.B1(n_1116),
.B2(n_845),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1038),
.B(n_1113),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1051),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1051),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1116),
.B(n_1118),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1218),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1191),
.B(n_1237),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1254),
.A2(n_1255),
.B1(n_1267),
.B2(n_1265),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1189),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1242),
.A2(n_1251),
.B(n_1175),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1197),
.A2(n_1181),
.B(n_1235),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1241),
.A2(n_1265),
.B1(n_1255),
.B2(n_1267),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1189),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1249),
.B(n_1172),
.Y(n_1282)
);

NOR2x1_ASAP7_75t_SL g1283 ( 
.A(n_1162),
.B(n_1263),
.Y(n_1283)
);

O2A1O1Ixp5_ASAP7_75t_L g1284 ( 
.A1(n_1271),
.A2(n_1253),
.B(n_1170),
.C(n_1239),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1162),
.A2(n_1164),
.B(n_1271),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1241),
.A2(n_1244),
.B1(n_1215),
.B2(n_1239),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1208),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1187),
.B(n_1268),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1259),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1245),
.B(n_1182),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1291)
);

AOI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1217),
.A2(n_1256),
.B(n_1263),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1174),
.B(n_1212),
.Y(n_1293)
);

INVx8_ASAP7_75t_L g1294 ( 
.A(n_1205),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1197),
.A2(n_1181),
.B(n_1183),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1261),
.B(n_1252),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1252),
.B(n_1258),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1258),
.A2(n_1200),
.B(n_1233),
.C(n_1244),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1226),
.B(n_1215),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1185),
.B(n_1202),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1201),
.B(n_1185),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1185),
.B(n_1257),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1205),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_L g1304 ( 
.A(n_1199),
.B(n_1262),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1213),
.B(n_1270),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1225),
.A2(n_1162),
.B1(n_1195),
.B2(n_1211),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1228),
.B(n_1229),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1161),
.B(n_1163),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1208),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1193),
.Y(n_1310)
);

NOR2xp67_ASAP7_75t_L g1311 ( 
.A(n_1209),
.B(n_1167),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1168),
.B(n_1169),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1195),
.A2(n_1194),
.B1(n_1184),
.B2(n_1206),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1236),
.B(n_1238),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1228),
.B(n_1229),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1173),
.A2(n_1179),
.B1(n_1177),
.B2(n_1247),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1246),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1250),
.Y(n_1318)
);

NOR2x1_ASAP7_75t_SL g1319 ( 
.A(n_1263),
.B(n_1188),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1260),
.B(n_1269),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1266),
.A2(n_1224),
.B1(n_1227),
.B2(n_1166),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1227),
.B(n_1214),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1224),
.A2(n_1227),
.B1(n_1166),
.B2(n_1196),
.Y(n_1323)
);

AND2x6_ASAP7_75t_L g1324 ( 
.A(n_1165),
.B(n_1243),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1193),
.Y(n_1325)
);

BUFx12f_ASAP7_75t_L g1326 ( 
.A(n_1240),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1196),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1186),
.A2(n_1219),
.B1(n_1264),
.B2(n_1240),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1186),
.A2(n_1219),
.B1(n_1264),
.B2(n_1232),
.Y(n_1329)
);

BUFx4f_ASAP7_75t_SL g1330 ( 
.A(n_1231),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1214),
.B(n_1178),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1178),
.B(n_1220),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1207),
.A2(n_1221),
.B(n_1220),
.C(n_1198),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1178),
.B(n_1222),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1216),
.B(n_1165),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1165),
.A2(n_1243),
.B1(n_1192),
.B2(n_1248),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1222),
.B(n_1160),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1204),
.B(n_1198),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1222),
.B(n_1203),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1222),
.B(n_1160),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1183),
.A2(n_1171),
.B(n_1234),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1223),
.B(n_1176),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1223),
.B(n_1180),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1176),
.B(n_1230),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1171),
.B(n_1234),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1307),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1288),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1307),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1298),
.A2(n_1279),
.B(n_1275),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1301),
.B(n_1339),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1286),
.A2(n_1298),
.B1(n_1282),
.B2(n_1293),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1334),
.B(n_1331),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1333),
.A2(n_1285),
.B(n_1337),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1322),
.B(n_1302),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1315),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1311),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1296),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1285),
.A2(n_1340),
.B(n_1343),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1272),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1272),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1315),
.B(n_1338),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1273),
.B(n_1290),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1316),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1335),
.B(n_1297),
.Y(n_1364)
);

BUFx12f_ASAP7_75t_L g1365 ( 
.A(n_1310),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1300),
.B(n_1318),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1300),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1317),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1338),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1305),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1313),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1304),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1314),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1320),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1287),
.A2(n_1309),
.B1(n_1327),
.B2(n_1299),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1321),
.B(n_1332),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1345),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1342),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1323),
.B(n_1308),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1278),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1324),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1312),
.B(n_1319),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1278),
.B(n_1344),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1295),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1336),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1278),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1287),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1295),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1284),
.B(n_1277),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1306),
.A2(n_1274),
.B1(n_1280),
.B2(n_1291),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1284),
.B(n_1277),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1283),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1383),
.B(n_1277),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1383),
.B(n_1295),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1369),
.B(n_1292),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1384),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1370),
.B(n_1324),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1359),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1384),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1361),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1370),
.B(n_1373),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1378),
.B(n_1352),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1359),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1352),
.B(n_1341),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1360),
.Y(n_1406)
);

INVxp67_ASAP7_75t_R g1407 ( 
.A(n_1389),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1388),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1369),
.B(n_1361),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1361),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1356),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1358),
.B(n_1329),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1387),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1369),
.B(n_1324),
.Y(n_1414)
);

INVx4_ASAP7_75t_L g1415 ( 
.A(n_1381),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1351),
.A2(n_1309),
.B1(n_1281),
.B2(n_1276),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1416),
.A2(n_1349),
.B1(n_1351),
.B2(n_1371),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_SL g1418 ( 
.A(n_1416),
.B(n_1375),
.C(n_1281),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1400),
.B(n_1376),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1412),
.A2(n_1349),
.B(n_1375),
.C(n_1363),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1407),
.B(n_1354),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1409),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1412),
.B(n_1372),
.C(n_1391),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1415),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1407),
.B(n_1354),
.Y(n_1425)
);

OAI221xp5_ASAP7_75t_L g1426 ( 
.A1(n_1411),
.A2(n_1390),
.B1(n_1392),
.B2(n_1366),
.C(n_1379),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1398),
.Y(n_1427)
);

INVx4_ASAP7_75t_L g1428 ( 
.A(n_1415),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1398),
.Y(n_1429)
);

AOI222xp33_ASAP7_75t_L g1430 ( 
.A1(n_1411),
.A2(n_1391),
.B1(n_1389),
.B2(n_1366),
.C1(n_1347),
.C2(n_1379),
.Y(n_1430)
);

OAI221xp5_ASAP7_75t_L g1431 ( 
.A1(n_1397),
.A2(n_1392),
.B1(n_1367),
.B2(n_1382),
.C(n_1385),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1403),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1414),
.B(n_1381),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1403),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1415),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1402),
.B(n_1377),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1407),
.B(n_1350),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1396),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1413),
.A2(n_1276),
.B1(n_1357),
.B2(n_1376),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1406),
.Y(n_1440)
);

OAI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1397),
.A2(n_1382),
.B1(n_1385),
.B2(n_1368),
.C(n_1376),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1404),
.A2(n_1368),
.B1(n_1374),
.B2(n_1362),
.C(n_1364),
.Y(n_1442)
);

OAI221xp5_ASAP7_75t_L g1443 ( 
.A1(n_1412),
.A2(n_1376),
.B1(n_1355),
.B2(n_1348),
.C(n_1346),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1402),
.Y(n_1444)
);

INVxp67_ASAP7_75t_SL g1445 ( 
.A(n_1401),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1401),
.B(n_1364),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1396),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1399),
.A2(n_1386),
.B(n_1380),
.Y(n_1448)
);

OAI221xp5_ASAP7_75t_L g1449 ( 
.A1(n_1400),
.A2(n_1376),
.B1(n_1348),
.B2(n_1355),
.C(n_1346),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1400),
.B(n_1350),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1402),
.B(n_1377),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1409),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1413),
.A2(n_1376),
.B1(n_1328),
.B2(n_1362),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1427),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1448),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1448),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1429),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1448),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1427),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1432),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1432),
.Y(n_1461)
);

NOR3xp33_ASAP7_75t_L g1462 ( 
.A(n_1417),
.B(n_1325),
.C(n_1415),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1423),
.A2(n_1380),
.B(n_1408),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1448),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1438),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1452),
.B(n_1394),
.Y(n_1466)
);

INVx4_ASAP7_75t_L g1467 ( 
.A(n_1428),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1424),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1438),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1424),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1445),
.B(n_1394),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1423),
.B(n_1405),
.Y(n_1472)
);

INVx4_ASAP7_75t_SL g1473 ( 
.A(n_1424),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1438),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1420),
.B(n_1414),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_L g1476 ( 
.A(n_1430),
.B(n_1404),
.C(n_1353),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1447),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1447),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1444),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1435),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1434),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1473),
.B(n_1452),
.Y(n_1482)
);

AND2x2_ASAP7_75t_SL g1483 ( 
.A(n_1462),
.B(n_1428),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1468),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1467),
.B(n_1428),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1476),
.B(n_1442),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1467),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1476),
.B(n_1450),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1468),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1454),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1457),
.B(n_1450),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1465),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1471),
.B(n_1446),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1454),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1457),
.B(n_1431),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1462),
.A2(n_1426),
.B1(n_1418),
.B2(n_1441),
.C(n_1449),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1471),
.B(n_1436),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1459),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1479),
.B(n_1453),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1459),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1479),
.B(n_1453),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1460),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1475),
.B(n_1421),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1472),
.B(n_1436),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1473),
.B(n_1437),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1460),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1463),
.B(n_1439),
.C(n_1443),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1473),
.B(n_1437),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1473),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1467),
.B(n_1365),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1472),
.B(n_1451),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1481),
.B(n_1421),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1473),
.B(n_1422),
.Y(n_1513)
);

NAND2xp33_ASAP7_75t_R g1514 ( 
.A(n_1463),
.B(n_1303),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1472),
.B(n_1451),
.Y(n_1515)
);

NAND2x1p5_ASAP7_75t_L g1516 ( 
.A(n_1467),
.B(n_1428),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1465),
.Y(n_1517)
);

AOI211xp5_ASAP7_75t_L g1518 ( 
.A1(n_1470),
.A2(n_1439),
.B(n_1433),
.C(n_1435),
.Y(n_1518)
);

NAND4xp25_ASAP7_75t_L g1519 ( 
.A(n_1467),
.B(n_1435),
.C(n_1415),
.D(n_1395),
.Y(n_1519)
);

AND2x4_ASAP7_75t_SL g1520 ( 
.A(n_1481),
.B(n_1414),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1470),
.B(n_1425),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1465),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1463),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1505),
.B(n_1473),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1486),
.B(n_1470),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1505),
.B(n_1480),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1508),
.B(n_1480),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1484),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1508),
.B(n_1480),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1482),
.B(n_1466),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1490),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1489),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1494),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1495),
.A2(n_1463),
.B(n_1419),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1499),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1483),
.B(n_1365),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1498),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1488),
.B(n_1461),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1496),
.B(n_1461),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1492),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1482),
.B(n_1466),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1492),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1518),
.A2(n_1393),
.B(n_1410),
.C(n_1464),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1500),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1501),
.B(n_1466),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1520),
.B(n_1422),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1502),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1506),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1510),
.B(n_1365),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1493),
.B(n_1463),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1517),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1510),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1491),
.B(n_1425),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1483),
.B(n_1294),
.Y(n_1554)
);

NAND2x1p5_ASAP7_75t_L g1555 ( 
.A(n_1487),
.B(n_1381),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1512),
.B(n_1440),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1520),
.B(n_1422),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1513),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1532),
.B(n_1503),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1536),
.B(n_1487),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1528),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1524),
.B(n_1487),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1524),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1558),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1558),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1526),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1535),
.B(n_1521),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1526),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1531),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1531),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1533),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1525),
.B(n_1504),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1538),
.B(n_1504),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1539),
.A2(n_1507),
.B1(n_1509),
.B2(n_1419),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1527),
.B(n_1513),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1527),
.B(n_1485),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1538),
.B(n_1545),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1529),
.B(n_1485),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1533),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1529),
.Y(n_1580)
);

OAI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1534),
.A2(n_1514),
.B1(n_1519),
.B2(n_1419),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1555),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1555),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1564),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1564),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1561),
.B(n_1552),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1565),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1565),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1566),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1563),
.B(n_1549),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1572),
.B(n_1556),
.Y(n_1591)
);

AOI222xp33_ASAP7_75t_L g1592 ( 
.A1(n_1574),
.A2(n_1543),
.B1(n_1554),
.B2(n_1523),
.C1(n_1547),
.C2(n_1544),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1580),
.Y(n_1593)
);

NOR3xp33_ASAP7_75t_L g1594 ( 
.A(n_1559),
.B(n_1523),
.C(n_1547),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1568),
.B(n_1567),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1581),
.A2(n_1516),
.B(n_1553),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1569),
.Y(n_1597)
);

AOI21xp33_ASAP7_75t_L g1598 ( 
.A1(n_1560),
.A2(n_1514),
.B(n_1544),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1575),
.A2(n_1530),
.B1(n_1541),
.B2(n_1516),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1562),
.B(n_1530),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1570),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1572),
.A2(n_1548),
.B1(n_1537),
.B2(n_1541),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1589),
.B(n_1577),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1585),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1584),
.B(n_1562),
.Y(n_1605)
);

NOR2x1_ASAP7_75t_L g1606 ( 
.A(n_1587),
.B(n_1583),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1588),
.B(n_1586),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1586),
.B(n_1577),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1600),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1590),
.B(n_1562),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1593),
.B(n_1575),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1598),
.A2(n_1575),
.B1(n_1576),
.B2(n_1578),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1608),
.A2(n_1609),
.B1(n_1607),
.B2(n_1602),
.C(n_1612),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1604),
.A2(n_1602),
.B1(n_1594),
.B2(n_1605),
.C(n_1595),
.Y(n_1614)
);

NOR3xp33_ASAP7_75t_L g1615 ( 
.A(n_1610),
.B(n_1601),
.C(n_1597),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1611),
.B(n_1591),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1603),
.A2(n_1599),
.B1(n_1596),
.B2(n_1573),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1606),
.B(n_1573),
.Y(n_1618)
);

NAND2xp33_ASAP7_75t_L g1619 ( 
.A(n_1606),
.B(n_1594),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1605),
.B(n_1571),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1605),
.B(n_1579),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1613),
.A2(n_1614),
.B1(n_1619),
.B2(n_1618),
.C(n_1617),
.Y(n_1622)
);

AOI31xp33_ASAP7_75t_L g1623 ( 
.A1(n_1616),
.A2(n_1592),
.A3(n_1576),
.B(n_1578),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1615),
.B(n_1582),
.Y(n_1624)
);

OAI21xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1620),
.A2(n_1583),
.B(n_1550),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1621),
.A2(n_1583),
.B1(n_1523),
.B2(n_1548),
.C(n_1537),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1624),
.Y(n_1627)
);

NAND2xp33_ASAP7_75t_SL g1628 ( 
.A(n_1623),
.B(n_1550),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1625),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1626),
.Y(n_1630)
);

OAI21xp33_ASAP7_75t_L g1631 ( 
.A1(n_1622),
.A2(n_1555),
.B(n_1551),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1624),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1629),
.B(n_1546),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1627),
.Y(n_1634)
);

OAI322xp33_ASAP7_75t_L g1635 ( 
.A1(n_1630),
.A2(n_1551),
.A3(n_1542),
.B1(n_1540),
.B2(n_1515),
.C1(n_1511),
.C2(n_1455),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1628),
.A2(n_1542),
.B1(n_1540),
.B2(n_1511),
.C(n_1515),
.Y(n_1636)
);

OAI21xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1629),
.A2(n_1557),
.B(n_1546),
.Y(n_1637)
);

INVxp33_ASAP7_75t_L g1638 ( 
.A(n_1633),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1634),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1637),
.B(n_1632),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1640),
.B(n_1631),
.C(n_1636),
.Y(n_1641)
);

OAI322xp33_ASAP7_75t_L g1642 ( 
.A1(n_1641),
.A2(n_1639),
.A3(n_1638),
.B1(n_1635),
.B2(n_1456),
.C1(n_1455),
.C2(n_1458),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1642),
.A2(n_1638),
.B1(n_1517),
.B2(n_1522),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1643),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1644),
.A2(n_1557),
.B1(n_1294),
.B2(n_1522),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1645),
.A2(n_1464),
.B(n_1458),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1645),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1647),
.A2(n_1294),
.B1(n_1330),
.B2(n_1456),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1646),
.A2(n_1497),
.B(n_1455),
.Y(n_1649)
);

OAI222xp33_ASAP7_75t_L g1650 ( 
.A1(n_1648),
.A2(n_1646),
.B1(n_1330),
.B2(n_1458),
.C1(n_1464),
.C2(n_1456),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1649),
.B(n_1469),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1651),
.Y(n_1652)
);

AOI22x1_ASAP7_75t_L g1653 ( 
.A1(n_1650),
.A2(n_1326),
.B1(n_1289),
.B2(n_1474),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1652),
.A2(n_1478),
.B1(n_1474),
.B2(n_1477),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1654),
.A2(n_1653),
.B1(n_1469),
.B2(n_1478),
.Y(n_1655)
);


endmodule