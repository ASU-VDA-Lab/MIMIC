module fake_jpeg_26877_n_383 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_383);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_383;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_38),
.Y(n_97)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_53),
.Y(n_83)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_52),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_13),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_13),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_12),
.Y(n_89)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_19),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_13),
.C(n_12),
.Y(n_88)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_22),
.B1(n_36),
.B2(n_18),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_86),
.B1(n_90),
.B2(n_96),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_68),
.B(n_84),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_17),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_21),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_17),
.B1(n_35),
.B2(n_31),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_89),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_40),
.A2(n_17),
.B1(n_35),
.B2(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_18),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_95),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_43),
.A2(n_18),
.B1(n_35),
.B2(n_31),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_101),
.Y(n_127)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_36),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_26),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_106),
.B(n_111),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_16),
.B1(n_20),
.B2(n_26),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_109),
.B(n_116),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_48),
.B1(n_55),
.B2(n_58),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_137),
.B1(n_144),
.B2(n_33),
.Y(n_152)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_53),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_133),
.C(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_26),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_24),
.Y(n_161)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_73),
.A2(n_19),
.B(n_21),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_33),
.B(n_28),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_39),
.B1(n_47),
.B2(n_44),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_132),
.B1(n_138),
.B2(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_128),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_69),
.Y(n_175)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_30),
.B1(n_36),
.B2(n_27),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_0),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_30),
.C(n_28),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_92),
.A2(n_33),
.B1(n_28),
.B2(n_24),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_140),
.B1(n_74),
.B2(n_70),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_71),
.A2(n_27),
.B1(n_20),
.B2(n_16),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_71),
.A2(n_97),
.B1(n_75),
.B2(n_92),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_94),
.B1(n_79),
.B2(n_93),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_93),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_141),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_75),
.A2(n_85),
.B1(n_94),
.B2(n_104),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_82),
.A2(n_16),
.B1(n_27),
.B2(n_20),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_106),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_153),
.B1(n_163),
.B2(n_136),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_79),
.B1(n_76),
.B2(n_87),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_111),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_156),
.B(n_162),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_170),
.B(n_179),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_81),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_158),
.B(n_161),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_159),
.Y(n_209)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_79),
.B1(n_87),
.B2(n_76),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_164),
.B(n_166),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_167),
.A2(n_122),
.B1(n_110),
.B2(n_121),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_103),
.C(n_93),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_175),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_141),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_103),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_87),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_127),
.B(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_132),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_117),
.B(n_76),
.C(n_78),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_166),
.A2(n_109),
.B1(n_116),
.B2(n_134),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_188),
.B1(n_211),
.B2(n_214),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_184),
.B(n_195),
.Y(n_233)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_193),
.Y(n_246)
);

OR2x2_ASAP7_75t_SL g187 ( 
.A(n_178),
.B(n_135),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_187),
.A2(n_198),
.B(n_202),
.Y(n_229)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_115),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_194),
.Y(n_230)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_115),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_196),
.B(n_11),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_142),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_133),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_207),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_124),
.B(n_133),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_147),
.B(n_150),
.Y(n_228)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_139),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_108),
.Y(n_206)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_129),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_218),
.B1(n_174),
.B2(n_145),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_162),
.A2(n_154),
.B1(n_156),
.B2(n_171),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_154),
.A2(n_113),
.B1(n_131),
.B2(n_112),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_159),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_215),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_170),
.A2(n_110),
.B1(n_78),
.B2(n_124),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_147),
.B1(n_150),
.B2(n_169),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_24),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_10),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_176),
.B1(n_168),
.B2(n_180),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_160),
.C(n_176),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_217),
.C(n_203),
.Y(n_264)
);

OAI32xp33_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_173),
.A3(n_164),
.B1(n_157),
.B2(n_145),
.Y(n_220)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_183),
.B1(n_207),
.B2(n_184),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_158),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_231),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_181),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_227),
.B(n_241),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_SL g262 ( 
.A1(n_228),
.A2(n_233),
.B(n_209),
.C(n_241),
.Y(n_262)
);

INVx4_ASAP7_75t_SL g231 ( 
.A(n_210),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_245),
.B1(n_196),
.B2(n_209),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_182),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_234),
.Y(n_267)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_30),
.B(n_172),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_187),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_169),
.B1(n_142),
.B2(n_139),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_243),
.B1(n_185),
.B2(n_208),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_142),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_252),
.Y(n_270)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_195),
.A2(n_139),
.B1(n_12),
.B2(n_11),
.Y(n_243)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_191),
.B(n_10),
.CI(n_1),
.CON(n_248),
.SN(n_248)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_213),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_194),
.B(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_1),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_1),
.Y(n_253)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_280),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_212),
.B1(n_215),
.B2(n_199),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_256),
.A2(n_258),
.B1(n_271),
.B2(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_259),
.B(n_250),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g287 ( 
.A1(n_262),
.A2(n_272),
.B(n_228),
.C(n_220),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_268),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_276),
.C(n_219),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_224),
.A2(n_202),
.B1(n_210),
.B2(n_213),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_275),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_224),
.A2(n_201),
.B1(n_193),
.B2(n_192),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_189),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_236),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_237),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_221),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_281),
.Y(n_293)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_229),
.B(n_228),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_284),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_229),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_285),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_290),
.C(n_255),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_299),
.B(n_262),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_288),
.A2(n_263),
.B1(n_279),
.B2(n_249),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_230),
.C(n_244),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_223),
.B(n_244),
.C(n_230),
.D(n_248),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_297),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_296),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_271),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_243),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_256),
.B(n_226),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_302),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_231),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_277),
.B(n_253),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_242),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_305),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_266),
.B(n_232),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_284),
.B(n_270),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_257),
.C(n_265),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_312),
.C(n_313),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_265),
.C(n_278),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_278),
.C(n_261),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_254),
.C(n_252),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_317),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_315),
.A2(n_319),
.B1(n_6),
.B2(n_7),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_258),
.B1(n_239),
.B2(n_248),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_275),
.C(n_280),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_298),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_225),
.B1(n_235),
.B2(n_8),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_SL g326 ( 
.A(n_308),
.B(n_291),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_326),
.B(n_327),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_292),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_333),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_308),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_331),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_282),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_303),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_298),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_334),
.B(n_338),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_321),
.A2(n_293),
.B(n_299),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_336),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_321),
.A2(n_287),
.B1(n_283),
.B2(n_235),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_337),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_294),
.Y(n_338)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_339),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_326),
.A2(n_316),
.B1(n_320),
.B2(n_325),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_324),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_337),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_353),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_318),
.B(n_314),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_349),
.A2(n_351),
.B(n_330),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_350),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_340),
.A2(n_331),
.B(n_338),
.Y(n_351)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_329),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_354),
.A2(n_360),
.B(n_8),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_344),
.B(n_322),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_355),
.B(n_359),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_323),
.Y(n_356)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_357),
.B(n_347),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_332),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_352),
.B(n_329),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_343),
.C(n_345),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_8),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_7),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_9),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_366),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_361),
.A2(n_345),
.B(n_8),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_362),
.B(n_7),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_367),
.B(n_369),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_368),
.A2(n_354),
.B1(n_358),
.B2(n_9),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_9),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_376),
.Y(n_378)
);

FAx1_ASAP7_75t_SL g375 ( 
.A(n_371),
.B(n_363),
.CI(n_364),
.CON(n_375),
.SN(n_375)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_375),
.B(n_367),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_377),
.A2(n_379),
.B(n_370),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_373),
.B(n_365),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_380),
.A2(n_374),
.B1(n_378),
.B2(n_376),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_375),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_9),
.Y(n_383)
);


endmodule