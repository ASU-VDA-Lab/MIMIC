module fake_jpeg_8234_n_249 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_14),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_43),
.Y(n_46)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_42),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_52),
.Y(n_68)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_33),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_24),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_28),
.B(n_26),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_34),
.B1(n_31),
.B2(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_65),
.B1(n_31),
.B2(n_18),
.Y(n_77)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_36),
.Y(n_78)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_34),
.B1(n_31),
.B2(n_26),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_71),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_69),
.B(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_80),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_86),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_42),
.B1(n_39),
.B2(n_50),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_42),
.B1(n_39),
.B2(n_29),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_38),
.C(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_25),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_44),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_89),
.Y(n_121)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_38),
.B(n_24),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_28),
.B(n_49),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_112),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_68),
.B(n_72),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_82),
.B1(n_96),
.B2(n_83),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_0),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_30),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_42),
.B1(n_39),
.B2(n_32),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_115),
.A2(n_123),
.B1(n_84),
.B2(n_83),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_74),
.B1(n_93),
.B2(n_84),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_23),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_67),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_79),
.A2(n_32),
.B1(n_21),
.B2(n_29),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_125),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_137),
.B(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_67),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_145),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_108),
.B(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_70),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_136),
.B(n_138),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_100),
.B1(n_72),
.B2(n_68),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_76),
.C(n_81),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_143),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_144),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_27),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_70),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_94),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_22),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_152),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_106),
.B1(n_118),
.B2(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_141),
.B1(n_151),
.B2(n_150),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_163),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_171),
.C(n_142),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_164),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_132),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_125),
.C(n_111),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_111),
.B(n_125),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_172),
.B1(n_156),
.B2(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_148),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_122),
.B(n_105),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_131),
.A2(n_122),
.B(n_105),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_107),
.B(n_124),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_127),
.A2(n_145),
.B(n_130),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_66),
.Y(n_183)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_181),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_1),
.B(n_2),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_170),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_152),
.A3(n_138),
.B1(n_107),
.B2(n_144),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_161),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_160),
.B(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_186),
.B1(n_188),
.B2(n_174),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_103),
.B1(n_96),
.B2(n_124),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_185),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_197)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_27),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_103),
.B1(n_92),
.B2(n_25),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_16),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_191),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_157),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_23),
.B1(n_21),
.B2(n_32),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_153),
.A2(n_17),
.B1(n_30),
.B2(n_22),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_166),
.A3(n_153),
.B1(n_163),
.B2(n_154),
.C1(n_161),
.C2(n_174),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_183),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_206),
.B1(n_1),
.B2(n_4),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_176),
.C(n_158),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_205),
.C(n_208),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_172),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_30),
.B1(n_15),
.B2(n_13),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_30),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_209),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_12),
.C(n_2),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_4),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_218),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_186),
.B(n_185),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_219),
.B1(n_221),
.B2(n_210),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_194),
.C(n_182),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_4),
.C(n_5),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_190),
.C(n_193),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_1),
.B(n_3),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_6),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_209),
.B1(n_202),
.B2(n_197),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_208),
.C(n_200),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_225),
.C(n_230),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_207),
.C(n_197),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_227),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_6),
.C(n_7),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_216),
.B1(n_218),
.B2(n_217),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_219),
.B(n_213),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_217),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_213),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_238),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_8),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_236),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_9),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_241),
.A2(n_236),
.B1(n_10),
.B2(n_11),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_239),
.Y(n_246)
);

OAI21x1_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_245),
.B(n_243),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_234),
.C(n_9),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_10),
.Y(n_249)
);


endmodule