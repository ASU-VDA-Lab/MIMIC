module fake_jpeg_12453_n_482 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_482);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_482;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_47),
.Y(n_137)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_51),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_53),
.B(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_55),
.Y(n_148)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_57),
.Y(n_128)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_24),
.Y(n_58)
);

CKINVDCx12_ASAP7_75t_R g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_60),
.Y(n_115)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_33),
.B(n_0),
.CON(n_64),
.SN(n_64)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_71),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_0),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_18),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_80),
.B(n_86),
.Y(n_141)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

CKINVDCx9p33_ASAP7_75t_R g83 ( 
.A(n_33),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_89),
.Y(n_110)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_90),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_44),
.B1(n_25),
.B2(n_18),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_101),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_44),
.B1(n_35),
.B2(n_30),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_103),
.A2(n_108),
.B1(n_114),
.B2(n_127),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_45),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_105),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_40),
.B1(n_30),
.B2(n_22),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_106),
.A2(n_116),
.B1(n_42),
.B2(n_28),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_44),
.B1(n_35),
.B2(n_30),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_38),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_111),
.B(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_76),
.B(n_26),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_59),
.A2(n_35),
.B1(n_22),
.B2(n_40),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_57),
.A2(n_22),
.B1(n_35),
.B2(n_37),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_34),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_117),
.B(n_118),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_61),
.C(n_37),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_36),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_124),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_36),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_25),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_129),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_62),
.A2(n_38),
.B1(n_26),
.B2(n_42),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_46),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_46),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_130),
.A2(n_12),
.B(n_14),
.C(n_95),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_48),
.B(n_46),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_56),
.B(n_43),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_84),
.B(n_43),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_10),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_63),
.A2(n_43),
.B1(n_42),
.B2(n_28),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_149),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_141),
.A2(n_73),
.B1(n_85),
.B2(n_87),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_150),
.A2(n_151),
.B1(n_166),
.B2(n_107),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_155),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_60),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_156),
.B(n_190),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_97),
.A2(n_28),
.B1(n_27),
.B2(n_68),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_159),
.A2(n_188),
.B(n_191),
.Y(n_228)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_97),
.A2(n_27),
.B(n_1),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_161),
.A2(n_99),
.B(n_98),
.Y(n_223)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_136),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_162),
.B(n_185),
.Y(n_213)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_168),
.A2(n_194),
.B1(n_196),
.B2(n_201),
.Y(n_216)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_97),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_204),
.Y(n_210)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_109),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_178),
.Y(n_207)
);

BUFx4f_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_174),
.Y(n_253)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_175),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_103),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_176),
.A2(n_131),
.B1(n_143),
.B2(n_94),
.Y(n_218)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_93),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_179),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_110),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_184),
.Y(n_211)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_105),
.B(n_6),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_195),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_96),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_193),
.B(n_198),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_114),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_92),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_96),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_120),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_200),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_105),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_108),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_202),
.A2(n_122),
.B(n_133),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_205),
.Y(n_251)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_131),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_187),
.A2(n_104),
.B1(n_94),
.B2(n_144),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_209),
.A2(n_224),
.B1(n_235),
.B2(n_242),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_218),
.B(n_222),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_156),
.A2(n_143),
.B(n_142),
.C(n_131),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g284 ( 
.A1(n_219),
.A2(n_245),
.B(n_172),
.C(n_233),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_171),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_178),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_223),
.A2(n_186),
.B(n_203),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_144),
.B1(n_102),
.B2(n_119),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_225),
.A2(n_234),
.B1(n_239),
.B2(n_250),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_174),
.B(n_100),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_233),
.B(n_222),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_150),
.A2(n_107),
.B1(n_102),
.B2(n_113),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_119),
.B1(n_146),
.B2(n_145),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_142),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_153),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_151),
.A2(n_146),
.B1(n_145),
.B2(n_100),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_184),
.A2(n_140),
.B1(n_145),
.B2(n_146),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_241),
.A2(n_154),
.B1(n_205),
.B2(n_167),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_199),
.A2(n_99),
.B1(n_98),
.B2(n_91),
.Y(n_242)
);

AOI32xp33_ASAP7_75t_L g245 ( 
.A1(n_188),
.A2(n_158),
.A3(n_152),
.B1(n_206),
.B2(n_192),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_173),
.B(n_133),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_257),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_169),
.A2(n_91),
.B1(n_122),
.B2(n_134),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_191),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_201),
.A2(n_159),
.B1(n_193),
.B2(n_185),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_254),
.A2(n_224),
.B1(n_235),
.B2(n_216),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_183),
.A2(n_133),
.B1(n_204),
.B2(n_191),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_255),
.A2(n_248),
.B1(n_230),
.B2(n_231),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_165),
.B(n_133),
.C(n_161),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_238),
.B(n_169),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_260),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_261),
.B(n_265),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_262),
.A2(n_270),
.B(n_273),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_229),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_266),
.Y(n_325)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_175),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_213),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_225),
.A2(n_160),
.B1(n_195),
.B2(n_191),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_267),
.A2(n_276),
.B1(n_302),
.B2(n_303),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_268),
.A2(n_295),
.B(n_246),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_207),
.B(n_177),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_269),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_155),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_272),
.B(n_281),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_210),
.B(n_163),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_277),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_164),
.C(n_170),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_275),
.B(n_208),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_227),
.A2(n_182),
.B1(n_181),
.B2(n_162),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_210),
.B(n_172),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_232),
.Y(n_278)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_213),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_212),
.Y(n_282)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_237),
.Y(n_283)
);

INVx3_ASAP7_75t_SL g330 ( 
.A(n_283),
.Y(n_330)
);

O2A1O1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_284),
.A2(n_292),
.B(n_301),
.C(n_280),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_249),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_288),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_209),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_292),
.Y(n_306)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_236),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_242),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_251),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_294),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_227),
.A2(n_223),
.B(n_219),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_254),
.A2(n_252),
.B1(n_228),
.B2(n_239),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_301),
.B1(n_208),
.B2(n_246),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_214),
.B(n_240),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_297),
.B(n_299),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_215),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_293),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_236),
.B(n_244),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_250),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_300),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_228),
.A2(n_245),
.B1(n_248),
.B2(n_218),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_231),
.A2(n_237),
.B1(n_244),
.B2(n_230),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_277),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_317),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_311),
.A2(n_338),
.B(n_296),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_340),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_217),
.B1(n_220),
.B2(n_243),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_217),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_315),
.Y(n_353)
);

AND2x6_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_271),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_295),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_320),
.B(n_333),
.Y(n_367)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_243),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_323),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_220),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_327),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_220),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_259),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_267),
.A2(n_298),
.B1(n_276),
.B2(n_273),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_303),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_268),
.A2(n_273),
.B(n_286),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_260),
.B(n_270),
.Y(n_339)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_281),
.A2(n_279),
.B(n_278),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_342),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_290),
.A2(n_302),
.B1(n_285),
.B2(n_294),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_343),
.A2(n_285),
.B1(n_290),
.B2(n_266),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_323),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_344),
.B(n_346),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_342),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_347),
.A2(n_307),
.B(n_340),
.Y(n_380)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_350),
.C(n_357),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_275),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_352),
.A2(n_362),
.B1(n_327),
.B2(n_306),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_329),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_304),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_376),
.Y(n_389)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_275),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_366),
.C(n_373),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_343),
.A2(n_262),
.B1(n_258),
.B2(n_264),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_291),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_324),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_368),
.B(n_371),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_311),
.A2(n_263),
.B(n_282),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_369),
.A2(n_307),
.B(n_315),
.Y(n_377)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_372),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_325),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_319),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_314),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_314),
.B(n_288),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_320),
.C(n_322),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_315),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_377),
.A2(n_380),
.B(n_391),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_367),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_382),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_364),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_383),
.A2(n_386),
.B1(n_390),
.B2(n_363),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_364),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_395),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_308),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_388),
.B(n_393),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_358),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_351),
.A2(n_312),
.B1(n_318),
.B2(n_333),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_332),
.C(n_317),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_396),
.C(n_401),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_345),
.B(n_324),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_341),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_332),
.C(n_321),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_345),
.B(n_335),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_400),
.B(n_375),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_306),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_351),
.A2(n_318),
.B1(n_337),
.B2(n_310),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_402),
.A2(n_362),
.B1(n_353),
.B2(n_352),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_403),
.A2(n_337),
.B1(n_305),
.B2(n_354),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_403),
.A2(n_356),
.B1(n_376),
.B2(n_353),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_404),
.A2(n_387),
.B1(n_391),
.B2(n_369),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_389),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_410),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_355),
.Y(n_407)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_407),
.Y(n_426)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_398),
.Y(n_409)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_409),
.Y(n_436)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_389),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_366),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_416),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_413),
.A2(n_420),
.B1(n_424),
.B2(n_326),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_381),
.B(n_355),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_411),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g415 ( 
.A1(n_383),
.A2(n_356),
.B(n_354),
.C(n_375),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_415),
.A2(n_380),
.B(n_377),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_374),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_402),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_397),
.A2(n_305),
.B1(n_347),
.B2(n_358),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_384),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_421),
.B(n_399),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_386),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_375),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_394),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_428),
.A2(n_434),
.B1(n_413),
.B2(n_406),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_429),
.A2(n_426),
.B(n_430),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_430),
.A2(n_440),
.B1(n_404),
.B2(n_410),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_396),
.C(n_379),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_439),
.C(n_442),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_392),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_432),
.B(n_435),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_441),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_401),
.C(n_398),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_399),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_394),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_433),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_447),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_425),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_445),
.B(n_451),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_439),
.B(n_412),
.C(n_414),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_427),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_452),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_450),
.A2(n_438),
.B1(n_418),
.B2(n_437),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_434),
.A2(n_405),
.B(n_415),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_453),
.B(n_442),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_405),
.C(n_407),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_454),
.B(n_455),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_436),
.A2(n_409),
.B(n_417),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_458),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_431),
.C(n_433),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_460),
.B(n_463),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_322),
.C(n_334),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_464),
.B(n_447),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_466),
.B(n_469),
.C(n_463),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_459),
.A2(n_452),
.B(n_454),
.Y(n_468)
);

AO221x1_ASAP7_75t_L g474 ( 
.A1(n_468),
.A2(n_470),
.B1(n_465),
.B2(n_457),
.C(n_448),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_455),
.C(n_448),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_462),
.A2(n_453),
.B(n_456),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_467),
.B(n_461),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_472),
.B(n_473),
.C(n_475),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_474),
.A2(n_471),
.B(n_385),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_385),
.C(n_334),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_477),
.A2(n_319),
.B(n_359),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_478),
.A2(n_479),
.B(n_330),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g479 ( 
.A(n_476),
.B(n_283),
.C(n_359),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_480),
.A2(n_330),
.B(n_283),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_330),
.Y(n_482)
);


endmodule