module fake_jpeg_31406_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_2),
.B(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_14),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_54),
.Y(n_103)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_20),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_47),
.Y(n_117)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_13),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_79),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_13),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_57),
.B(n_60),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_62),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_70),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_17),
.B(n_0),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_27),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_74),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_35),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_78),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_1),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_34),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_82),
.Y(n_115)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_85),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_86),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_48),
.B(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_44),
.A2(n_45),
.B1(n_77),
.B2(n_75),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_97),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_26),
.B1(n_43),
.B2(n_32),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_136),
.B1(n_69),
.B2(n_55),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_21),
.B1(n_42),
.B2(n_29),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_105),
.A2(n_118),
.B1(n_8),
.B2(n_10),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_59),
.A2(n_24),
.B1(n_40),
.B2(n_34),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_130),
.B1(n_37),
.B2(n_18),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_43),
.B1(n_32),
.B2(n_39),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_43),
.B1(n_32),
.B2(n_39),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_66),
.A2(n_42),
.B1(n_21),
.B2(n_29),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_74),
.A2(n_32),
.B1(n_39),
.B2(n_38),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_119),
.A2(n_135),
.B1(n_114),
.B2(n_97),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_31),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_131),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_48),
.A2(n_16),
.B(n_31),
.C(n_33),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_21),
.B(n_66),
.C(n_54),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_80),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_63),
.B(n_16),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_67),
.A2(n_38),
.B1(n_37),
.B2(n_42),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_49),
.A2(n_26),
.B1(n_37),
.B2(n_29),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_138),
.B(n_142),
.Y(n_205)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_140),
.A2(n_153),
.B1(n_162),
.B2(n_173),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_141),
.A2(n_174),
.B1(n_162),
.B2(n_168),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_98),
.A2(n_54),
.B(n_35),
.C(n_83),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_35),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_175),
.Y(n_192)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_145),
.Y(n_222)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

BUFx2_ASAP7_75t_SL g148 ( 
.A(n_89),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_91),
.A2(n_50),
.B1(n_52),
.B2(n_82),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_152),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_52),
.B1(n_35),
.B2(n_5),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_155),
.A2(n_177),
.B1(n_178),
.B2(n_180),
.Y(n_217)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_156),
.Y(n_189)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_90),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_159),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_111),
.B(n_6),
.Y(n_159)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_100),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_6),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_165),
.Y(n_196)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_6),
.Y(n_165)
);

CKINVDCx12_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_168),
.Y(n_202)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_118),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_170),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_101),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_115),
.B(n_7),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_179),
.Y(n_214)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_172),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_104),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_119),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_136),
.A2(n_11),
.B1(n_95),
.B2(n_108),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_96),
.A2(n_11),
.B1(n_108),
.B2(n_134),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_103),
.B(n_11),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_182),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_103),
.B(n_105),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_183),
.A2(n_124),
.B1(n_102),
.B2(n_99),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_124),
.B1(n_118),
.B2(n_133),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_185),
.A2(n_206),
.B1(n_199),
.B2(n_208),
.Y(n_245)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_123),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_207),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_219),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_211),
.B1(n_146),
.B2(n_161),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_144),
.A2(n_110),
.B(n_89),
.C(n_88),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_181),
.B(n_149),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_102),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_208),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_140),
.A2(n_133),
.B1(n_125),
.B2(n_121),
.Y(n_206)
);

AOI32xp33_ASAP7_75t_L g207 ( 
.A1(n_160),
.A2(n_101),
.A3(n_125),
.B1(n_121),
.B2(n_94),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_110),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_183),
.A2(n_94),
.B1(n_174),
.B2(n_176),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_176),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_156),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_152),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_137),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_142),
.B(n_153),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_224),
.A2(n_220),
.B1(n_217),
.B2(n_200),
.Y(n_260)
);

NOR2x1_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_173),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_226),
.A2(n_237),
.B(n_241),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_228),
.A2(n_227),
.B1(n_241),
.B2(n_248),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_231),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_238),
.B(n_242),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_170),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_143),
.B1(n_180),
.B2(n_147),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_245),
.B1(n_250),
.B2(n_253),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_150),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_256),
.C(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_202),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_254),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_167),
.B(n_145),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_157),
.B(n_164),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_192),
.A2(n_143),
.B(n_147),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_204),
.A2(n_154),
.B(n_180),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_154),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_230),
.B(n_242),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_195),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_246),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_218),
.B(n_184),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_219),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_249),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_197),
.A2(n_211),
.B1(n_219),
.B2(n_224),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_184),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_197),
.A2(n_206),
.B1(n_216),
.B2(n_198),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_214),
.B(n_215),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_257),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_196),
.B(n_197),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_207),
.B(n_194),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_223),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_189),
.B(n_194),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_259),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_220),
.B1(n_222),
.B2(n_210),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_243),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_222),
.B1(n_213),
.B2(n_212),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_266),
.A2(n_273),
.B1(n_288),
.B2(n_257),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_231),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_269),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_212),
.B1(n_193),
.B2(n_186),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_210),
.A3(n_193),
.B1(n_223),
.B2(n_189),
.C1(n_186),
.C2(n_209),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_276),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_277),
.B(n_285),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_209),
.C(n_234),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_287),
.C(n_285),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_228),
.A2(n_260),
.B1(n_227),
.B2(n_232),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_235),
.B1(n_239),
.B2(n_249),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_291),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_286),
.B(n_243),
.Y(n_298)
);

XOR2x1_ASAP7_75t_L g286 ( 
.A(n_225),
.B(n_237),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_225),
.B(n_256),
.C(n_246),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_233),
.B1(n_226),
.B2(n_238),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_244),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_229),
.B(n_226),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_290),
.B(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_294),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_269),
.B(n_272),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_295),
.A2(n_286),
.B1(n_276),
.B2(n_289),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_296),
.A2(n_301),
.B1(n_316),
.B2(n_279),
.Y(n_326)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_298),
.B(n_307),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_303),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_254),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_252),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_305),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_282),
.B(n_272),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_291),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_306),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_287),
.C(n_278),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_312),
.C(n_275),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_282),
.B(n_283),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_313),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_277),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_275),
.B(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_268),
.Y(n_314)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_280),
.B1(n_289),
.B2(n_274),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_261),
.A2(n_288),
.B1(n_273),
.B2(n_281),
.Y(n_316)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_309),
.Y(n_318)
);

INVx13_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_319),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_299),
.A2(n_261),
.B1(n_311),
.B2(n_281),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_325),
.A2(n_293),
.B1(n_313),
.B2(n_305),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_326),
.A2(n_331),
.B1(n_338),
.B2(n_315),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_332),
.C(n_336),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_267),
.B1(n_266),
.B2(n_270),
.Y(n_330)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_301),
.A2(n_265),
.B1(n_270),
.B2(n_284),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_286),
.C(n_280),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_295),
.B(n_331),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_267),
.C(n_271),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_296),
.A2(n_271),
.B1(n_316),
.B2(n_295),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_317),
.C(n_298),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_322),
.C(n_329),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_340),
.A2(n_346),
.B(n_326),
.Y(n_359)
);

OAI22x1_ASAP7_75t_L g341 ( 
.A1(n_335),
.A2(n_293),
.B1(n_294),
.B2(n_299),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_341),
.A2(n_343),
.B1(n_348),
.B2(n_356),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_338),
.A2(n_317),
.B(n_302),
.Y(n_345)
);

AOI21x1_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_357),
.B(n_340),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_327),
.A2(n_319),
.B(n_325),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_321),
.A2(n_310),
.B1(n_297),
.B2(n_314),
.Y(n_348)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_349),
.Y(n_360)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_351),
.Y(n_371)
);

FAx1_ASAP7_75t_SL g352 ( 
.A(n_321),
.B(n_322),
.CI(n_332),
.CON(n_352),
.SN(n_352)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_357),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_344),
.Y(n_358)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_354),
.Y(n_364)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_333),
.Y(n_355)
);

INVx11_ASAP7_75t_L g363 ( 
.A(n_355),
.Y(n_363)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_362),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_359),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_346),
.A2(n_339),
.B(n_319),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_336),
.C(n_337),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_368),
.C(n_352),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_334),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_366),
.B(n_345),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_323),
.C(n_324),
.Y(n_368)
);

NAND4xp25_ASAP7_75t_SL g369 ( 
.A(n_341),
.B(n_350),
.C(n_343),
.D(n_347),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_369),
.B(n_346),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_350),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_375),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_361),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_342),
.C(n_349),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_358),
.C(n_366),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_363),
.B(n_355),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_380),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_369),
.A2(n_342),
.B1(n_354),
.B2(n_351),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_379),
.A2(n_360),
.B1(n_371),
.B2(n_370),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_359),
.A2(n_348),
.B1(n_346),
.B2(n_356),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_368),
.A2(n_350),
.B(n_347),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_367),
.B(n_371),
.Y(n_387)
);

XOR2x1_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_362),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_385),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_391),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_373),
.A2(n_361),
.B1(n_360),
.B2(n_367),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_390),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_389),
.B(n_377),
.C(n_374),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_364),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_392),
.B(n_394),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_377),
.Y(n_394)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_386),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_396),
.A2(n_373),
.B1(n_384),
.B2(n_382),
.Y(n_401)
);

OAI221xp5_ASAP7_75t_L g398 ( 
.A1(n_393),
.A2(n_385),
.B1(n_364),
.B2(n_363),
.C(n_383),
.Y(n_398)
);

AOI21xp33_ASAP7_75t_L g403 ( 
.A1(n_398),
.A2(n_396),
.B(n_397),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_395),
.A2(n_388),
.B(n_375),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_401),
.C(n_395),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_402),
.B(n_400),
.C(n_350),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_403),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_347),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_405),
.Y(n_407)
);


endmodule