module fake_jpeg_8737_n_32 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_32);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_32;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_15;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_6),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_7),
.B1(n_9),
.B2(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_12),
.A2(n_1),
.B(n_16),
.Y(n_23)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_19),
.A3(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_24)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_26),
.B1(n_21),
.B2(n_17),
.Y(n_28)
);

MAJx2_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_26),
.C(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_30),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_15),
.B(n_20),
.C(n_29),
.Y(n_32)
);


endmodule