module real_aes_7213_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g463 ( .A1(n_0), .A2(n_164), .B(n_464), .C(n_467), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_1), .B(n_458), .Y(n_469) );
INVx1_ASAP7_75t_L g427 ( .A(n_2), .Y(n_427) );
INVx1_ASAP7_75t_L g213 ( .A(n_3), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_4), .B(n_152), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_5), .A2(n_104), .B1(n_737), .B2(n_746), .C1(n_761), .C2(n_767), .Y(n_103) );
OAI211xp5_ASAP7_75t_L g746 ( .A1(n_5), .A2(n_747), .B(n_757), .C(n_760), .Y(n_746) );
OAI211xp5_ASAP7_75t_L g757 ( .A1(n_5), .A2(n_749), .B(n_754), .C(n_758), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_6), .A2(n_442), .B(n_512), .Y(n_511) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_7), .A2(n_10), .B1(n_422), .B2(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_7), .Y(n_753) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_8), .A2(n_169), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_9), .A2(n_38), .B1(n_125), .B2(n_137), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g108 ( .A1(n_10), .A2(n_109), .B1(n_110), .B2(n_422), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_10), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_11), .B(n_169), .Y(n_202) );
AND2x6_ASAP7_75t_L g140 ( .A(n_12), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_13), .A2(n_140), .B(n_445), .C(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_14), .B(n_39), .Y(n_428) );
INVx1_ASAP7_75t_L g121 ( .A(n_15), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_16), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g207 ( .A(n_17), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_18), .B(n_152), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_19), .B(n_167), .Y(n_185) );
AO32x2_ASAP7_75t_L g161 ( .A1(n_20), .A2(n_162), .A3(n_166), .B1(n_168), .B2(n_169), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_21), .A2(n_57), .B1(n_729), .B2(n_730), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_21), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_22), .B(n_125), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_23), .B(n_167), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_24), .A2(n_55), .B1(n_125), .B2(n_137), .Y(n_165) );
AOI22xp33_ASAP7_75t_SL g178 ( .A1(n_25), .A2(n_82), .B1(n_125), .B2(n_129), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_26), .B(n_125), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_27), .A2(n_168), .B(n_445), .C(n_447), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_28), .A2(n_168), .B(n_445), .C(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_29), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_30), .B(n_117), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_31), .A2(n_442), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_32), .B(n_117), .Y(n_159) );
INVx2_ASAP7_75t_L g127 ( .A(n_33), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_34), .A2(n_476), .B(n_477), .C(n_481), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_35), .B(n_125), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_36), .B(n_117), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_37), .B(n_132), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_40), .B(n_441), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_41), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_42), .B(n_152), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_43), .B(n_442), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_44), .A2(n_476), .B(n_481), .C(n_503), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_45), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_45), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_46), .B(n_125), .Y(n_195) );
INVx1_ASAP7_75t_L g465 ( .A(n_47), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_48), .A2(n_91), .B1(n_137), .B2(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g504 ( .A(n_49), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_50), .B(n_125), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_51), .B(n_125), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_52), .B(n_744), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_53), .B(n_442), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_54), .B(n_200), .Y(n_199) );
AOI22xp33_ASAP7_75t_SL g189 ( .A1(n_56), .A2(n_61), .B1(n_125), .B2(n_129), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_57), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_58), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_59), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_60), .B(n_125), .Y(n_226) );
INVx1_ASAP7_75t_L g141 ( .A(n_62), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_63), .B(n_442), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_64), .B(n_458), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_65), .A2(n_200), .B(n_210), .C(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_66), .B(n_125), .Y(n_214) );
INVx1_ASAP7_75t_L g120 ( .A(n_67), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_68), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_69), .B(n_152), .Y(n_479) );
AO32x2_ASAP7_75t_L g174 ( .A1(n_70), .A2(n_168), .A3(n_169), .B1(n_175), .B2(n_179), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_71), .B(n_153), .Y(n_535) );
INVx1_ASAP7_75t_L g225 ( .A(n_72), .Y(n_225) );
INVx1_ASAP7_75t_L g150 ( .A(n_73), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_74), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_75), .B(n_449), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_76), .A2(n_445), .B(n_481), .C(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_77), .B(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_77), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_78), .B(n_129), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_79), .Y(n_513) );
INVx1_ASAP7_75t_L g741 ( .A(n_80), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_81), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_83), .B(n_137), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_84), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_85), .B(n_129), .Y(n_156) );
AOI222xp33_ASAP7_75t_L g105 ( .A1(n_86), .A2(n_106), .B1(n_724), .B2(n_725), .C1(n_731), .C2(n_733), .Y(n_105) );
INVx2_ASAP7_75t_L g118 ( .A(n_87), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_88), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_89), .B(n_139), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_90), .B(n_129), .Y(n_196) );
OR2x2_ASAP7_75t_L g425 ( .A(n_92), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g723 ( .A(n_92), .Y(n_723) );
OR2x2_ASAP7_75t_L g745 ( .A(n_92), .B(n_736), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_93), .A2(n_102), .B1(n_129), .B2(n_130), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_94), .B(n_442), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_95), .Y(n_478) );
INVxp67_ASAP7_75t_L g516 ( .A(n_96), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_97), .B(n_129), .Y(n_223) );
INVx1_ASAP7_75t_L g491 ( .A(n_98), .Y(n_491) );
INVx1_ASAP7_75t_L g531 ( .A(n_99), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_100), .B(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g506 ( .A(n_101), .B(n_117), .Y(n_506) );
INVxp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22x1_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_423), .B1(n_429), .B2(n_720), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_108), .A2(n_430), .B1(n_720), .B2(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_109), .A2(n_110), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_344), .Y(n_110) );
NAND5xp2_ASAP7_75t_L g111 ( .A(n_112), .B(n_263), .C(n_278), .D(n_304), .E(n_326), .Y(n_111) );
NOR2xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_243), .Y(n_112) );
OAI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_180), .B1(n_216), .B2(n_232), .C(n_233), .Y(n_113) );
NOR2xp33_ASAP7_75t_SL g114 ( .A(n_115), .B(n_170), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_115), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_SL g420 ( .A(n_115), .Y(n_420) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_143), .Y(n_115) );
INVx1_ASAP7_75t_L g260 ( .A(n_116), .Y(n_260) );
AND2x2_ASAP7_75t_L g262 ( .A(n_116), .B(n_161), .Y(n_262) );
AND2x2_ASAP7_75t_L g272 ( .A(n_116), .B(n_160), .Y(n_272) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_116), .Y(n_290) );
INVx1_ASAP7_75t_L g300 ( .A(n_116), .Y(n_300) );
OR2x2_ASAP7_75t_L g338 ( .A(n_116), .B(n_237), .Y(n_338) );
INVx2_ASAP7_75t_L g388 ( .A(n_116), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_116), .B(n_236), .Y(n_405) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_142), .Y(n_116) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_117), .A2(n_147), .B(n_159), .Y(n_146) );
INVx2_ASAP7_75t_L g179 ( .A(n_117), .Y(n_179) );
INVx1_ASAP7_75t_L g455 ( .A(n_117), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_117), .A2(n_474), .B(n_475), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_117), .A2(n_501), .B(n_502), .Y(n_500) );
AND2x2_ASAP7_75t_SL g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AND2x2_ASAP7_75t_L g167 ( .A(n_118), .B(n_119), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_134), .B(n_140), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_128), .B(n_131), .Y(n_123) );
INVx3_ASAP7_75t_L g149 ( .A(n_125), .Y(n_149) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_125), .Y(n_493) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g137 ( .A(n_126), .Y(n_137) );
BUFx3_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
AND2x6_ASAP7_75t_L g445 ( .A(n_126), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g130 ( .A(n_127), .Y(n_130) );
INVx1_ASAP7_75t_L g201 ( .A(n_127), .Y(n_201) );
INVx2_ASAP7_75t_L g208 ( .A(n_129), .Y(n_208) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx3_ASAP7_75t_L g153 ( .A(n_133), .Y(n_153) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_133), .Y(n_158) );
AND2x2_ASAP7_75t_L g443 ( .A(n_133), .B(n_201), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_133), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_138), .Y(n_134) );
O2A1O1Ixp5_ASAP7_75t_L g224 ( .A1(n_138), .A2(n_212), .B(n_225), .C(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_139), .A2(n_163), .B1(n_164), .B2(n_165), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g175 ( .A1(n_139), .A2(n_153), .B1(n_176), .B2(n_178), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_139), .A2(n_164), .B1(n_188), .B2(n_189), .Y(n_187) );
INVx4_ASAP7_75t_L g466 ( .A(n_139), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g147 ( .A1(n_140), .A2(n_148), .B(n_154), .Y(n_147) );
BUFx3_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_140), .A2(n_194), .B(n_197), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_140), .A2(n_206), .B(n_211), .Y(n_205) );
AND2x4_ASAP7_75t_L g442 ( .A(n_140), .B(n_443), .Y(n_442) );
INVx4_ASAP7_75t_SL g468 ( .A(n_140), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_140), .B(n_443), .Y(n_532) );
NOR2xp67_ASAP7_75t_L g143 ( .A(n_144), .B(n_160), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_145), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_145), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_SL g320 ( .A(n_145), .B(n_260), .Y(n_320) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
INVx2_ASAP7_75t_L g237 ( .A(n_146), .Y(n_237) );
OR2x2_ASAP7_75t_L g299 ( .A(n_146), .B(n_300), .Y(n_299) );
O2A1O1Ixp5_ASAP7_75t_SL g148 ( .A1(n_149), .A2(n_150), .B(n_151), .C(n_152), .Y(n_148) );
INVx2_ASAP7_75t_L g164 ( .A(n_152), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_152), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_152), .A2(n_222), .B(n_223), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_152), .B(n_516), .Y(n_515) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_157), .Y(n_154) );
INVx1_ASAP7_75t_L g210 ( .A(n_157), .Y(n_210) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g449 ( .A(n_158), .Y(n_449) );
AND2x2_ASAP7_75t_L g238 ( .A(n_160), .B(n_174), .Y(n_238) );
AND2x2_ASAP7_75t_L g255 ( .A(n_160), .B(n_235), .Y(n_255) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g173 ( .A(n_161), .B(n_174), .Y(n_173) );
BUFx2_ASAP7_75t_L g258 ( .A(n_161), .Y(n_258) );
AND2x2_ASAP7_75t_L g387 ( .A(n_161), .B(n_388), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_164), .A2(n_198), .B(n_199), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_164), .A2(n_212), .B(n_213), .C(n_214), .Y(n_211) );
INVx2_ASAP7_75t_L g204 ( .A(n_166), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_166), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_167), .Y(n_169) );
NAND3xp33_ASAP7_75t_L g186 ( .A(n_168), .B(n_187), .C(n_190), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_168), .A2(n_221), .B(n_224), .Y(n_220) );
INVx4_ASAP7_75t_L g190 ( .A(n_169), .Y(n_190) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_169), .A2(n_193), .B(n_202), .Y(n_192) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_169), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_169), .A2(n_522), .B(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g232 ( .A(n_170), .Y(n_232) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_173), .Y(n_170) );
AND2x2_ASAP7_75t_L g350 ( .A(n_171), .B(n_238), .Y(n_350) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g351 ( .A(n_172), .B(n_262), .Y(n_351) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_173), .A2(n_319), .B(n_321), .C(n_323), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_173), .B(n_319), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_173), .A2(n_249), .B1(n_392), .B2(n_393), .C(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g235 ( .A(n_174), .Y(n_235) );
INVx1_ASAP7_75t_L g271 ( .A(n_174), .Y(n_271) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_174), .Y(n_280) );
INVx2_ASAP7_75t_L g467 ( .A(n_177), .Y(n_467) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_177), .Y(n_480) );
INVx1_ASAP7_75t_L g452 ( .A(n_179), .Y(n_452) );
INVx1_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_191), .Y(n_181) );
AND2x2_ASAP7_75t_L g297 ( .A(n_182), .B(n_242), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_182), .B(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_183), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g389 ( .A(n_183), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g421 ( .A(n_183), .Y(n_421) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx3_ASAP7_75t_L g251 ( .A(n_184), .Y(n_251) );
AND2x2_ASAP7_75t_L g277 ( .A(n_184), .B(n_231), .Y(n_277) );
NOR2x1_ASAP7_75t_L g286 ( .A(n_184), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g293 ( .A(n_184), .B(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
INVx1_ASAP7_75t_L g229 ( .A(n_185), .Y(n_229) );
AO21x1_ASAP7_75t_L g228 ( .A1(n_187), .A2(n_190), .B(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g458 ( .A(n_190), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_190), .B(n_483), .Y(n_482) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_190), .A2(n_488), .B(n_495), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_190), .B(n_496), .Y(n_495) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_190), .A2(n_530), .B(n_537), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_191), .B(n_333), .Y(n_368) );
INVx1_ASAP7_75t_SL g372 ( .A(n_191), .Y(n_372) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_203), .Y(n_191) );
INVx3_ASAP7_75t_L g231 ( .A(n_192), .Y(n_231) );
AND2x2_ASAP7_75t_L g242 ( .A(n_192), .B(n_219), .Y(n_242) );
AND2x2_ASAP7_75t_L g264 ( .A(n_192), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g309 ( .A(n_192), .B(n_303), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_192), .B(n_241), .Y(n_390) );
INVx2_ASAP7_75t_L g212 ( .A(n_200), .Y(n_212) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g230 ( .A(n_203), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g241 ( .A(n_203), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_203), .B(n_219), .Y(n_266) );
AND2x2_ASAP7_75t_L g302 ( .A(n_203), .B(n_303), .Y(n_302) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_215), .Y(n_203) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_204), .A2(n_220), .B(n_227), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_209), .C(n_210), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_208), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_208), .A2(n_535), .B(n_536), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_210), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_212), .A2(n_448), .B(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_230), .Y(n_217) );
INVx1_ASAP7_75t_L g282 ( .A(n_218), .Y(n_282) );
AND2x2_ASAP7_75t_L g324 ( .A(n_218), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_218), .B(n_245), .Y(n_330) );
AOI21xp5_ASAP7_75t_SL g404 ( .A1(n_218), .A2(n_236), .B(n_259), .Y(n_404) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_228), .Y(n_218) );
OR2x2_ASAP7_75t_L g247 ( .A(n_219), .B(n_228), .Y(n_247) );
AND2x2_ASAP7_75t_L g294 ( .A(n_219), .B(n_231), .Y(n_294) );
INVx2_ASAP7_75t_L g303 ( .A(n_219), .Y(n_303) );
INVx1_ASAP7_75t_L g409 ( .A(n_219), .Y(n_409) );
AND2x2_ASAP7_75t_L g333 ( .A(n_228), .B(n_303), .Y(n_333) );
INVx1_ASAP7_75t_L g358 ( .A(n_228), .Y(n_358) );
AND2x2_ASAP7_75t_L g267 ( .A(n_230), .B(n_251), .Y(n_267) );
AND2x2_ASAP7_75t_L g279 ( .A(n_230), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_SL g397 ( .A(n_230), .Y(n_397) );
INVx2_ASAP7_75t_L g287 ( .A(n_231), .Y(n_287) );
AND2x2_ASAP7_75t_L g325 ( .A(n_231), .B(n_241), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_231), .B(n_409), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_238), .B(n_239), .Y(n_233) );
AND2x2_ASAP7_75t_L g340 ( .A(n_234), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g394 ( .A(n_234), .Y(n_394) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
INVx1_ASAP7_75t_L g314 ( .A(n_235), .Y(n_314) );
BUFx2_ASAP7_75t_L g413 ( .A(n_235), .Y(n_413) );
BUFx2_ASAP7_75t_L g284 ( .A(n_236), .Y(n_284) );
AND2x2_ASAP7_75t_L g386 ( .A(n_236), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g369 ( .A(n_237), .Y(n_369) );
AND2x4_ASAP7_75t_L g296 ( .A(n_238), .B(n_259), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_238), .B(n_320), .Y(n_332) );
AOI32xp33_ASAP7_75t_L g256 ( .A1(n_239), .A2(n_257), .A3(n_259), .B1(n_261), .B2(n_262), .Y(n_256) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
INVx3_ASAP7_75t_L g245 ( .A(n_240), .Y(n_245) );
OR2x2_ASAP7_75t_L g381 ( .A(n_240), .B(n_337), .Y(n_381) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g250 ( .A(n_241), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g357 ( .A(n_241), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g249 ( .A(n_242), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g261 ( .A(n_242), .B(n_251), .Y(n_261) );
INVx1_ASAP7_75t_L g382 ( .A(n_242), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_242), .B(n_357), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_248), .B(n_252), .C(n_256), .Y(n_243) );
OAI322xp33_ASAP7_75t_L g352 ( .A1(n_244), .A2(n_289), .A3(n_353), .B1(n_355), .B2(n_359), .C1(n_360), .C2(n_364), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVxp67_ASAP7_75t_L g317 ( .A(n_245), .Y(n_317) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g371 ( .A(n_247), .B(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_247), .B(n_287), .Y(n_418) );
INVxp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g310 ( .A(n_250), .Y(n_310) );
OR2x2_ASAP7_75t_L g396 ( .A(n_251), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_254), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g305 ( .A(n_255), .B(n_284), .Y(n_305) );
AND2x2_ASAP7_75t_L g376 ( .A(n_255), .B(n_289), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_255), .B(n_363), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_257), .A2(n_264), .B1(n_267), .B2(n_268), .C(n_273), .Y(n_263) );
OR2x2_ASAP7_75t_L g274 ( .A(n_257), .B(n_270), .Y(n_274) );
AND2x2_ASAP7_75t_L g362 ( .A(n_257), .B(n_363), .Y(n_362) );
AOI32xp33_ASAP7_75t_L g401 ( .A1(n_257), .A2(n_287), .A3(n_402), .B1(n_403), .B2(n_406), .Y(n_401) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_258), .B(n_294), .C(n_317), .Y(n_335) );
AND2x2_ASAP7_75t_L g361 ( .A(n_258), .B(n_354), .Y(n_361) );
INVxp67_ASAP7_75t_L g341 ( .A(n_259), .Y(n_341) );
BUFx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_262), .B(n_314), .Y(n_370) );
INVx2_ASAP7_75t_L g380 ( .A(n_262), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_262), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g349 ( .A(n_265), .Y(n_349) );
OR2x2_ASAP7_75t_L g275 ( .A(n_266), .B(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_268), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_271), .Y(n_354) );
AND2x2_ASAP7_75t_L g313 ( .A(n_272), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g359 ( .A(n_272), .Y(n_359) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_272), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AOI21xp33_ASAP7_75t_SL g298 ( .A1(n_274), .A2(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g392 ( .A(n_277), .B(n_302), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_281), .B(n_291), .C(n_298), .Y(n_278) );
AND2x2_ASAP7_75t_L g322 ( .A(n_280), .B(n_290), .Y(n_322) );
INVx2_ASAP7_75t_L g337 ( .A(n_280), .Y(n_337) );
OR2x2_ASAP7_75t_L g375 ( .A(n_280), .B(n_338), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_280), .B(n_418), .Y(n_417) );
AOI211xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_283), .B(n_285), .C(n_288), .Y(n_281) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_284), .B(n_322), .Y(n_321) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_285), .A2(n_380), .B(n_404), .C(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_286), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g343 ( .A(n_287), .B(n_333), .Y(n_343) );
INVx1_ASAP7_75t_L g348 ( .A(n_287), .Y(n_348) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVxp33_ASAP7_75t_L g399 ( .A(n_293), .Y(n_399) );
AND2x2_ASAP7_75t_L g378 ( .A(n_294), .B(n_357), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_299), .A2(n_361), .B(n_362), .Y(n_360) );
OAI322xp33_ASAP7_75t_L g379 ( .A1(n_301), .A2(n_380), .A3(n_381), .B1(n_382), .B2(n_383), .C1(n_385), .C2(n_389), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_311), .B2(n_315), .C(n_318), .Y(n_304) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g356 ( .A(n_309), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g400 ( .A(n_313), .Y(n_400) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_316), .B(n_336), .Y(n_402) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g365 ( .A(n_325), .B(n_333), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B1(n_331), .B2(n_333), .C(n_334), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_329), .A2(n_346), .B1(n_350), .B2(n_351), .C(n_352), .Y(n_345) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVxp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_333), .B(n_348), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_339), .B2(n_342), .Y(n_334) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx2_ASAP7_75t_SL g363 ( .A(n_338), .Y(n_363) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND5xp2_ASAP7_75t_L g344 ( .A(n_345), .B(n_366), .C(n_391), .D(n_401), .E(n_411), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_347), .B(n_349), .Y(n_346) );
NOR4xp25_ASAP7_75t_L g419 ( .A(n_348), .B(n_354), .C(n_420), .D(n_421), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_351), .A2(n_412), .B1(n_414), .B2(n_416), .C(n_419), .Y(n_411) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g410 ( .A(n_357), .Y(n_410) );
OAI322xp33_ASAP7_75t_L g367 ( .A1(n_361), .A2(n_368), .A3(n_369), .B1(n_370), .B2(n_371), .C1(n_373), .C2(n_377), .Y(n_367) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_367), .B(n_379), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g412 ( .A(n_387), .B(n_413), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B1(n_399), .B2(n_400), .Y(n_395) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g732 ( .A(n_424), .Y(n_732) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g722 ( .A(n_426), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g736 ( .A(n_426), .Y(n_736) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_431), .B(n_675), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_610), .Y(n_431) );
NAND4xp25_ASAP7_75t_SL g432 ( .A(n_433), .B(n_555), .C(n_579), .D(n_602), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_497), .B1(n_527), .B2(n_539), .C(n_542), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_470), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_436), .A2(n_456), .B1(n_498), .B2(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_436), .B(n_471), .Y(n_613) );
AND2x2_ASAP7_75t_L g632 ( .A(n_436), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_436), .B(n_616), .Y(n_702) );
AND2x4_ASAP7_75t_L g436 ( .A(n_437), .B(n_456), .Y(n_436) );
AND2x2_ASAP7_75t_L g570 ( .A(n_437), .B(n_471), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_437), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g593 ( .A(n_437), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g598 ( .A(n_437), .B(n_457), .Y(n_598) );
INVx2_ASAP7_75t_L g630 ( .A(n_437), .Y(n_630) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_437), .Y(n_674) );
AND2x2_ASAP7_75t_L g691 ( .A(n_437), .B(n_568), .Y(n_691) );
INVx5_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g609 ( .A(n_438), .B(n_568), .Y(n_609) );
AND2x4_ASAP7_75t_L g623 ( .A(n_438), .B(n_456), .Y(n_623) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_438), .Y(n_627) );
AND2x2_ASAP7_75t_L g647 ( .A(n_438), .B(n_562), .Y(n_647) );
AND2x2_ASAP7_75t_L g697 ( .A(n_438), .B(n_472), .Y(n_697) );
AND2x2_ASAP7_75t_L g707 ( .A(n_438), .B(n_457), .Y(n_707) );
OR2x6_ASAP7_75t_L g438 ( .A(n_439), .B(n_453), .Y(n_438) );
AOI21xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_444), .B(n_452), .Y(n_439) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx5_ASAP7_75t_L g462 ( .A(n_445), .Y(n_462) );
INVx2_ASAP7_75t_L g451 ( .A(n_449), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_451), .A2(n_478), .B(n_479), .C(n_480), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_451), .A2(n_480), .B(n_504), .C(n_505), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x2_ASAP7_75t_L g563 ( .A(n_456), .B(n_471), .Y(n_563) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_456), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_456), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g653 ( .A(n_456), .Y(n_653) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g541 ( .A(n_457), .B(n_486), .Y(n_541) );
AND2x2_ASAP7_75t_L g568 ( .A(n_457), .B(n_487), .Y(n_568) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_469), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_462), .B(n_463), .C(n_468), .Y(n_460) );
INVx2_ASAP7_75t_L g476 ( .A(n_462), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_462), .A2(n_468), .B(n_513), .C(n_514), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g481 ( .A(n_468), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_470), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_484), .Y(n_470) );
OR2x2_ASAP7_75t_L g594 ( .A(n_471), .B(n_485), .Y(n_594) );
AND2x2_ASAP7_75t_L g631 ( .A(n_471), .B(n_541), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_471), .B(n_562), .Y(n_642) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_471), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_471), .B(n_598), .Y(n_715) );
INVx5_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g540 ( .A(n_472), .Y(n_540) );
AND2x2_ASAP7_75t_L g549 ( .A(n_472), .B(n_485), .Y(n_549) );
AND2x2_ASAP7_75t_L g665 ( .A(n_472), .B(n_560), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_472), .B(n_598), .Y(n_687) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_482), .Y(n_472) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_485), .Y(n_633) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_486), .Y(n_585) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g562 ( .A(n_487), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_494), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_498), .B(n_575), .Y(n_694) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_499), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g546 ( .A(n_499), .B(n_547), .Y(n_546) );
INVx5_ASAP7_75t_SL g554 ( .A(n_499), .Y(n_554) );
OR2x2_ASAP7_75t_L g577 ( .A(n_499), .B(n_547), .Y(n_577) );
OR2x2_ASAP7_75t_L g587 ( .A(n_499), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g650 ( .A(n_499), .B(n_509), .Y(n_650) );
AND2x2_ASAP7_75t_SL g688 ( .A(n_499), .B(n_508), .Y(n_688) );
NOR4xp25_ASAP7_75t_L g709 ( .A(n_499), .B(n_630), .C(n_710), .D(n_711), .Y(n_709) );
AND2x2_ASAP7_75t_L g719 ( .A(n_499), .B(n_551), .Y(n_719) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .Y(n_499) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g544 ( .A(n_508), .B(n_540), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_508), .B(n_546), .Y(n_713) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_518), .Y(n_508) );
OR2x2_ASAP7_75t_L g553 ( .A(n_509), .B(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g560 ( .A(n_509), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_509), .B(n_529), .Y(n_572) );
INVxp67_ASAP7_75t_L g575 ( .A(n_509), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_509), .B(n_547), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_509), .B(n_519), .Y(n_641) );
AND2x2_ASAP7_75t_L g656 ( .A(n_509), .B(n_551), .Y(n_656) );
OR2x2_ASAP7_75t_L g685 ( .A(n_509), .B(n_519), .Y(n_685) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_517), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_518), .B(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_518), .B(n_554), .Y(n_693) );
OR2x2_ASAP7_75t_L g714 ( .A(n_518), .B(n_591), .Y(n_714) );
INVx1_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g528 ( .A(n_519), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g551 ( .A(n_519), .B(n_547), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_519), .B(n_529), .Y(n_566) );
AND2x2_ASAP7_75t_L g636 ( .A(n_519), .B(n_560), .Y(n_636) );
AND2x2_ASAP7_75t_L g670 ( .A(n_519), .B(n_554), .Y(n_670) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_520), .B(n_554), .Y(n_573) );
AND2x2_ASAP7_75t_L g601 ( .A(n_520), .B(n_529), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_527), .B(n_609), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_528), .A2(n_616), .B1(n_652), .B2(n_669), .C(n_671), .Y(n_668) );
INVx5_ASAP7_75t_SL g547 ( .A(n_529), .Y(n_547) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
OAI33xp33_ASAP7_75t_L g567 ( .A1(n_540), .A2(n_568), .A3(n_569), .B1(n_571), .B2(n_574), .B3(n_578), .Y(n_567) );
OR2x2_ASAP7_75t_L g583 ( .A(n_540), .B(n_584), .Y(n_583) );
AOI322xp5_ASAP7_75t_L g692 ( .A1(n_540), .A2(n_609), .A3(n_616), .B1(n_693), .B2(n_694), .C1(n_695), .C2(n_698), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_540), .B(n_568), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_SL g716 ( .A1(n_540), .A2(n_568), .B(n_717), .C(n_719), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_541), .A2(n_556), .B1(n_561), .B2(n_564), .C(n_567), .Y(n_555) );
INVx1_ASAP7_75t_L g648 ( .A(n_541), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_541), .B(n_697), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_545), .B1(n_548), .B2(n_550), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g625 ( .A(n_546), .B(n_560), .Y(n_625) );
AND2x2_ASAP7_75t_L g683 ( .A(n_546), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g591 ( .A(n_547), .B(n_554), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_547), .B(n_560), .Y(n_619) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_549), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_549), .B(n_627), .Y(n_681) );
OAI321xp33_ASAP7_75t_L g700 ( .A1(n_549), .A2(n_622), .A3(n_701), .B1(n_702), .B2(n_703), .C(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g667 ( .A(n_550), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_551), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g606 ( .A(n_551), .B(n_554), .Y(n_606) );
AOI321xp33_ASAP7_75t_L g664 ( .A1(n_551), .A2(n_568), .A3(n_665), .B1(n_666), .B2(n_667), .C(n_668), .Y(n_664) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g581 ( .A(n_553), .B(n_566), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_554), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_554), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_554), .B(n_640), .Y(n_677) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g600 ( .A(n_558), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g565 ( .A(n_559), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g673 ( .A(n_560), .Y(n_673) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_563), .B(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g596 ( .A(n_568), .Y(n_596) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_570), .B(n_605), .Y(n_654) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OR2x2_ASAP7_75t_L g618 ( .A(n_573), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g663 ( .A(n_573), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_574), .A2(n_621), .B1(n_624), .B2(n_626), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g718 ( .A(n_577), .B(n_641), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_582), .B1(n_586), .B2(n_592), .C(n_595), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx2_ASAP7_75t_L g616 ( .A(n_585), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_SL g662 ( .A(n_588), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_590), .B(n_640), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_590), .A2(n_658), .B(n_660), .Y(n_657) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g703 ( .A(n_591), .B(n_685), .Y(n_703) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_SL g605 ( .A(n_594), .Y(n_605) );
AOI21xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_599), .Y(n_595) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g649 ( .A(n_601), .B(n_650), .Y(n_649) );
INVxp67_ASAP7_75t_L g711 ( .A(n_601), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_606), .B(n_607), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_605), .B(n_623), .Y(n_659) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g680 ( .A(n_609), .Y(n_680) );
NAND5xp2_ASAP7_75t_L g610 ( .A(n_611), .B(n_628), .C(n_637), .D(n_657), .E(n_664), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .B(n_617), .C(n_620), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g652 ( .A(n_616), .Y(n_652) );
CKINVDCx16_ASAP7_75t_R g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_624), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g666 ( .A(n_626), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g628 ( .A1(n_629), .A2(n_632), .B(n_634), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_629), .A2(n_683), .B1(n_686), .B2(n_688), .C(n_689), .Y(n_682) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AOI321xp33_ASAP7_75t_L g637 ( .A1(n_630), .A2(n_638), .A3(n_642), .B1(n_643), .B2(n_649), .C(n_651), .Y(n_637) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g708 ( .A(n_642), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_644), .B(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g660 ( .A(n_645), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
NOR2xp67_ASAP7_75t_SL g672 ( .A(n_646), .B(n_653), .Y(n_672) );
AOI321xp33_ASAP7_75t_SL g704 ( .A1(n_649), .A2(n_705), .A3(n_706), .B1(n_707), .B2(n_708), .C(n_709), .Y(n_704) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_654), .C(n_655), .Y(n_651) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_662), .B(n_670), .Y(n_699) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .C(n_674), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_700), .C(n_712), .Y(n_675) );
OAI211xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_678), .B(n_682), .C(n_692), .Y(n_676) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_680), .B(n_681), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_681), .A2(n_713), .B1(n_714), .B2(n_715), .C(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g701 ( .A(n_683), .Y(n_701) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g705 ( .A(n_703), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
CKINVDCx14_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_723), .B(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx3_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .Y(n_738) );
NOR2xp33_ASAP7_75t_SL g739 ( .A(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_SL g766 ( .A(n_740), .Y(n_766) );
INVx1_ASAP7_75t_L g765 ( .A(n_742), .Y(n_765) );
OA21x2_ASAP7_75t_L g768 ( .A1(n_742), .A2(n_766), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g748 ( .A(n_744), .B(n_749), .C(n_754), .Y(n_748) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g759 ( .A(n_745), .Y(n_759) );
BUFx2_ASAP7_75t_L g769 ( .A(n_745), .Y(n_769) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g756 ( .A(n_750), .Y(n_756) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
endmodule