module real_aes_2446_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g521 ( .A(n_0), .B(n_218), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_1), .B(n_109), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_2), .Y(n_125) );
INVx1_ASAP7_75t_L g152 ( .A(n_3), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_4), .B(n_524), .Y(n_543) );
NAND2xp33_ASAP7_75t_SL g514 ( .A(n_5), .B(n_173), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_6), .B(n_186), .Y(n_209) );
INVx1_ASAP7_75t_L g506 ( .A(n_7), .Y(n_506) );
INVx1_ASAP7_75t_L g243 ( .A(n_8), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_9), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_10), .Y(n_260) );
AND2x2_ASAP7_75t_L g541 ( .A(n_11), .B(n_142), .Y(n_541) );
INVx2_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_13), .B(n_108), .C(n_110), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_13), .Y(n_120) );
INVx1_ASAP7_75t_L g219 ( .A(n_14), .Y(n_219) );
AOI221x1_ASAP7_75t_L g509 ( .A1(n_15), .A2(n_175), .B1(n_510), .B2(n_512), .C(n_513), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_16), .B(n_524), .Y(n_577) );
INVx1_ASAP7_75t_L g106 ( .A(n_17), .Y(n_106) );
INVx1_ASAP7_75t_L g216 ( .A(n_18), .Y(n_216) );
INVx1_ASAP7_75t_SL g164 ( .A(n_19), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_20), .B(n_167), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_21), .A2(n_101), .B1(n_103), .B2(n_111), .Y(n_100) );
AOI33xp33_ASAP7_75t_L g234 ( .A1(n_22), .A2(n_50), .A3(n_149), .B1(n_160), .B2(n_235), .B3(n_236), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_23), .A2(n_512), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_24), .B(n_218), .Y(n_546) );
AOI221xp5_ASAP7_75t_SL g586 ( .A1(n_25), .A2(n_40), .B1(n_512), .B2(n_524), .C(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g253 ( .A(n_26), .Y(n_253) );
OR2x2_ASAP7_75t_L g144 ( .A(n_27), .B(n_88), .Y(n_144) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_27), .A2(n_88), .B(n_143), .Y(n_177) );
INVxp67_ASAP7_75t_L g508 ( .A(n_28), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_29), .B(n_221), .Y(n_581) );
AND2x2_ASAP7_75t_L g535 ( .A(n_30), .B(n_141), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_31), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_32), .A2(n_512), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_33), .B(n_221), .Y(n_588) );
AND2x2_ASAP7_75t_L g154 ( .A(n_34), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g159 ( .A(n_34), .Y(n_159) );
AND2x2_ASAP7_75t_L g173 ( .A(n_34), .B(n_152), .Y(n_173) );
INVxp67_ASAP7_75t_L g110 ( .A(n_35), .Y(n_110) );
OR2x6_ASAP7_75t_L g122 ( .A(n_35), .B(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_36), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_37), .B(n_147), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_38), .A2(n_176), .B1(n_182), .B2(n_186), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_39), .B(n_191), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_41), .A2(n_80), .B1(n_157), .B2(n_512), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_42), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_43), .B(n_218), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g789 ( .A1(n_44), .A2(n_788), .B1(n_790), .B2(n_792), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_45), .B(n_193), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_46), .B(n_167), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_47), .Y(n_185) );
AND2x2_ASAP7_75t_L g525 ( .A(n_48), .B(n_141), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_49), .B(n_141), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_51), .B(n_167), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_52), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_52), .A2(n_62), .B1(n_432), .B2(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g150 ( .A(n_53), .Y(n_150) );
INVx1_ASAP7_75t_L g169 ( .A(n_53), .Y(n_169) );
AND2x2_ASAP7_75t_L g285 ( .A(n_54), .B(n_141), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g241 ( .A1(n_55), .A2(n_73), .B1(n_147), .B2(n_157), .C(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_56), .B(n_147), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_57), .B(n_524), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_58), .B(n_176), .Y(n_262) );
AOI21xp5_ASAP7_75t_SL g198 ( .A1(n_59), .A2(n_157), .B(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g562 ( .A(n_60), .B(n_141), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_61), .B(n_221), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_62), .Y(n_807) );
INVx1_ASAP7_75t_L g212 ( .A(n_63), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_64), .B(n_218), .Y(n_560) );
AND2x2_ASAP7_75t_SL g582 ( .A(n_65), .B(n_142), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_66), .A2(n_512), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g283 ( .A(n_67), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_68), .B(n_221), .Y(n_547) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_69), .B(n_193), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_70), .A2(n_157), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g155 ( .A(n_71), .Y(n_155) );
INVx1_ASAP7_75t_L g171 ( .A(n_71), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_72), .B(n_147), .Y(n_237) );
AND2x2_ASAP7_75t_L g174 ( .A(n_74), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g213 ( .A(n_75), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_76), .A2(n_157), .B(n_163), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_77), .A2(n_157), .B(n_188), .C(n_192), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_78), .A2(n_83), .B1(n_147), .B2(n_524), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_79), .B(n_524), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_81), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_82), .B(n_175), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_84), .A2(n_157), .B1(n_232), .B2(n_233), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_85), .B(n_218), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_86), .B(n_218), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_87), .A2(n_512), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g200 ( .A(n_89), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_90), .B(n_221), .Y(n_559) );
AND2x2_ASAP7_75t_L g238 ( .A(n_91), .B(n_175), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_92), .A2(n_251), .B(n_252), .C(n_254), .Y(n_250) );
INVxp67_ASAP7_75t_L g511 ( .A(n_93), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_94), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_95), .B(n_221), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_96), .A2(n_512), .B(n_579), .Y(n_578) );
BUFx2_ASAP7_75t_L g115 ( .A(n_97), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_98), .B(n_167), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_99), .Y(n_788) );
BUFx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx3_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_SL g104 ( .A(n_105), .B(n_107), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_106), .B(n_124), .Y(n_123) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_126), .B(n_796), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_114), .B(n_797), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_117), .A2(n_798), .B(n_808), .Y(n_797) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_125), .Y(n_117) );
BUFx2_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g808 ( .A(n_119), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x6_ASAP7_75t_SL g496 ( .A(n_120), .B(n_122), .Y(n_496) );
OR2x6_ASAP7_75t_SL g787 ( .A(n_120), .B(n_121), .Y(n_787) );
OR2x2_ASAP7_75t_L g795 ( .A(n_120), .B(n_122), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_788), .B(n_789), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_495), .B1(n_497), .B2(n_785), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_130), .A2(n_495), .B1(n_498), .B2(n_791), .Y(n_790) );
AND3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_489), .C(n_492), .Y(n_130) );
NAND5xp2_ASAP7_75t_L g131 ( .A(n_132), .B(n_389), .C(n_419), .D(n_433), .E(n_459), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI21xp33_ASAP7_75t_L g489 ( .A1(n_133), .A2(n_432), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g803 ( .A(n_133), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_338), .Y(n_133) );
NOR3xp33_ASAP7_75t_SL g134 ( .A(n_135), .B(n_286), .C(n_320), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_203), .B(n_225), .C(n_264), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_178), .Y(n_136) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_138), .B(n_276), .Y(n_341) );
AND2x2_ASAP7_75t_L g428 ( .A(n_138), .B(n_206), .Y(n_428) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g224 ( .A(n_139), .B(n_195), .Y(n_224) );
INVx1_ASAP7_75t_L g266 ( .A(n_139), .Y(n_266) );
INVx2_ASAP7_75t_L g271 ( .A(n_139), .Y(n_271) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_139), .Y(n_299) );
INVx1_ASAP7_75t_L g313 ( .A(n_139), .Y(n_313) );
AND2x2_ASAP7_75t_L g317 ( .A(n_139), .B(n_208), .Y(n_317) );
AND2x2_ASAP7_75t_L g398 ( .A(n_139), .B(n_207), .Y(n_398) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_145), .B(n_174), .Y(n_139) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_140), .A2(n_529), .B(n_535), .Y(n_528) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_140), .A2(n_556), .B(n_562), .Y(n_555) );
AO21x2_ASAP7_75t_L g593 ( .A1(n_140), .A2(n_529), .B(n_535), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_141), .Y(n_140) );
OA21x2_ASAP7_75t_L g585 ( .A1(n_141), .A2(n_586), .B(n_590), .Y(n_585) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x4_ASAP7_75t_L g186 ( .A(n_143), .B(n_144), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_156), .Y(n_145) );
INVx1_ASAP7_75t_L g263 ( .A(n_147), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_147), .A2(n_157), .B1(n_505), .B2(n_507), .Y(n_504) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_153), .Y(n_147) );
INVx1_ASAP7_75t_L g183 ( .A(n_148), .Y(n_183) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
OR2x6_ASAP7_75t_L g165 ( .A(n_149), .B(n_161), .Y(n_165) );
INVxp33_ASAP7_75t_L g235 ( .A(n_149), .Y(n_235) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g162 ( .A(n_150), .B(n_152), .Y(n_162) );
AND2x4_ASAP7_75t_L g221 ( .A(n_150), .B(n_170), .Y(n_221) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g512 ( .A(n_154), .B(n_162), .Y(n_512) );
INVx2_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
AND2x6_ASAP7_75t_L g218 ( .A(n_155), .B(n_168), .Y(n_218) );
INVxp67_ASAP7_75t_L g261 ( .A(n_157), .Y(n_261) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
NOR2x1p5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx1_ASAP7_75t_L g236 ( .A(n_160), .Y(n_236) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_SL g163 ( .A1(n_164), .A2(n_165), .B(n_166), .C(n_172), .Y(n_163) );
INVx2_ASAP7_75t_L g191 ( .A(n_165), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_165), .A2(n_172), .B(n_200), .C(n_201), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_165), .A2(n_212), .B1(n_213), .B2(n_214), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_SL g242 ( .A1(n_165), .A2(n_172), .B(n_243), .C(n_244), .Y(n_242) );
INVxp67_ASAP7_75t_L g251 ( .A(n_165), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g282 ( .A1(n_165), .A2(n_172), .B(n_283), .C(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g214 ( .A(n_167), .Y(n_214) );
AND2x4_ASAP7_75t_L g524 ( .A(n_167), .B(n_173), .Y(n_524) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_170), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_172), .A2(n_189), .B(n_190), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_172), .B(n_186), .Y(n_222) );
INVx1_ASAP7_75t_L g232 ( .A(n_172), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_172), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_172), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_172), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_172), .A2(n_559), .B(n_560), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_172), .A2(n_580), .B(n_581), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_172), .A2(n_588), .B(n_589), .Y(n_587) );
INVx5_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_173), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_175), .A2(n_250), .B1(n_255), .B2(n_256), .Y(n_249) );
INVx3_ASAP7_75t_L g256 ( .A(n_175), .Y(n_256) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_176), .B(n_259), .Y(n_258) );
AOI21x1_ASAP7_75t_L g517 ( .A1(n_176), .A2(n_518), .B(n_525), .Y(n_517) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_177), .Y(n_193) );
AND2x4_ASAP7_75t_SL g178 ( .A(n_179), .B(n_194), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g223 ( .A(n_180), .Y(n_223) );
AND2x2_ASAP7_75t_L g267 ( .A(n_180), .B(n_208), .Y(n_267) );
AND2x2_ASAP7_75t_L g288 ( .A(n_180), .B(n_195), .Y(n_288) );
INVx1_ASAP7_75t_L g311 ( .A(n_180), .Y(n_311) );
AND2x4_ASAP7_75t_L g378 ( .A(n_180), .B(n_207), .Y(n_378) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_187), .Y(n_180) );
NOR3xp33_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .C(n_185), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_186), .A2(n_198), .B(n_202), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_186), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_186), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_186), .B(n_511), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_186), .B(n_214), .C(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_186), .A2(n_543), .B(n_544), .Y(n_542) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_192), .A2(n_230), .B(n_238), .Y(n_229) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_192), .A2(n_230), .B(n_238), .Y(n_293) );
AOI21x1_ASAP7_75t_L g550 ( .A1(n_192), .A2(n_551), .B(n_554), .Y(n_550) );
INVx2_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_193), .A2(n_241), .B(n_245), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_193), .A2(n_577), .B(n_578), .Y(n_576) );
AND2x4_ASAP7_75t_L g394 ( .A(n_194), .B(n_311), .Y(n_394) );
OR2x2_ASAP7_75t_L g435 ( .A(n_194), .B(n_436), .Y(n_435) );
NOR2xp67_ASAP7_75t_SL g454 ( .A(n_194), .B(n_327), .Y(n_454) );
NOR2x1_ASAP7_75t_L g472 ( .A(n_194), .B(n_386), .Y(n_472) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2x1_ASAP7_75t_SL g272 ( .A(n_195), .B(n_208), .Y(n_272) );
AND2x4_ASAP7_75t_L g310 ( .A(n_195), .B(n_311), .Y(n_310) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_195), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_195), .B(n_270), .Y(n_348) );
INVx2_ASAP7_75t_L g362 ( .A(n_195), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_195), .B(n_314), .Y(n_384) );
AND2x2_ASAP7_75t_L g476 ( .A(n_195), .B(n_334), .Y(n_476) );
OR2x6_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2x1_ASAP7_75t_L g204 ( .A(n_205), .B(n_224), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_206), .B(n_313), .Y(n_327) );
AND2x2_ASAP7_75t_SL g336 ( .A(n_206), .B(n_316), .Y(n_336) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_223), .Y(n_206) );
INVx1_ASAP7_75t_L g314 ( .A(n_207), .Y(n_314) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g334 ( .A(n_208), .Y(n_334) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_215), .B(n_222), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_214), .B(n_253), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B1(n_219), .B2(n_220), .Y(n_215) );
INVxp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVxp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g367 ( .A(n_223), .Y(n_367) );
INVx2_ASAP7_75t_SL g412 ( .A(n_224), .Y(n_412) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_246), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_227), .B(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g358 ( .A(n_227), .Y(n_358) );
AND2x2_ASAP7_75t_L g482 ( .A(n_227), .B(n_307), .Y(n_482) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_239), .Y(n_227) );
AND2x4_ASAP7_75t_L g295 ( .A(n_228), .B(n_277), .Y(n_295) );
INVx1_ASAP7_75t_L g306 ( .A(n_228), .Y(n_306) );
AND2x2_ASAP7_75t_L g337 ( .A(n_228), .B(n_292), .Y(n_337) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_229), .B(n_240), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_229), .B(n_278), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_231), .B(n_237), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVxp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g275 ( .A(n_240), .Y(n_275) );
AND2x4_ASAP7_75t_L g343 ( .A(n_240), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g355 ( .A(n_240), .Y(n_355) );
INVx1_ASAP7_75t_L g397 ( .A(n_240), .Y(n_397) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_240), .Y(n_409) );
AND2x2_ASAP7_75t_L g425 ( .A(n_240), .B(n_248), .Y(n_425) );
BUFx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g372 ( .A(n_247), .B(n_330), .Y(n_372) );
INVx1_ASAP7_75t_SL g374 ( .A(n_247), .Y(n_374) );
AND2x2_ASAP7_75t_L g395 ( .A(n_247), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g274 ( .A(n_248), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g302 ( .A(n_248), .Y(n_302) );
INVx2_ASAP7_75t_L g308 ( .A(n_248), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_248), .B(n_278), .Y(n_323) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_257), .Y(n_248) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_256), .A2(n_279), .B(n_285), .Y(n_278) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_256), .A2(n_279), .B(n_285), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .B1(n_262), .B2(n_263), .Y(n_257) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .B(n_273), .Y(n_264) );
INVx1_ASAP7_75t_L g404 ( .A(n_265), .Y(n_404) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g324 ( .A(n_267), .Y(n_324) );
AND2x2_ASAP7_75t_L g380 ( .A(n_267), .B(n_316), .Y(n_380) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
INVx1_ASAP7_75t_L g294 ( .A(n_269), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_269), .B(n_310), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_269), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g401 ( .A(n_269), .B(n_394), .Y(n_401) );
AND2x2_ASAP7_75t_L g475 ( .A(n_269), .B(n_476), .Y(n_475) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_270), .Y(n_463) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_271), .Y(n_383) );
AND2x2_ASAP7_75t_L g296 ( .A(n_272), .B(n_297), .Y(n_296) );
OAI21xp33_ASAP7_75t_L g484 ( .A1(n_272), .A2(n_485), .B(n_487), .Y(n_484) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx3_ASAP7_75t_L g370 ( .A(n_274), .Y(n_370) );
NAND2x1_ASAP7_75t_SL g414 ( .A(n_274), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g417 ( .A(n_274), .B(n_295), .Y(n_417) );
AND2x2_ASAP7_75t_L g329 ( .A(n_276), .B(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g466 ( .A(n_276), .B(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g477 ( .A(n_276), .B(n_425), .Y(n_477) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2x1p5_ASAP7_75t_L g353 ( .A(n_277), .B(n_354), .Y(n_353) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g408 ( .A(n_278), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
OAI21xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_300), .B(n_303), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B1(n_295), .B2(n_296), .Y(n_287) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_288), .Y(n_345) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_294), .Y(n_289) );
AND2x2_ASAP7_75t_L g318 ( .A(n_290), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g424 ( .A(n_290), .B(n_425), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_290), .A2(n_443), .B1(n_444), .B2(n_445), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_290), .B(n_451), .Y(n_450) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g307 ( .A(n_292), .B(n_308), .Y(n_307) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_292), .B(n_308), .Y(n_388) );
NOR2x1_ASAP7_75t_L g396 ( .A(n_292), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g344 ( .A(n_293), .Y(n_344) );
AND2x2_ASAP7_75t_L g352 ( .A(n_293), .B(n_308), .Y(n_352) );
INVx1_ASAP7_75t_L g415 ( .A(n_293), .Y(n_415) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2x1_ASAP7_75t_L g333 ( .A(n_298), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g445 ( .A(n_301), .B(n_330), .Y(n_445) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g319 ( .A(n_302), .Y(n_319) );
AND2x2_ASAP7_75t_L g342 ( .A(n_302), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g430 ( .A(n_302), .B(n_337), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_309), .B1(n_315), .B2(n_318), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g438 ( .A(n_305), .B(n_439), .Y(n_438) );
NAND2x1p5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x2_ASAP7_75t_L g468 ( .A(n_308), .B(n_355), .Y(n_468) );
AND2x2_ASAP7_75t_SL g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx2_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
OAI21xp33_ASAP7_75t_SL g481 ( .A1(n_310), .A2(n_482), .B(n_483), .Y(n_481) );
AND2x4_ASAP7_75t_SL g312 ( .A(n_313), .B(n_314), .Y(n_312) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_313), .Y(n_471) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_SL g413 ( .A1(n_316), .A2(n_414), .B(n_416), .C(n_418), .Y(n_413) );
AND2x2_ASAP7_75t_SL g365 ( .A(n_317), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g418 ( .A(n_317), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_317), .B(n_394), .Y(n_458) );
INVx1_ASAP7_75t_SL g325 ( .A(n_318), .Y(n_325) );
AND2x2_ASAP7_75t_L g406 ( .A(n_319), .B(n_343), .Y(n_406) );
INVx1_ASAP7_75t_L g451 ( .A(n_319), .Y(n_451) );
OAI221xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_324), .B1(n_325), .B2(n_326), .C(n_328), .Y(n_320) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_321), .Y(n_440) );
INVx2_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g488 ( .A(n_323), .B(n_331), .Y(n_488) );
OR2x2_ASAP7_75t_L g347 ( .A(n_324), .B(n_348), .Y(n_347) );
NOR2x1_ASAP7_75t_L g360 ( .A(n_324), .B(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_324), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g486 ( .A(n_324), .B(n_383), .Y(n_486) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI32xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .A3(n_335), .B1(n_336), .B2(n_337), .Y(n_328) );
INVx1_ASAP7_75t_L g349 ( .A(n_330), .Y(n_349) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_332), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g444 ( .A(n_333), .Y(n_444) );
OAI22xp33_ASAP7_75t_SL g426 ( .A1(n_335), .A2(n_427), .B1(n_429), .B2(n_431), .Y(n_426) );
INVx1_ASAP7_75t_L g457 ( .A(n_336), .Y(n_457) );
AOI211x1_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_345), .B(n_346), .C(n_363), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_340), .B(n_425), .Y(n_431) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g387 ( .A(n_343), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g453 ( .A(n_343), .Y(n_453) );
OAI222xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B1(n_350), .B2(n_356), .C1(n_357), .C2(n_359), .Y(n_346) );
INVxp67_ASAP7_75t_L g443 ( .A(n_347), .Y(n_443) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_351), .B(n_436), .Y(n_483) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g399 ( .A(n_352), .B(n_396), .Y(n_399) );
INVx3_ASAP7_75t_L g439 ( .A(n_354), .Y(n_439) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g377 ( .A(n_362), .B(n_378), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_368), .B1(n_371), .B2(n_376), .C(n_379), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_365), .A2(n_422), .B(n_424), .Y(n_421) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g375 ( .A(n_369), .Y(n_375) );
OR2x2_ASAP7_75t_L g479 ( .A(n_370), .B(n_415), .Y(n_479) );
NOR2xp67_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_373), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_376), .A2(n_405), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_377), .A2(n_449), .B(n_456), .Y(n_455) );
INVx4_ASAP7_75t_L g386 ( .A(n_378), .Y(n_386) );
OAI31xp33_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_381), .A3(n_385), .B(n_387), .Y(n_379) );
INVx1_ASAP7_75t_L g437 ( .A(n_381), .Y(n_437) );
NOR2x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g411 ( .A(n_386), .Y(n_411) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_402), .Y(n_389) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_390), .B(n_402), .C(n_421), .D(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_400), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B1(n_398), .B2(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g462 ( .A(n_394), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_395), .B(n_415), .Y(n_423) );
INVx1_ASAP7_75t_SL g436 ( .A(n_398), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_413), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_407), .B2(n_410), .Y(n_403) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2x1_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_412), .A2(n_475), .B1(n_477), .B2(n_478), .Y(n_474) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_426), .C(n_432), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g491 ( .A(n_426), .Y(n_491) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g492 ( .A1(n_432), .A2(n_493), .B(n_494), .Y(n_492) );
INVxp33_ASAP7_75t_L g493 ( .A(n_433), .Y(n_493) );
AND2x2_ASAP7_75t_L g802 ( .A(n_433), .B(n_459), .Y(n_802) );
NOR2xp67_ASAP7_75t_L g433 ( .A(n_434), .B(n_441), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_438), .B2(n_440), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_438), .A2(n_461), .B(n_464), .Y(n_460) );
INVx2_ASAP7_75t_L g448 ( .A(n_439), .Y(n_448) );
NAND3xp33_ASAP7_75t_SL g441 ( .A(n_442), .B(n_446), .C(n_455), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_449), .B1(n_452), .B2(n_454), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVxp33_ASAP7_75t_SL g494 ( .A(n_459), .Y(n_494) );
NOR3x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_473), .C(n_480), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_481), .B(n_484), .Y(n_480) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g804 ( .A(n_490), .Y(n_804) );
CKINVDCx11_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_662), .Y(n_498) );
NOR4xp25_ASAP7_75t_L g499 ( .A(n_500), .B(n_605), .C(n_644), .D(n_651), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_526), .B1(n_563), .B2(n_572), .C(n_591), .Y(n_500) );
OR2x2_ASAP7_75t_L g735 ( .A(n_501), .B(n_597), .Y(n_735) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g650 ( .A(n_502), .B(n_575), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_502), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_SL g715 ( .A(n_502), .B(n_716), .Y(n_715) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_515), .Y(n_502) );
AND2x4_ASAP7_75t_SL g574 ( .A(n_503), .B(n_575), .Y(n_574) );
INVx3_ASAP7_75t_L g596 ( .A(n_503), .Y(n_596) );
AND2x2_ASAP7_75t_L g631 ( .A(n_503), .B(n_604), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_503), .B(n_516), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_503), .B(n_598), .Y(n_683) );
OR2x2_ASAP7_75t_L g761 ( .A(n_503), .B(n_575), .Y(n_761) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .Y(n_503) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g583 ( .A(n_516), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_516), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g609 ( .A(n_516), .Y(n_609) );
OR2x2_ASAP7_75t_L g614 ( .A(n_516), .B(n_598), .Y(n_614) );
AND2x2_ASAP7_75t_L g627 ( .A(n_516), .B(n_585), .Y(n_627) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_516), .Y(n_630) );
INVx1_ASAP7_75t_L g642 ( .A(n_516), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_516), .B(n_596), .Y(n_707) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_527), .B(n_536), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g571 ( .A(n_528), .B(n_555), .Y(n_571) );
AND2x4_ASAP7_75t_L g601 ( .A(n_528), .B(n_540), .Y(n_601) );
INVx2_ASAP7_75t_L g635 ( .A(n_528), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_528), .B(n_555), .Y(n_693) );
AND2x2_ASAP7_75t_L g740 ( .A(n_528), .B(n_569), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
AOI222xp33_ASAP7_75t_L g728 ( .A1(n_536), .A2(n_600), .B1(n_643), .B2(n_703), .C1(n_729), .C2(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_548), .Y(n_537) );
AND2x2_ASAP7_75t_L g647 ( .A(n_538), .B(n_567), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_538), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g776 ( .A(n_538), .B(n_616), .Y(n_776) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_539), .A2(n_607), .B(n_611), .Y(n_606) );
AND2x2_ASAP7_75t_L g687 ( .A(n_539), .B(n_570), .Y(n_687) );
OR2x2_ASAP7_75t_L g712 ( .A(n_539), .B(n_571), .Y(n_712) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx5_ASAP7_75t_L g566 ( .A(n_540), .Y(n_566) );
AND2x2_ASAP7_75t_L g653 ( .A(n_540), .B(n_635), .Y(n_653) );
AND2x2_ASAP7_75t_L g679 ( .A(n_540), .B(n_555), .Y(n_679) );
OR2x2_ASAP7_75t_L g682 ( .A(n_540), .B(n_569), .Y(n_682) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_540), .Y(n_700) );
AND2x4_ASAP7_75t_SL g757 ( .A(n_540), .B(n_634), .Y(n_757) );
OR2x2_ASAP7_75t_L g766 ( .A(n_540), .B(n_593), .Y(n_766) );
OR2x6_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g599 ( .A(n_548), .Y(n_599) );
AOI221xp5_ASAP7_75t_SL g717 ( .A1(n_548), .A2(n_601), .B1(n_718), .B2(n_720), .C(n_721), .Y(n_717) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_555), .Y(n_548) );
OR2x2_ASAP7_75t_L g656 ( .A(n_549), .B(n_626), .Y(n_656) );
OR2x2_ASAP7_75t_L g666 ( .A(n_549), .B(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g692 ( .A(n_549), .B(n_693), .Y(n_692) );
AND2x4_ASAP7_75t_L g698 ( .A(n_549), .B(n_617), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_549), .B(n_681), .Y(n_710) );
INVx2_ASAP7_75t_L g723 ( .A(n_549), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_549), .B(n_601), .Y(n_744) );
AND2x2_ASAP7_75t_L g748 ( .A(n_549), .B(n_570), .Y(n_748) );
AND2x2_ASAP7_75t_L g756 ( .A(n_549), .B(n_757), .Y(n_756) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g569 ( .A(n_550), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_555), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g600 ( .A(n_555), .B(n_569), .Y(n_600) );
INVx2_ASAP7_75t_L g617 ( .A(n_555), .Y(n_617) );
AND2x4_ASAP7_75t_L g634 ( .A(n_555), .B(n_635), .Y(n_634) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_555), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g746 ( .A(n_565), .B(n_568), .Y(n_746) );
AND2x4_ASAP7_75t_L g592 ( .A(n_566), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g633 ( .A(n_566), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g660 ( .A(n_566), .B(n_600), .Y(n_660) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
AND2x2_ASAP7_75t_L g764 ( .A(n_568), .B(n_765), .Y(n_764) );
BUFx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g616 ( .A(n_569), .B(n_617), .Y(n_616) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_570), .A2(n_637), .B(n_643), .Y(n_636) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_583), .Y(n_573) );
INVx1_ASAP7_75t_SL g690 ( .A(n_574), .Y(n_690) );
AND2x2_ASAP7_75t_L g720 ( .A(n_574), .B(n_630), .Y(n_720) );
AND2x4_ASAP7_75t_L g731 ( .A(n_574), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g597 ( .A(n_575), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g604 ( .A(n_575), .Y(n_604) );
AND2x4_ASAP7_75t_L g610 ( .A(n_575), .B(n_596), .Y(n_610) );
INVx2_ASAP7_75t_L g621 ( .A(n_575), .Y(n_621) );
INVx1_ASAP7_75t_L g670 ( .A(n_575), .Y(n_670) );
OR2x2_ASAP7_75t_L g691 ( .A(n_575), .B(n_675), .Y(n_691) );
OR2x2_ASAP7_75t_L g705 ( .A(n_575), .B(n_585), .Y(n_705) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_575), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_575), .B(n_627), .Y(n_777) );
OR2x6_ASAP7_75t_L g575 ( .A(n_576), .B(n_582), .Y(n_575) );
INVx1_ASAP7_75t_L g622 ( .A(n_583), .Y(n_622) );
AND2x2_ASAP7_75t_L g755 ( .A(n_583), .B(n_621), .Y(n_755) );
AND2x2_ASAP7_75t_L g780 ( .A(n_583), .B(n_610), .Y(n_780) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g598 ( .A(n_585), .Y(n_598) );
BUFx3_ASAP7_75t_L g640 ( .A(n_585), .Y(n_640) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_585), .Y(n_667) );
INVx1_ASAP7_75t_L g676 ( .A(n_585), .Y(n_676) );
AOI33xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .A3(n_599), .B1(n_600), .B2(n_601), .B3(n_602), .Y(n_591) );
AOI21x1_ASAP7_75t_SL g694 ( .A1(n_592), .A2(n_616), .B(n_678), .Y(n_694) );
INVx2_ASAP7_75t_L g724 ( .A(n_592), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_592), .B(n_723), .Y(n_730) );
AND2x2_ASAP7_75t_L g678 ( .A(n_593), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g641 ( .A(n_596), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g742 ( .A(n_597), .Y(n_742) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_598), .Y(n_732) );
OAI32xp33_ASAP7_75t_L g781 ( .A1(n_599), .A2(n_601), .A3(n_777), .B1(n_782), .B2(n_784), .Y(n_781) );
AND2x2_ASAP7_75t_L g699 ( .A(n_600), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g689 ( .A(n_601), .Y(n_689) );
AND2x2_ASAP7_75t_L g754 ( .A(n_601), .B(n_698), .Y(n_754) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_615), .B1(n_618), .B2(n_632), .C(n_636), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_609), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_610), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_610), .B(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_610), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g659 ( .A(n_614), .Y(n_659) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_623), .C(n_628), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g721 ( .A1(n_620), .A2(n_682), .B1(n_722), .B2(n_725), .Y(n_721) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g625 ( .A(n_621), .Y(n_625) );
NOR2x1p5_ASAP7_75t_L g639 ( .A(n_621), .B(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_621), .Y(n_661) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI322xp33_ASAP7_75t_L g688 ( .A1(n_624), .A2(n_666), .A3(n_689), .B1(n_690), .B2(n_691), .C1(n_692), .C2(n_694), .Y(n_688) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_626), .A2(n_645), .B(n_646), .C(n_648), .Y(n_644) );
OR2x2_ASAP7_75t_L g736 ( .A(n_626), .B(n_690), .Y(n_736) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g643 ( .A(n_627), .B(n_631), .Y(n_643) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g649 ( .A(n_633), .B(n_650), .Y(n_649) );
INVx3_ASAP7_75t_SL g681 ( .A(n_634), .Y(n_681) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_638), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_SL g685 ( .A(n_641), .Y(n_685) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_642), .Y(n_727) );
OR2x6_ASAP7_75t_SL g782 ( .A(n_645), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g772 ( .A1(n_650), .A2(n_773), .B(n_774), .C(n_781), .Y(n_772) );
O2A1O1Ixp33_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_654), .B(n_657), .C(n_661), .Y(n_651) );
OAI211xp5_ASAP7_75t_SL g663 ( .A1(n_652), .A2(n_664), .B(n_671), .C(n_695), .Y(n_663) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_708), .C(n_752), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_667), .Y(n_759) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g714 ( .A(n_670), .Y(n_714) );
NOR3xp33_ASAP7_75t_SL g671 ( .A(n_672), .B(n_684), .C(n_688), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_677), .B1(n_680), .B2(n_683), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g716 ( .A(n_676), .Y(n_716) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_676), .Y(n_783) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_SL g769 ( .A(n_682), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
OR2x2_ASAP7_75t_L g719 ( .A(n_685), .B(n_705), .Y(n_719) );
OR2x2_ASAP7_75t_L g770 ( .A(n_685), .B(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g768 ( .A(n_693), .Y(n_768) );
OR2x2_ASAP7_75t_L g784 ( .A(n_693), .B(n_723), .Y(n_784) );
OAI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_699), .B(n_701), .Y(n_695) );
OAI31xp33_ASAP7_75t_L g709 ( .A1(n_696), .A2(n_710), .A3(n_711), .B(n_713), .Y(n_709) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g741 ( .A(n_706), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND4xp25_ASAP7_75t_SL g708 ( .A(n_709), .B(n_717), .C(n_728), .D(n_733), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_716), .Y(n_751) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_737), .B1(n_741), .B2(n_743), .C(n_745), .Y(n_733) );
NAND2xp33_ASAP7_75t_SL g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g778 ( .A(n_737), .Y(n_778) );
AND2x2_ASAP7_75t_SL g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g773 ( .A(n_747), .Y(n_773) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_753), .B(n_772), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B1(n_756), .B2(n_758), .C(n_762), .Y(n_753) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
AOI21xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_767), .B(n_770), .Y(n_762) );
INVxp33_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_786), .Y(n_791) );
CKINVDCx11_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
INVx3_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI22xp33_ASAP7_75t_SL g798 ( .A1(n_799), .A2(n_800), .B1(n_805), .B2(n_806), .Y(n_798) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NAND3x1_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .C(n_804), .Y(n_801) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
endmodule