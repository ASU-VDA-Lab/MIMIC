module fake_jpeg_507_n_597 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_597);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_597;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_18),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_59),
.Y(n_153)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g146 ( 
.A(n_61),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_66),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_70),
.Y(n_135)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_75),
.Y(n_147)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_87),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_20),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_76),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_77),
.Y(n_193)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_78),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_80),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_81),
.A2(n_26),
.B1(n_47),
.B2(n_43),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_82),
.Y(n_197)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_84),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_33),
.B(n_2),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_89),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_92),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_24),
.B(n_2),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_102),
.Y(n_143)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_95),
.Y(n_179)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_96),
.Y(n_216)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_98),
.Y(n_187)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_99),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

INVx11_ASAP7_75t_SL g101 ( 
.A(n_25),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_3),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_25),
.Y(n_104)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_109),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_33),
.B(n_4),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_111),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_33),
.B(n_4),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

CKINVDCx11_ASAP7_75t_R g114 ( 
.A(n_33),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_21),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_29),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_121),
.Y(n_169)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_118),
.B(n_123),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_21),
.Y(n_119)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_24),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_124),
.B(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_27),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_125),
.B(n_126),
.Y(n_183)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_27),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_59),
.B(n_55),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_128),
.B(n_130),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_35),
.B(n_28),
.C(n_47),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_82),
.B(n_35),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_131),
.B(n_154),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_38),
.B1(n_54),
.B2(n_44),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_132),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_103),
.A2(n_88),
.B1(n_116),
.B2(n_36),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_134),
.A2(n_16),
.B(n_132),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_62),
.A2(n_51),
.B1(n_44),
.B2(n_40),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_62),
.A2(n_51),
.B1(n_40),
.B2(n_36),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_141),
.B(n_177),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_60),
.A2(n_117),
.B1(n_76),
.B2(n_90),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_142),
.A2(n_164),
.B1(n_182),
.B2(n_207),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_30),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_90),
.B(n_32),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_155),
.B(n_162),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_32),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_43),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_163),
.B(n_174),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_L g164 ( 
.A1(n_69),
.A2(n_41),
.B1(n_28),
.B2(n_26),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_95),
.B(n_41),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_120),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_65),
.B(n_42),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_178),
.B(n_184),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_100),
.A2(n_42),
.B1(n_23),
.B2(n_9),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_124),
.B(n_23),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_67),
.B(n_6),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_16),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_96),
.B(n_6),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_194),
.B(n_198),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_79),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_217),
.B1(n_159),
.B2(n_152),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_97),
.B(n_8),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_85),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_206),
.B(n_214),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_91),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_100),
.A2(n_113),
.B1(n_105),
.B2(n_98),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_209),
.A2(n_211),
.B1(n_213),
.B2(n_181),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_61),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_210),
.A2(n_211),
.B1(n_182),
.B2(n_134),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_66),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_66),
.A2(n_71),
.B1(n_13),
.B2(n_14),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_71),
.B(n_10),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_89),
.A2(n_15),
.B1(n_16),
.B2(n_92),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_15),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_218),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_219),
.B(n_250),
.Y(n_321)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_148),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_220),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g327 ( 
.A(n_221),
.B(n_269),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_222),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_143),
.B(n_150),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_223),
.B(n_255),
.Y(n_310)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_224),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_187),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_225),
.B(n_242),
.C(n_244),
.Y(n_339)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_226),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_130),
.A2(n_200),
.B(n_169),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_228),
.A2(n_292),
.B(n_208),
.Y(n_317)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_151),
.Y(n_229)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_229),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_230),
.A2(n_235),
.B1(n_248),
.B2(n_218),
.Y(n_330)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_186),
.B(n_203),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_234),
.B(n_288),
.Y(n_340)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_237),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_156),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_239),
.Y(n_308)
);

OR2x2_ASAP7_75t_SL g240 ( 
.A(n_133),
.B(n_149),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_240),
.Y(n_300)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_157),
.Y(n_242)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_156),
.Y(n_243)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_161),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_246),
.Y(n_337)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_247),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_166),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_248),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_147),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_251),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_252),
.A2(n_167),
.B1(n_176),
.B2(n_204),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_165),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_253),
.Y(n_341)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_254),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_129),
.B(n_190),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_256),
.Y(n_347)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_257),
.Y(n_349)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_259),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_168),
.B(n_170),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_260),
.B(n_275),
.Y(n_315)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_160),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_271),
.Y(n_312)
);

BUFx12_ASAP7_75t_L g262 ( 
.A(n_146),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_262),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_158),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_263),
.B(n_267),
.Y(n_334)
);

AND2x2_ASAP7_75t_SL g266 ( 
.A(n_212),
.B(n_173),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_144),
.C(n_195),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_146),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_175),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_135),
.B(n_145),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_160),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_153),
.B(n_191),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_272),
.B(n_276),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_165),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_273),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_164),
.B(n_200),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_175),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_197),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_278),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_153),
.B(n_191),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_171),
.B(n_173),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_279),
.B(n_281),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_186),
.B(n_203),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_280),
.B(n_282),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_179),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_197),
.Y(n_283)
);

NOR3xp33_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_285),
.C(n_286),
.Y(n_320)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_167),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_171),
.Y(n_286)
);

AO22x2_ASAP7_75t_L g287 ( 
.A1(n_215),
.A2(n_172),
.B1(n_209),
.B2(n_142),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_136),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_173),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_266),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_139),
.A2(n_213),
.B(n_137),
.C(n_193),
.Y(n_292)
);

AO22x2_ASAP7_75t_L g293 ( 
.A1(n_172),
.A2(n_195),
.B1(n_144),
.B2(n_193),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_293),
.A2(n_192),
.B1(n_205),
.B2(n_284),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_295),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_223),
.B(n_179),
.C(n_176),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_299),
.B(n_304),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_302),
.A2(n_289),
.B1(n_245),
.B2(n_293),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_204),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_275),
.A2(n_192),
.B1(n_205),
.B2(n_208),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_313),
.A2(n_331),
.B1(n_350),
.B2(n_280),
.Y(n_353)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_288),
.A2(n_264),
.A3(n_228),
.B1(n_219),
.B2(n_260),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_338),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_317),
.A2(n_329),
.B(n_333),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_322),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_235),
.A2(n_227),
.B1(n_258),
.B2(n_265),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_324),
.A2(n_330),
.B1(n_257),
.B2(n_226),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_236),
.A2(n_252),
.B1(n_233),
.B2(n_274),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_255),
.A2(n_221),
.B1(n_287),
.B2(n_248),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_332),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_292),
.A2(n_287),
.B1(n_280),
.B2(n_218),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_266),
.B(n_240),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_232),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_345),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_287),
.A2(n_261),
.B1(n_271),
.B2(n_282),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_329),
.A2(n_220),
.B1(n_285),
.B2(n_243),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_352),
.A2(n_353),
.B1(n_366),
.B2(n_367),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_331),
.A2(n_269),
.B1(n_247),
.B2(n_253),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_354),
.A2(n_371),
.B1(n_374),
.B2(n_295),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_241),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_364),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_290),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_357),
.B(n_368),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_327),
.A2(n_234),
.B(n_293),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_358),
.A2(n_390),
.B(n_394),
.Y(n_410)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_344),
.Y(n_360)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_361),
.Y(n_409)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_325),
.Y(n_362)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_362),
.Y(n_414)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_363),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_311),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_297),
.B(n_237),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_378),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_315),
.A2(n_222),
.B1(n_273),
.B2(n_238),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_293),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_370),
.B(n_373),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_315),
.A2(n_302),
.B1(n_317),
.B2(n_313),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_304),
.B(n_299),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_340),
.A2(n_256),
.B1(n_239),
.B2(n_259),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_297),
.B(n_232),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_375),
.B(n_376),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_296),
.B(n_262),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_312),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_312),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_381),
.Y(n_420)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_325),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_307),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_333),
.A2(n_262),
.B1(n_340),
.B2(n_316),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_384),
.A2(n_391),
.B1(n_320),
.B2(n_335),
.Y(n_412)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_386),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_334),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_387),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_303),
.B(n_321),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_388),
.B(n_389),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_332),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_296),
.B(n_323),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_337),
.A2(n_314),
.B1(n_338),
.B2(n_300),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_308),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_392),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_312),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_393),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_328),
.B(n_298),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_371),
.A2(n_337),
.B1(n_319),
.B2(n_348),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_398),
.A2(n_402),
.B1(n_379),
.B2(n_383),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_400),
.B(n_412),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_353),
.A2(n_348),
.B1(n_298),
.B2(n_309),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_372),
.C(n_373),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_405),
.B(n_408),
.C(n_411),
.Y(n_433)
);

OAI32xp33_ASAP7_75t_L g406 ( 
.A1(n_351),
.A2(n_346),
.A3(n_342),
.B1(n_336),
.B2(n_349),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_413),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_359),
.B(n_372),
.C(n_357),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_351),
.B(n_346),
.Y(n_411)
);

OAI32xp33_ASAP7_75t_L g413 ( 
.A1(n_368),
.A2(n_342),
.A3(n_336),
.B1(n_349),
.B2(n_305),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_365),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_425),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_356),
.A2(n_335),
.B(n_308),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_419),
.A2(n_423),
.B(n_428),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_356),
.A2(n_318),
.B(n_347),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_384),
.B(n_389),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_426),
.C(n_405),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_394),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_318),
.C(n_305),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_377),
.A2(n_301),
.B1(n_341),
.B2(n_294),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_427),
.A2(n_354),
.B1(n_367),
.B2(n_377),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_391),
.A2(n_347),
.B(n_306),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_419),
.A2(n_358),
.B(n_393),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_434),
.A2(n_456),
.B(n_455),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_435),
.A2(n_441),
.B1(n_443),
.B2(n_446),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_425),
.B(n_386),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_436),
.B(n_444),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_448),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_411),
.C(n_424),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_445),
.C(n_454),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_420),
.Y(n_439)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_440),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_400),
.A2(n_352),
.B1(n_366),
.B2(n_363),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_395),
.B(n_380),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_361),
.C(n_360),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_398),
.B1(n_407),
.B2(n_402),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_414),
.Y(n_447)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_388),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_407),
.A2(n_378),
.B1(n_374),
.B2(n_364),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_449),
.A2(n_404),
.B1(n_403),
.B2(n_415),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_395),
.B(n_410),
.Y(n_450)
);

AOI21xp33_ASAP7_75t_L g469 ( 
.A1(n_450),
.A2(n_452),
.B(n_453),
.Y(n_469)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_414),
.Y(n_451)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_376),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_401),
.B(n_390),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_397),
.B(n_375),
.C(n_355),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_423),
.A2(n_392),
.B(n_362),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_401),
.B(n_381),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_457),
.A2(n_430),
.B1(n_341),
.B2(n_294),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_397),
.B(n_422),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_459),
.C(n_461),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_406),
.B(n_385),
.Y(n_459)
);

OA22x2_ASAP7_75t_L g460 ( 
.A1(n_412),
.A2(n_382),
.B1(n_369),
.B2(n_301),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_460),
.B(n_462),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_326),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_399),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_464),
.A2(n_485),
.B1(n_460),
.B2(n_430),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_404),
.Y(n_465)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_465),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_433),
.B(n_415),
.C(n_409),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_470),
.B(n_480),
.C(n_488),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_426),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_445),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_432),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_473),
.B(n_487),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_418),
.Y(n_474)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_474),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_431),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_477),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_462),
.B(n_417),
.Y(n_478)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_478),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_442),
.A2(n_428),
.B1(n_399),
.B2(n_409),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_479),
.A2(n_482),
.B1(n_449),
.B2(n_441),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_437),
.B(n_429),
.C(n_417),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_442),
.A2(n_421),
.B1(n_427),
.B2(n_429),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_447),
.Y(n_483)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_483),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_442),
.A2(n_421),
.B1(n_413),
.B2(n_396),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_451),
.Y(n_486)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_486),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_456),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_396),
.C(n_306),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_431),
.Y(n_489)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_489),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_491),
.A2(n_455),
.B(n_434),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_460),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_497),
.C(n_467),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_448),
.C(n_454),
.Y(n_497)
);

OAI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_498),
.A2(n_504),
.B1(n_514),
.B2(n_485),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_459),
.Y(n_499)
);

CKINVDCx14_ASAP7_75t_R g533 ( 
.A(n_499),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_480),
.B(n_458),
.Y(n_500)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_500),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_503),
.A2(n_463),
.B(n_469),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_465),
.B(n_461),
.Y(n_506)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_506),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_470),
.B(n_326),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_507),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_446),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_510),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_468),
.B(n_443),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_512),
.A2(n_479),
.B1(n_466),
.B2(n_486),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_482),
.A2(n_460),
.B1(n_369),
.B2(n_382),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_491),
.A2(n_416),
.B(n_294),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_515),
.A2(n_463),
.B(n_487),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_478),
.Y(n_516)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_516),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_489),
.A2(n_307),
.B1(n_416),
.B2(n_473),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_517),
.A2(n_476),
.B1(n_481),
.B2(n_416),
.Y(n_534)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_518),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_519),
.B(n_503),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_505),
.B(n_475),
.Y(n_521)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_521),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_522),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_524),
.B(n_525),
.Y(n_540)
);

AOI322xp5_ASAP7_75t_L g525 ( 
.A1(n_513),
.A2(n_474),
.A3(n_475),
.B1(n_477),
.B2(n_484),
.C1(n_466),
.C2(n_464),
.Y(n_525)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_526),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_488),
.C(n_472),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_527),
.B(n_529),
.C(n_536),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_483),
.Y(n_528)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_528),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_494),
.B(n_467),
.C(n_468),
.Y(n_529)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_534),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_502),
.B(n_476),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_535),
.B(n_506),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_493),
.B(n_481),
.C(n_497),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g538 ( 
.A1(n_518),
.A2(n_501),
.B(n_495),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_538),
.A2(n_548),
.B(n_549),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_532),
.B(n_508),
.Y(n_543)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_543),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_521),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_544),
.B(n_530),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_526),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_504),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_547),
.A2(n_531),
.B(n_520),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_535),
.A2(n_495),
.B(n_502),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_527),
.B(n_536),
.C(n_524),
.Y(n_552)
);

NOR2xp67_ASAP7_75t_SL g562 ( 
.A(n_552),
.B(n_510),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_529),
.C(n_523),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_553),
.B(n_557),
.Y(n_572)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_554),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_542),
.A2(n_551),
.B1(n_514),
.B2(n_537),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_558),
.B(n_561),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_523),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_559),
.B(n_560),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_539),
.B(n_519),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_551),
.A2(n_501),
.B1(n_498),
.B2(n_496),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_562),
.B(n_546),
.C(n_549),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_540),
.B(n_520),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_563),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_541),
.A2(n_533),
.B1(n_531),
.B2(n_501),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_564),
.B(n_537),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_538),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_566),
.B(n_554),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_567),
.A2(n_568),
.B1(n_557),
.B2(n_561),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_563),
.B(n_546),
.C(n_539),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_569),
.B(n_570),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_538),
.C(n_550),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_515),
.C(n_517),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_571),
.B(n_555),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_576),
.B(n_556),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_578),
.B(n_581),
.Y(n_587)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_572),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_579),
.B(n_580),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_574),
.A2(n_555),
.B(n_560),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_582),
.B(n_583),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_573),
.B(n_574),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_584),
.B(n_568),
.C(n_575),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_585),
.B(n_588),
.Y(n_590)
);

BUFx24_ASAP7_75t_SL g588 ( 
.A(n_577),
.Y(n_588)
);

OAI21xp33_ASAP7_75t_L g591 ( 
.A1(n_587),
.A2(n_586),
.B(n_589),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_591),
.A2(n_592),
.B(n_545),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_586),
.A2(n_579),
.B(n_583),
.Y(n_592)
);

OAI21xp33_ASAP7_75t_L g595 ( 
.A1(n_593),
.A2(n_594),
.B(n_528),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_590),
.B(n_511),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_595),
.B(n_509),
.C(n_571),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_596),
.B(n_534),
.Y(n_597)
);


endmodule