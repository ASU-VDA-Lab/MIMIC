module fake_jpeg_16684_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_43),
.B(n_47),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_29),
.B(n_16),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_0),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_61),
.B1(n_21),
.B2(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_1),
.C(n_2),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_17),
.B1(n_37),
.B2(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_15),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_34),
.B1(n_17),
.B2(n_19),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_81),
.B1(n_32),
.B2(n_28),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_57),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_34),
.B1(n_19),
.B2(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_75),
.B1(n_79),
.B2(n_35),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_34),
.B1(n_19),
.B2(n_37),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_20),
.B1(n_24),
.B2(n_35),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_21),
.B1(n_18),
.B2(n_26),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_42),
.A2(n_18),
.B1(n_26),
.B2(n_28),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_35),
.B1(n_23),
.B2(n_32),
.Y(n_98)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_56),
.B1(n_39),
.B2(n_41),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_63),
.B1(n_67),
.B2(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_95),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_98),
.B1(n_101),
.B2(n_103),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_114),
.B1(n_117),
.B2(n_63),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_61),
.A3(n_43),
.B1(n_45),
.B2(n_62),
.Y(n_97)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_83),
.A3(n_63),
.B1(n_26),
.B2(n_36),
.Y(n_118)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_102),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_50),
.B1(n_52),
.B2(n_39),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_55),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_83),
.B1(n_78),
.B2(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_105),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

BUFx2_ASAP7_75t_SL g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_47),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_113),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_57),
.B(n_49),
.C(n_70),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_112),
.A2(n_85),
.B(n_36),
.C(n_27),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_24),
.B1(n_20),
.B2(n_32),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_41),
.B1(n_48),
.B2(n_76),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_54),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_116),
.B(n_77),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_30),
.B1(n_26),
.B2(n_28),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_126),
.B(n_128),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_139),
.B1(n_96),
.B2(n_107),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_28),
.B(n_85),
.Y(n_126)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_101),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_94),
.B1(n_114),
.B2(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_103),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_150),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_153),
.B1(n_130),
.B2(n_129),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_100),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_104),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_148),
.Y(n_162)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_97),
.A3(n_92),
.B1(n_112),
.B2(n_91),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_155),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_113),
.C(n_105),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_137),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_115),
.B1(n_112),
.B2(n_91),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_141),
.B1(n_147),
.B2(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_116),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_102),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_152),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_98),
.A3(n_116),
.B1(n_109),
.B2(n_106),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_159),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_108),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_176),
.B1(n_120),
.B2(n_130),
.Y(n_195)
);

OAI221xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_131),
.B1(n_132),
.B2(n_128),
.C(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_161),
.B(n_31),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_168),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_121),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_170),
.C(n_173),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_132),
.Y(n_170)
);

CKINVDCx12_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_139),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_157),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_175),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_121),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_121),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_178),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_146),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_153),
.B1(n_152),
.B2(n_151),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_195),
.B1(n_48),
.B2(n_51),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_90),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_149),
.B1(n_150),
.B2(n_148),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_166),
.B1(n_172),
.B2(n_163),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_134),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_194),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_99),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_201),
.B(n_202),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_129),
.B1(n_136),
.B2(n_123),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_203),
.B1(n_162),
.B2(n_168),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_163),
.B(n_136),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_199),
.B(n_172),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_123),
.C(n_125),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_174),
.C(n_171),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_179),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_129),
.B(n_89),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_125),
.B1(n_96),
.B2(n_89),
.Y(n_203)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_199),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_208),
.B1(n_183),
.B2(n_192),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_166),
.B1(n_173),
.B2(n_174),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_212),
.C(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_179),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_77),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_31),
.B(n_38),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_214),
.A2(n_219),
.B1(n_202),
.B2(n_184),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_77),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_93),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_2),
.B(n_3),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_191),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_223),
.B(n_224),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_199),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_219),
.A2(n_198),
.B1(n_195),
.B2(n_203),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_233),
.B1(n_220),
.B2(n_221),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_230),
.Y(n_254)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_231),
.C(n_234),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_190),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_189),
.C(n_184),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_185),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_185),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_245)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_201),
.C(n_187),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_210),
.B(n_222),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_SL g258 ( 
.A1(n_246),
.A2(n_249),
.B(n_224),
.C(n_223),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_226),
.CI(n_236),
.CON(n_247),
.SN(n_247)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_27),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_210),
.B(n_211),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_238),
.A2(n_205),
.B1(n_217),
.B2(n_204),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_251),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_217),
.B1(n_204),
.B2(n_215),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_214),
.B(n_216),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_255),
.B(n_256),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_230),
.C(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_84),
.C(n_65),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_SL g255 ( 
.A(n_232),
.B(n_218),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_213),
.B(n_191),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_250),
.B1(n_245),
.B2(n_254),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_247),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_269),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_197),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_264),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_SL g263 ( 
.A1(n_241),
.A2(n_191),
.A3(n_15),
.B1(n_13),
.B2(n_11),
.C1(n_27),
.C2(n_36),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_265),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_15),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_84),
.C(n_65),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_267),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_53),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_44),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_243),
.A2(n_11),
.B1(n_13),
.B2(n_38),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_270),
.A2(n_252),
.B1(n_246),
.B2(n_249),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_244),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_276),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_279),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_256),
.Y(n_276)
);

NAND2x1_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_258),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_242),
.C(n_254),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_93),
.C(n_65),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_245),
.B1(n_253),
.B2(n_76),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_282),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_5),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_2),
.B(n_3),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_51),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_74),
.B(n_38),
.Y(n_287)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_74),
.B(n_51),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_4),
.B(n_5),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_271),
.A3(n_277),
.B1(n_274),
.B2(n_281),
.C1(n_280),
.C2(n_44),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_4),
.B(n_5),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_4),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_295),
.B(n_6),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_283),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_299),
.B(n_289),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_5),
.B(n_6),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_293),
.B(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_301),
.B(n_304),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_300),
.A2(n_292),
.B(n_297),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_302),
.A2(n_286),
.B(n_8),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_305),
.C(n_306),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_7),
.B(n_8),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_311),
.C(n_308),
.Y(n_312)
);

AOI221xp5_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_7),
.B1(n_9),
.B2(n_301),
.C(n_298),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_7),
.Y(n_313)
);


endmodule