module fake_netlist_6_1831_n_783 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_783);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_783;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_575;
wire n_368;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_601;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_153;
wire n_758;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_600;
wire n_464;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_6),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_136),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_92),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_75),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_30),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_31),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_1),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_10),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_10),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_2),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_39),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_3),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_33),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_64),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_48),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_16),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_45),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_66),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_121),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_133),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_44),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_94),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_90),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_112),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_57),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_16),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_141),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_131),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_114),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_43),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_142),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_49),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_89),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_54),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_117),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_24),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_99),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_71),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_88),
.Y(n_201)
);

BUFx8_ASAP7_75t_SL g202 ( 
.A(n_155),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_146),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_27),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_0),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_0),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_1),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_28),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_L g216 ( 
.A(n_145),
.B(n_2),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

BUFx8_ASAP7_75t_SL g221 ( 
.A(n_164),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_151),
.B(n_3),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_29),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_4),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_149),
.B(n_4),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_152),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_160),
.B(n_5),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_168),
.B(n_5),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_167),
.B(n_32),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_149),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_149),
.B(n_195),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_6),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_233),
.A2(n_227),
.B1(n_238),
.B2(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_201),
.B1(n_200),
.B2(n_150),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_196),
.B1(n_192),
.B2(n_179),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_231),
.B1(n_219),
.B2(n_243),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_210),
.B(n_153),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_176),
.B1(n_191),
.B2(n_189),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_210),
.B(n_154),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_205),
.A2(n_184),
.B1(n_188),
.B2(n_187),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_210),
.B(n_159),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_204),
.A2(n_175),
.B1(n_183),
.B2(n_181),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_204),
.A2(n_180),
.B1(n_173),
.B2(n_172),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_161),
.B1(n_170),
.B2(n_9),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

BUFx6f_ASAP7_75t_SL g266 ( 
.A(n_212),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_211),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_211),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_207),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_195),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_205),
.A2(n_195),
.B1(n_12),
.B2(n_13),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_206),
.A2(n_195),
.B1(n_12),
.B2(n_13),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_213),
.A2(n_195),
.B1(n_14),
.B2(n_15),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_213),
.A2(n_195),
.B1(n_14),
.B2(n_15),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_206),
.A2(n_11),
.B1(n_17),
.B2(n_18),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_212),
.B(n_34),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_216),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_222),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_209),
.B(n_35),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_209),
.A2(n_241),
.B1(n_208),
.B2(n_229),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_221),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

AO22x2_ASAP7_75t_L g286 ( 
.A1(n_223),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_228),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_229),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_234),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_234),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_234),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g292 ( 
.A1(n_208),
.A2(n_41),
.B1(n_42),
.B2(n_46),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_228),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g295 ( 
.A(n_250),
.B(n_223),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_245),
.A2(n_223),
.B(n_217),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_247),
.A2(n_217),
.B(n_242),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_258),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_242),
.Y(n_301)
);

NAND2x1p5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_214),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_251),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_263),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_242),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_254),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_256),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_214),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_253),
.Y(n_319)
);

NAND2xp33_ASAP7_75t_SL g320 ( 
.A(n_266),
.B(n_264),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_266),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_245),
.A2(n_252),
.B(n_255),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_248),
.B(n_242),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_248),
.B(n_214),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_265),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_271),
.B(n_214),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_259),
.B(n_244),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_259),
.B(n_228),
.Y(n_336)
);

INVxp33_ASAP7_75t_SL g337 ( 
.A(n_262),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_273),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_273),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_276),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_249),
.B(n_202),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_277),
.B(n_218),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_276),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_262),
.B(n_244),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_267),
.B(n_230),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_268),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_275),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_254),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_R g351 ( 
.A(n_245),
.B(n_47),
.Y(n_351)
);

NAND2x1p5_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_230),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_261),
.B(n_230),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_246),
.B(n_202),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_261),
.B(n_230),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_275),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_282),
.B(n_235),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_282),
.B(n_235),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_275),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_296),
.B(n_226),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_345),
.Y(n_361)
);

AND2x2_ASAP7_75t_SL g362 ( 
.A(n_307),
.B(n_357),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_303),
.Y(n_364)
);

AND2x4_ASAP7_75t_SL g365 ( 
.A(n_345),
.B(n_235),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_318),
.B(n_235),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_306),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_236),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

NOR2x1_ASAP7_75t_L g372 ( 
.A(n_307),
.B(n_327),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_236),
.Y(n_374)
);

INVx3_ASAP7_75t_SL g375 ( 
.A(n_322),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_236),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_300),
.B(n_50),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_304),
.Y(n_379)
);

AND2x2_ASAP7_75t_SL g380 ( 
.A(n_338),
.B(n_226),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_339),
.B(n_340),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_239),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_304),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_317),
.B(n_236),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_299),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_305),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_308),
.B(n_220),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_301),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_350),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_315),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_321),
.B(n_327),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_294),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_344),
.B(n_343),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_312),
.B(n_239),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_297),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_336),
.B(n_239),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_334),
.B(n_346),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_347),
.B(n_239),
.Y(n_401)
);

BUFx4_ASAP7_75t_SL g402 ( 
.A(n_348),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_220),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_295),
.B(n_237),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_336),
.B(n_220),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_335),
.B(n_237),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_326),
.B(n_237),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_314),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_356),
.B(n_51),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_359),
.B(n_237),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_352),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_332),
.B(n_330),
.Y(n_415)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_311),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_330),
.B(n_52),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_309),
.B(n_53),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_316),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_298),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_333),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_325),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_333),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_337),
.B(n_55),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_323),
.B(n_56),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_328),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

BUFx8_ASAP7_75t_L g428 ( 
.A(n_324),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_302),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_362),
.B(n_302),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_419),
.Y(n_431)
);

BUFx4f_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_370),
.B(n_342),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_407),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_354),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_362),
.B(n_320),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_379),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_398),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_392),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_362),
.B(n_58),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_59),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_428),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_351),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_351),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_407),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_361),
.B(n_394),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_407),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_407),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_361),
.B(n_60),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_363),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_400),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_401),
.B(n_61),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_398),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_394),
.B(n_62),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_394),
.B(n_65),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_401),
.B(n_67),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_403),
.B(n_68),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_400),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_412),
.B(n_69),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_364),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_381),
.Y(n_469)
);

AND2x2_ASAP7_75t_SL g470 ( 
.A(n_424),
.B(n_70),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_72),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_403),
.B(n_74),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_415),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_364),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_414),
.B(n_423),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_373),
.B(n_429),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_414),
.B(n_76),
.Y(n_478)
);

BUFx4f_ASAP7_75t_L g479 ( 
.A(n_377),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_415),
.B(n_78),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_80),
.Y(n_481)
);

AND2x2_ASAP7_75t_SL g482 ( 
.A(n_380),
.B(n_414),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_393),
.B(n_81),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_381),
.Y(n_484)
);

CKINVDCx8_ASAP7_75t_R g485 ( 
.A(n_377),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_372),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_441),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_474),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_396),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_441),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_451),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_451),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_454),
.Y(n_494)
);

BUFx4_ASAP7_75t_SL g495 ( 
.A(n_444),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_434),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_451),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_431),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_476),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_434),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_472),
.Y(n_501)
);

NAND2x1p5_ASAP7_75t_L g502 ( 
.A(n_472),
.B(n_377),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_447),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_434),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_447),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_456),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_479),
.A2(n_423),
.B1(n_380),
.B2(n_421),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_465),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_437),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_444),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_430),
.A2(n_426),
.B1(n_425),
.B2(n_380),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_435),
.Y(n_512)
);

BUFx8_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_470),
.A2(n_423),
.B1(n_421),
.B2(n_425),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_469),
.B(n_396),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_438),
.Y(n_516)
);

BUFx5_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_437),
.Y(n_518)
);

BUFx8_ASAP7_75t_L g519 ( 
.A(n_443),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_437),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_472),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_437),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_484),
.B(n_389),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_476),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_440),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_449),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_449),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_436),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_480),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_449),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_458),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_510),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_514),
.A2(n_485),
.B1(n_430),
.B2(n_479),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_517),
.A2(n_470),
.B1(n_482),
.B2(n_428),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_510),
.Y(n_536)
);

CKINVDCx11_ASAP7_75t_R g537 ( 
.A(n_487),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_495),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_511),
.A2(n_485),
.B1(n_479),
.B2(n_432),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_486),
.A2(n_445),
.B1(n_446),
.B2(n_442),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_489),
.Y(n_541)
);

OAI22x1_ASAP7_75t_L g542 ( 
.A1(n_529),
.A2(n_512),
.B1(n_486),
.B2(n_530),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_487),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_501),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_490),
.A2(n_377),
.B1(n_481),
.B2(n_471),
.Y(n_545)
);

BUFx12f_ASAP7_75t_L g546 ( 
.A(n_523),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_523),
.A2(n_418),
.B1(n_477),
.B2(n_481),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_502),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_491),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_498),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_506),
.Y(n_551)
);

OAI22xp33_ASAP7_75t_L g552 ( 
.A1(n_515),
.A2(n_467),
.B1(n_432),
.B2(n_408),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_494),
.A2(n_432),
.B1(n_429),
.B2(n_481),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_503),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_501),
.Y(n_555)
);

INVx6_ASAP7_75t_L g556 ( 
.A(n_509),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_503),
.Y(n_557)
);

OAI22xp33_ASAP7_75t_L g558 ( 
.A1(n_494),
.A2(n_471),
.B1(n_466),
.B2(n_452),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_491),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_508),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_509),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_490),
.A2(n_428),
.B1(n_382),
.B2(n_466),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_505),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_516),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_492),
.A2(n_471),
.B1(n_466),
.B2(n_454),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_526),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_502),
.A2(n_449),
.B1(n_452),
.B2(n_453),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_492),
.A2(n_454),
.B1(n_460),
.B2(n_459),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_507),
.A2(n_452),
.B1(n_453),
.B2(n_459),
.Y(n_569)
);

CKINVDCx11_ASAP7_75t_R g570 ( 
.A(n_488),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_493),
.A2(n_452),
.B1(n_453),
.B2(n_459),
.Y(n_571)
);

CKINVDCx6p67_ASAP7_75t_R g572 ( 
.A(n_509),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_505),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_532),
.A2(n_428),
.B1(n_382),
.B2(n_360),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_517),
.A2(n_519),
.B1(n_513),
.B2(n_460),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_493),
.Y(n_576)
);

OAI21xp33_ASAP7_75t_L g577 ( 
.A1(n_547),
.A2(n_387),
.B(n_409),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_570),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_535),
.A2(n_519),
.B1(n_412),
.B2(n_513),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_535),
.A2(n_519),
.B1(n_513),
.B2(n_517),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_576),
.B(n_390),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_560),
.B(n_409),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_534),
.A2(n_517),
.B1(n_460),
.B2(n_478),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_550),
.Y(n_584)
);

CKINVDCx11_ASAP7_75t_R g585 ( 
.A(n_533),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_564),
.Y(n_586)
);

BUFx12f_ASAP7_75t_L g587 ( 
.A(n_537),
.Y(n_587)
);

INVx5_ASAP7_75t_SL g588 ( 
.A(n_572),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_574),
.A2(n_517),
.B1(n_497),
.B2(n_524),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_539),
.A2(n_546),
.B1(n_517),
.B2(n_536),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_540),
.B(n_517),
.Y(n_591)
);

BUFx5_ASAP7_75t_L g592 ( 
.A(n_566),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_SL g593 ( 
.A1(n_549),
.A2(n_478),
.B1(n_499),
.B2(n_524),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_554),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_540),
.B(n_497),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_543),
.A2(n_525),
.B1(n_499),
.B2(n_360),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_557),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_568),
.A2(n_525),
.B1(n_453),
.B2(n_509),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_559),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_563),
.Y(n_600)
);

OAI21xp33_ASAP7_75t_L g601 ( 
.A1(n_574),
.A2(n_562),
.B(n_542),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_562),
.A2(n_462),
.B1(n_473),
.B2(n_365),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_573),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_541),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_575),
.A2(n_365),
.B1(n_457),
.B2(n_461),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_541),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_575),
.A2(n_365),
.B1(n_483),
.B2(n_405),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_544),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_545),
.A2(n_565),
.B1(n_552),
.B2(n_558),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_558),
.A2(n_509),
.B1(n_501),
.B2(n_521),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_544),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_569),
.A2(n_521),
.B1(n_369),
.B2(n_374),
.Y(n_612)
);

BUFx12f_ASAP7_75t_L g613 ( 
.A(n_538),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_571),
.A2(n_521),
.B1(n_376),
.B2(n_427),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_555),
.Y(n_615)
);

NOR2x1_ASAP7_75t_R g616 ( 
.A(n_556),
.B(n_402),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_555),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_553),
.Y(n_618)
);

OAI222xp33_ASAP7_75t_L g619 ( 
.A1(n_552),
.A2(n_399),
.B1(n_417),
.B2(n_406),
.C1(n_368),
.C2(n_366),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_551),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_SL g621 ( 
.A1(n_548),
.A2(n_417),
.B1(n_496),
.B2(n_527),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_548),
.A2(n_531),
.B1(n_528),
.B2(n_527),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_551),
.A2(n_405),
.B1(n_411),
.B2(n_404),
.Y(n_623)
);

OAI21xp33_ASAP7_75t_SL g624 ( 
.A1(n_567),
.A2(n_504),
.B(n_518),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_556),
.A2(n_427),
.B1(n_528),
.B2(n_527),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_601),
.A2(n_411),
.B1(n_405),
.B2(n_395),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_609),
.A2(n_596),
.B1(n_579),
.B2(n_593),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_580),
.A2(n_375),
.B1(n_556),
.B2(n_561),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_577),
.A2(n_411),
.B1(n_395),
.B2(n_386),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_590),
.A2(n_395),
.B1(n_386),
.B2(n_368),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_SL g631 ( 
.A1(n_598),
.A2(n_561),
.B1(n_531),
.B2(n_528),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_583),
.A2(n_395),
.B1(n_386),
.B2(n_385),
.Y(n_632)
);

AOI221xp5_ASAP7_75t_L g633 ( 
.A1(n_619),
.A2(n_384),
.B1(n_420),
.B2(n_386),
.C(n_385),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_589),
.A2(n_385),
.B1(n_388),
.B2(n_420),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_591),
.B(n_488),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_595),
.A2(n_388),
.B1(n_367),
.B2(n_416),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_582),
.A2(n_388),
.B1(n_367),
.B2(n_416),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_618),
.A2(n_367),
.B1(n_416),
.B2(n_375),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_594),
.B(n_500),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_621),
.B(n_488),
.Y(n_640)
);

BUFx6f_ASAP7_75t_SL g641 ( 
.A(n_578),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_597),
.B(n_500),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_598),
.A2(n_375),
.B1(n_475),
.B2(n_468),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_591),
.A2(n_416),
.B1(n_383),
.B2(n_379),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_600),
.B(n_603),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_602),
.A2(n_416),
.B1(n_383),
.B2(n_410),
.Y(n_646)
);

AOI221xp5_ASAP7_75t_L g647 ( 
.A1(n_581),
.A2(n_413),
.B1(n_397),
.B2(n_475),
.C(n_468),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_584),
.B(n_520),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_586),
.B(n_488),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_607),
.A2(n_416),
.B1(n_383),
.B2(n_504),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_605),
.A2(n_416),
.B1(n_504),
.B2(n_518),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_578),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_599),
.A2(n_606),
.B1(n_604),
.B2(n_620),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_585),
.A2(n_416),
.B1(n_518),
.B2(n_371),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_592),
.A2(n_416),
.B1(n_371),
.B2(n_364),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_623),
.A2(n_561),
.B1(n_520),
.B2(n_528),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_592),
.A2(n_578),
.B1(n_610),
.B2(n_612),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_622),
.A2(n_528),
.B1(n_527),
.B2(n_522),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_592),
.A2(n_371),
.B1(n_364),
.B2(n_439),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_610),
.A2(n_531),
.B1(n_527),
.B2(n_522),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_608),
.B(n_455),
.Y(n_661)
);

OAI222xp33_ASAP7_75t_L g662 ( 
.A1(n_625),
.A2(n_464),
.B1(n_439),
.B2(n_448),
.C1(n_455),
.C2(n_371),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_592),
.A2(n_464),
.B1(n_439),
.B2(n_488),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_592),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_611),
.B(n_448),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_645),
.B(n_592),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_664),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_635),
.B(n_649),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_635),
.B(n_615),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_649),
.B(n_617),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_664),
.B(n_631),
.Y(n_671)
);

OAI21xp33_ASAP7_75t_L g672 ( 
.A1(n_627),
.A2(n_614),
.B(n_624),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_648),
.B(n_614),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_657),
.A2(n_588),
.B1(n_625),
.B2(n_587),
.Y(n_674)
);

NAND3xp33_ASAP7_75t_L g675 ( 
.A(n_626),
.B(n_531),
.C(n_522),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_643),
.B(n_531),
.C(n_522),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_SL g677 ( 
.A(n_641),
.B(n_522),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_639),
.B(n_616),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_642),
.B(n_588),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_660),
.B(n_588),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_640),
.B(n_464),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_640),
.B(n_82),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_630),
.A2(n_613),
.B1(n_463),
.B2(n_378),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_643),
.A2(n_463),
.B1(n_378),
.B2(n_86),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_644),
.B(n_84),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_652),
.B(n_85),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_653),
.B(n_87),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_661),
.B(n_91),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_665),
.B(n_652),
.Y(n_689)
);

AND2x2_ASAP7_75t_SL g690 ( 
.A(n_632),
.B(n_463),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_634),
.B(n_93),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_628),
.A2(n_463),
.B1(n_378),
.B2(n_97),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_651),
.A2(n_378),
.B1(n_96),
.B2(n_98),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_658),
.B(n_95),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_638),
.B(n_378),
.C(n_101),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_636),
.B(n_100),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_R g697 ( 
.A(n_682),
.B(n_641),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_667),
.Y(n_698)
);

OAI211xp5_ASAP7_75t_L g699 ( 
.A1(n_672),
.A2(n_687),
.B(n_673),
.C(n_682),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_695),
.B(n_647),
.C(n_637),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_668),
.B(n_656),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_667),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_670),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_674),
.A2(n_641),
.B1(n_650),
.B2(n_654),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_692),
.A2(n_646),
.B1(n_629),
.B2(n_633),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_684),
.A2(n_655),
.B1(n_659),
.B2(n_663),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_676),
.B(n_688),
.C(n_666),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_678),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_669),
.B(n_104),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_689),
.B(n_106),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_L g711 ( 
.A(n_679),
.B(n_662),
.C(n_109),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_671),
.B(n_107),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_671),
.B(n_110),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_681),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_702),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_703),
.B(n_681),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_714),
.B(n_680),
.Y(n_717)
);

NAND4xp75_ASAP7_75t_L g718 ( 
.A(n_713),
.B(n_694),
.C(n_680),
.D(n_686),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_702),
.Y(n_719)
);

NOR2x1_ASAP7_75t_L g720 ( 
.A(n_707),
.B(n_699),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_714),
.B(n_694),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_698),
.B(n_690),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_708),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_701),
.Y(n_724)
);

XNOR2x2_ASAP7_75t_L g725 ( 
.A(n_700),
.B(n_675),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_701),
.B(n_690),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_719),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_724),
.B(n_713),
.Y(n_728)
);

XNOR2xp5_ASAP7_75t_L g729 ( 
.A(n_718),
.B(n_708),
.Y(n_729)
);

XNOR2x1_ASAP7_75t_L g730 ( 
.A(n_720),
.B(n_712),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_715),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_724),
.B(n_721),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_730),
.A2(n_729),
.B1(n_718),
.B2(n_697),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_730),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_732),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_732),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_736),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_735),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_734),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_733),
.Y(n_740)
);

AOI22x1_ASAP7_75t_L g741 ( 
.A1(n_739),
.A2(n_725),
.B1(n_726),
.B2(n_727),
.Y(n_741)
);

OA22x2_ASAP7_75t_L g742 ( 
.A1(n_739),
.A2(n_728),
.B1(n_726),
.B2(n_725),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_740),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_743),
.Y(n_744)
);

OAI221xp5_ASAP7_75t_L g745 ( 
.A1(n_741),
.A2(n_737),
.B1(n_738),
.B2(n_723),
.C(n_704),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_742),
.A2(n_723),
.B1(n_722),
.B2(n_677),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_743),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_744),
.A2(n_677),
.B1(n_722),
.B2(n_721),
.Y(n_748)
);

NOR2x1_ASAP7_75t_L g749 ( 
.A(n_747),
.B(n_686),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_746),
.B(n_731),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_745),
.B(n_717),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_744),
.A2(n_710),
.B1(n_711),
.B2(n_709),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_751),
.A2(n_716),
.B1(n_715),
.B2(n_705),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_750),
.B(n_696),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_749),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_748),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_752),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_750),
.B(n_691),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_755),
.Y(n_759)
);

AO22x2_ASAP7_75t_L g760 ( 
.A1(n_757),
.A2(n_696),
.B1(n_685),
.B2(n_683),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_756),
.A2(n_685),
.B1(n_706),
.B2(n_693),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_758),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_753),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_759),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_762),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_763),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_761),
.B(n_754),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_760),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_765),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_766),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_764),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_SL g772 ( 
.A1(n_768),
.A2(n_760),
.B1(n_115),
.B2(n_116),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_770),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_769),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_771),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_775),
.A2(n_767),
.B1(n_772),
.B2(n_119),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_774),
.A2(n_767),
.B1(n_118),
.B2(n_120),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_773),
.A2(n_111),
.B1(n_122),
.B2(n_123),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_776),
.Y(n_779)
);

OA22x2_ASAP7_75t_L g780 ( 
.A1(n_779),
.A2(n_777),
.B1(n_778),
.B2(n_126),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_780),
.Y(n_781)
);

AOI221xp5_ASAP7_75t_L g782 ( 
.A1(n_781),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.C(n_128),
.Y(n_782)
);

AOI211xp5_ASAP7_75t_L g783 ( 
.A1(n_782),
.A2(n_130),
.B(n_132),
.C(n_134),
.Y(n_783)
);


endmodule