module real_jpeg_30351_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_0),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_0),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_1),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_18)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_1),
.A2(n_23),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_1),
.A2(n_23),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_2),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_5),
.B(n_62),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_5),
.A2(n_104),
.A3(n_111),
.B1(n_113),
.B2(n_118),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_5),
.A2(n_119),
.B1(n_145),
.B2(n_149),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_5),
.A2(n_74),
.B1(n_183),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_6),
.A2(n_98),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_7),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_7),
.A2(n_52),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_8),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

INVx2_ASAP7_75t_R g84 ( 
.A(n_8),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_8),
.A2(n_84),
.B1(n_165),
.B2(n_168),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_10),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_11),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_11),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_178),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_176),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_101),
.Y(n_14)
);

NOR2xp67_ASAP7_75t_SL g177 ( 
.A(n_15),
.B(n_101),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_60),
.C(n_73),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_16),
.A2(n_60),
.B1(n_61),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_16),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_28),
.B1(n_49),
.B2(n_58),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_18),
.A2(n_172),
.B1(n_234),
.B2(n_237),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_22),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_28),
.Y(n_172)
);

AO21x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_37),
.B(n_41),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_36),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_37),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_43),
.Y(n_129)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_43),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_43),
.Y(n_231)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_49),
.Y(n_173)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_58),
.B(n_119),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_58),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_59),
.Y(n_171)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AO21x2_ASAP7_75t_L g135 ( 
.A1(n_63),
.A2(n_113),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_65),
.Y(n_170)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_73),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_78),
.B1(n_88),
.B2(n_93),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_74),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_74),
.A2(n_125),
.B1(n_183),
.B2(n_189),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_78),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_87),
.Y(n_195)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_88),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_123),
.B1(n_124),
.B2(n_127),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_133),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_122),
.B1(n_131),
.B2(n_132),
.Y(n_102)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_119),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_119),
.B(n_226),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_SL g234 ( 
.A1(n_119),
.A2(n_225),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_123),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_208)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_163),
.B1(n_174),
.B2(n_175),
.Y(n_133)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_144),
.B1(n_152),
.B2(n_153),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_241),
.B(n_246),
.Y(n_178)
);

AOI22x1_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_207),
.B1(n_239),
.B2(n_240),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_197),
.B(n_206),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_196),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_182),
.B(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_233),
.B2(n_238),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_213),
.B(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_224),
.B1(n_230),
.B2(n_232),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);


endmodule