module fake_jpeg_12645_n_194 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_17),
.Y(n_58)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_23),
.B1(n_22),
.B2(n_31),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_37),
.B1(n_23),
.B2(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_61),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_33),
.B1(n_16),
.B2(n_19),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_21),
.B1(n_26),
.B2(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_19),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_68),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_43),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_16),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_69),
.A2(n_82),
.B1(n_84),
.B2(n_50),
.Y(n_103)
);

AOI32xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_21),
.A3(n_40),
.B1(n_44),
.B2(n_30),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_49),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_76),
.C(n_59),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_45),
.C(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_35),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_31),
.B1(n_28),
.B2(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_33),
.B1(n_37),
.B2(n_48),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_30),
.B(n_21),
.C(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_86),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_26),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_62),
.C(n_63),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_97),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_104),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_62),
.C(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_11),
.Y(n_101)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_75),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_85),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_69),
.B1(n_68),
.B2(n_86),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_122),
.B1(n_123),
.B2(n_94),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_115),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_14),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_99),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_67),
.B(n_1),
.Y(n_120)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_124),
.B(n_126),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_87),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_78),
.B1(n_74),
.B2(n_79),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_75),
.B1(n_56),
.B2(n_51),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_67),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_50),
.B(n_2),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_115),
.A2(n_87),
.B1(n_93),
.B2(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_136),
.B1(n_123),
.B2(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_138),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_124),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_122),
.C(n_18),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_141),
.B1(n_109),
.B2(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_94),
.B1(n_106),
.B2(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_104),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_104),
.B1(n_39),
.B2(n_18),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_135),
.A2(n_119),
.B1(n_113),
.B2(n_125),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_147),
.B1(n_148),
.B2(n_5),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_134),
.B(n_137),
.C(n_127),
.D(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_11),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_152),
.B1(n_131),
.B2(n_130),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_3),
.C(n_5),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_157),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_160),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_138),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_162),
.B(n_163),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_137),
.B(n_131),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_10),
.C(n_12),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_152),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_154),
.B(n_145),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_155),
.B1(n_12),
.B2(n_13),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_166),
.A2(n_168),
.B1(n_6),
.B2(n_7),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_176),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_148),
.B1(n_155),
.B2(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_173),
.A2(n_174),
.B1(n_166),
.B2(n_162),
.Y(n_179)
);

AOI31xp67_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_5),
.A3(n_6),
.B(n_7),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_175),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_160),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_8),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_178),
.B1(n_182),
.B2(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_163),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_170),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_184),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_186),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_183),
.B(n_186),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_189),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_190),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_192),
.Y(n_194)
);


endmodule