module fake_jpeg_15562_n_302 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_SL g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_14),
.B(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_33),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_59),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_31),
.B1(n_34),
.B2(n_30),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_30),
.B1(n_33),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_33),
.B1(n_25),
.B2(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_16),
.B1(n_15),
.B2(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_24),
.B1(n_25),
.B2(n_23),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_25),
.B1(n_23),
.B2(n_20),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_42),
.B1(n_39),
.B2(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_20),
.B1(n_19),
.B2(n_29),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_38),
.B(n_46),
.C(n_39),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_24),
.B1(n_20),
.B2(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_53),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_69),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_46),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_46),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_67),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_41),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_40),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_62),
.B(n_48),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_38),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_44),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_64),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_101),
.B(n_70),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_44),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_99),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_106),
.B(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_29),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_57),
.B1(n_38),
.B2(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_75),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_63),
.B(n_18),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_116),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_82),
.B(n_72),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_92),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_117),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_123),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_72),
.B(n_82),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_120),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_82),
.C(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_84),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_126),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_84),
.C(n_78),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_95),
.C(n_97),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_158),
.C(n_109),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_147),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_152),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_110),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_151),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_111),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_127),
.B(n_101),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_94),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_157),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_130),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_105),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_105),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_153),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_185),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_120),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_106),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_168),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_115),
.B1(n_120),
.B2(n_124),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_169),
.B1(n_174),
.B2(n_175),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_125),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_115),
.B1(n_127),
.B2(n_114),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_138),
.C(n_134),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_114),
.B1(n_112),
.B2(n_116),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_113),
.B1(n_117),
.B2(n_84),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_182),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_121),
.B1(n_95),
.B2(n_131),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_180),
.B1(n_137),
.B2(n_101),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_121),
.B1(n_89),
.B2(n_103),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_186),
.Y(n_207)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_189),
.C(n_190),
.Y(n_217)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_99),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_119),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_192),
.B(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_136),
.C(n_144),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_195),
.C(n_196),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_136),
.C(n_144),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_137),
.C(n_140),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_198),
.B(n_73),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_203),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_174),
.B(n_133),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_171),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_205),
.B(n_103),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_133),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_208),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_98),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_71),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_204),
.A2(n_182),
.B1(n_179),
.B2(n_168),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_211),
.A2(n_216),
.B1(n_78),
.B2(n_70),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_199),
.A2(n_166),
.B1(n_173),
.B2(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_195),
.B1(n_193),
.B2(n_197),
.Y(n_216)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_222),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_224),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_180),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_228),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_173),
.B1(n_186),
.B2(n_176),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_191),
.A2(n_139),
.B(n_143),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_226),
.A2(n_83),
.B(n_170),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_229),
.Y(n_243)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_192),
.B(n_208),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_219),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_216),
.C(n_217),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_234),
.C(n_221),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_225),
.A2(n_185),
.B1(n_170),
.B2(n_148),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_241),
.B1(n_0),
.B2(n_1),
.Y(n_251)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_214),
.A3(n_217),
.B1(n_210),
.B2(n_223),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_0),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_143),
.C(n_147),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_245),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_78),
.B1(n_71),
.B2(n_69),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_71),
.B1(n_57),
.B2(n_24),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_57),
.B1(n_63),
.B2(n_22),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_257),
.C(n_239),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_212),
.C(n_213),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_255),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_256),
.B(n_247),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_245),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_22),
.B(n_21),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_11),
.C(n_1),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_29),
.C(n_22),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_21),
.B1(n_17),
.B2(n_16),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_258),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_17),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_252),
.B(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_238),
.B1(n_236),
.B2(n_230),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_270),
.B1(n_15),
.B2(n_2),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_236),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_18),
.Y(n_279)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_246),
.B1(n_2),
.B2(n_3),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_241),
.C(n_242),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_18),
.B(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_277),
.C(n_278),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_267),
.A2(n_21),
.B(n_16),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_283)
);

NOR3xp33_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_0),
.C(n_2),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_266),
.C(n_263),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_279),
.C(n_275),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_268),
.C(n_264),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_265),
.C(n_4),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_3),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_288),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_3),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_289),
.C(n_292),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_293),
.B(n_5),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_4),
.B(n_5),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_10),
.C(n_5),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_10),
.B(n_5),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_4),
.B(n_6),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_6),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_302)
);


endmodule