module fake_jpeg_7478_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_18),
.B1(n_35),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_42),
.B1(n_19),
.B2(n_17),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_18),
.B1(n_35),
.B2(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_19),
.B1(n_17),
.B2(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_78),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_42),
.B1(n_18),
.B2(n_21),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_22),
.B1(n_34),
.B2(n_31),
.Y(n_112)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_42),
.B1(n_47),
.B2(n_44),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_81),
.B1(n_83),
.B2(n_31),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_86),
.B1(n_20),
.B2(n_21),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_80),
.B(n_84),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_39),
.B1(n_19),
.B2(n_17),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_37),
.B1(n_39),
.B2(n_20),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_68),
.B1(n_64),
.B2(n_59),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_50),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_111),
.C(n_121),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_109),
.B1(n_112),
.B2(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_37),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_113),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_41),
.C(n_44),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_87),
.B1(n_88),
.B2(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_R g115 ( 
.A(n_77),
.B(n_39),
.Y(n_115)
);

XNOR2x2_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_36),
.Y(n_147)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_119),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_71),
.A2(n_34),
.B1(n_22),
.B2(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_48),
.C(n_44),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_68),
.B1(n_64),
.B2(n_59),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_58),
.B1(n_92),
.B2(n_25),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g131 ( 
.A(n_104),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_75),
.B1(n_76),
.B2(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_132),
.A2(n_120),
.B1(n_116),
.B2(n_108),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_90),
.B1(n_89),
.B2(n_96),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_150),
.B1(n_99),
.B2(n_103),
.Y(n_177)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_141),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_75),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_120),
.B(n_47),
.Y(n_184)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_145),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_115),
.B(n_114),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_147),
.B(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_96),
.C(n_94),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_127),
.C(n_102),
.Y(n_163)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_152),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_91),
.B1(n_94),
.B2(n_58),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_91),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_102),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_138),
.B(n_139),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_160),
.B(n_162),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_112),
.B(n_25),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_122),
.B(n_125),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_143),
.C(n_146),
.Y(n_188)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_177),
.Y(n_190)
);

OAI22x1_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_27),
.B1(n_99),
.B2(n_23),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_175),
.B1(n_123),
.B2(n_140),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_170),
.B(n_172),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_36),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_182),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_28),
.B(n_29),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_184),
.B(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_24),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_48),
.B(n_47),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_182),
.B1(n_180),
.B2(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_192),
.C(n_198),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_189),
.B(n_191),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_164),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_149),
.Y(n_192)
);

AOI22x1_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_139),
.B1(n_133),
.B2(n_148),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_175),
.B1(n_181),
.B2(n_123),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_195),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_145),
.C(n_136),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_29),
.B(n_30),
.C(n_33),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_214),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_133),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_208),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_217),
.B(n_28),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_184),
.B(n_187),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_162),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_211),
.B1(n_213),
.B2(n_215),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_48),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_154),
.B1(n_108),
.B2(n_153),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_166),
.B1(n_175),
.B2(n_165),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_41),
.C(n_140),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_171),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_171),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_167),
.C(n_179),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_218),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_165),
.B1(n_178),
.B2(n_177),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_222),
.B1(n_228),
.B2(n_234),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_220),
.A2(n_221),
.B1(n_227),
.B2(n_209),
.Y(n_256)
);

OAI22x1_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_169),
.B1(n_159),
.B2(n_185),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_199),
.A2(n_177),
.B1(n_170),
.B2(n_167),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_232),
.B(n_238),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_158),
.B1(n_185),
.B2(n_161),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_190),
.A2(n_158),
.B1(n_160),
.B2(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_181),
.B(n_161),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_231),
.B(n_243),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_214),
.B(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_23),
.B1(n_26),
.B2(n_41),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_23),
.B1(n_26),
.B2(n_2),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_24),
.B(n_23),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_0),
.B(n_1),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_200),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_16),
.C(n_15),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_209),
.B(n_168),
.CI(n_26),
.CON(n_244),
.SN(n_244)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_210),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_188),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_224),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_208),
.C(n_212),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_249),
.C(n_255),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_212),
.C(n_198),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_217),
.B1(n_202),
.B2(n_203),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_252),
.A2(n_263),
.B1(n_235),
.B2(n_229),
.Y(n_284)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_234),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_192),
.C(n_206),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_206),
.C(n_205),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_260),
.B(n_229),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_0),
.C(n_2),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_266),
.C(n_239),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_0),
.C(n_2),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_274),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_241),
.B(n_242),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_270),
.B1(n_281),
.B2(n_284),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_278),
.C(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_233),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_271),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g272 ( 
.A(n_251),
.B(n_224),
.CI(n_221),
.CON(n_272),
.SN(n_272)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_272),
.B(n_282),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_238),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_265),
.Y(n_291)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_279),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_235),
.C(n_220),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_227),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_280),
.A2(n_246),
.B1(n_245),
.B2(n_263),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_231),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_244),
.B(n_12),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_269),
.C(n_295),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_292),
.B1(n_296),
.B2(n_284),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_257),
.B(n_256),
.C(n_261),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_290),
.A2(n_282),
.B(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_271),
.A2(n_264),
.B1(n_257),
.B2(n_250),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_249),
.B(n_238),
.Y(n_293)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_280),
.A2(n_244),
.B1(n_247),
.B2(n_13),
.Y(n_296)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_12),
.C(n_11),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_3),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_268),
.A2(n_11),
.B(n_10),
.Y(n_299)
);

OAI321xp33_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_10),
.A3(n_276),
.B1(n_272),
.B2(n_6),
.C(n_7),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_295),
.A2(n_281),
.B1(n_267),
.B2(n_275),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_301),
.B1(n_289),
.B2(n_308),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_312),
.B(n_299),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_278),
.B(n_273),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_304),
.A2(n_307),
.B(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_302),
.C(n_310),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_294),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_306),
.A2(n_290),
.B(n_289),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_4),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_3),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_287),
.A2(n_3),
.B(n_4),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_314),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_316),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_321),
.C(n_6),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_300),
.B(n_290),
.CI(n_5),
.CON(n_318),
.SN(n_318)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_303),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_290),
.Y(n_320)
);

AOI21xp33_ASAP7_75t_SL g324 ( 
.A1(n_320),
.A2(n_4),
.B(n_5),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_9),
.B1(n_5),
.B2(n_6),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_324),
.A2(n_315),
.B(n_318),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_8),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_313),
.A2(n_8),
.B1(n_9),
.B2(n_317),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_322),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_8),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_9),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_330),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_332),
.B(n_333),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_329),
.C(n_325),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

NAND3xp33_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_323),
.C(n_335),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_339),
.B(n_323),
.CI(n_9),
.CON(n_340),
.SN(n_340)
);


endmodule