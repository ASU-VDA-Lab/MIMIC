module fake_jpeg_14563_n_303 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_33),
.B1(n_27),
.B2(n_16),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_33),
.B1(n_16),
.B2(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_27),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_49),
.Y(n_58)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_61),
.Y(n_86)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_68),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_24),
.B(n_17),
.C(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_65),
.Y(n_97)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_72),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_38),
.B1(n_32),
.B2(n_16),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_77),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_19),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_37),
.Y(n_77)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_17),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_20),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_93),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_39),
.B1(n_53),
.B2(n_47),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_39),
.B1(n_53),
.B2(n_47),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_33),
.B1(n_43),
.B2(n_15),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_38),
.B1(n_32),
.B2(n_31),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_48),
.B(n_22),
.C(n_20),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_26),
.B(n_29),
.Y(n_112)
);

NAND2x1_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_41),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_79),
.B(n_35),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_74),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_103),
.B1(n_26),
.B2(n_29),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_102),
.B(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_32),
.B1(n_38),
.B2(n_31),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_76),
.B1(n_63),
.B2(n_55),
.Y(n_122)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_66),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_111),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_110),
.B(n_28),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_86),
.B(n_64),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_126),
.B(n_25),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_115),
.B(n_118),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_36),
.C(n_73),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_85),
.C(n_82),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_103),
.B1(n_76),
.B2(n_112),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_63),
.B1(n_80),
.B2(n_84),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_125),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_23),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_61),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_96),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_18),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_92),
.C(n_103),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_143),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_132),
.B(n_111),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_147),
.B1(n_149),
.B2(n_42),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_137),
.B(n_151),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_144),
.C(n_154),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_97),
.B1(n_81),
.B2(n_105),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_0),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_104),
.A3(n_97),
.B1(n_101),
.B2(n_98),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_101),
.B1(n_67),
.B2(n_68),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_116),
.B1(n_108),
.B2(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_91),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_36),
.C(n_95),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_91),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_119),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_164),
.B1(n_109),
.B2(n_131),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_122),
.A2(n_121),
.B1(n_124),
.B2(n_126),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_28),
.B1(n_18),
.B2(n_54),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_36),
.B(n_23),
.C(n_21),
.D(n_28),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_73),
.A3(n_21),
.B1(n_28),
.B2(n_23),
.C1(n_14),
.C2(n_18),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_109),
.A2(n_69),
.B1(n_42),
.B2(n_35),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_165),
.A2(n_167),
.B1(n_145),
.B2(n_150),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_166),
.B(n_184),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_25),
.B1(n_113),
.B2(n_119),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_154),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_177),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_188),
.B1(n_159),
.B2(n_145),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_175),
.B(n_186),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_10),
.Y(n_177)
);

NAND2x1_ASAP7_75t_SL g178 ( 
.A(n_153),
.B(n_113),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_141),
.B(n_163),
.Y(n_197)
);

OA22x2_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_42),
.B1(n_99),
.B2(n_54),
.Y(n_179)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_13),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_185),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_13),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_194),
.Y(n_204)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_12),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_190),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_12),
.Y(n_190)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_192),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_140),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_155),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_217),
.B1(n_164),
.B2(n_18),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_146),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_146),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_211),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_142),
.C(n_147),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_214),
.C(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_150),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_161),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_151),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_218),
.B(n_171),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_219),
.B(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_167),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_224),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_221),
.A2(n_228),
.B1(n_236),
.B2(n_237),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_210),
.A2(n_188),
.B1(n_183),
.B2(n_193),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_197),
.B1(n_215),
.B2(n_212),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_211),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_226),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_216),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_210),
.A2(n_196),
.B1(n_199),
.B2(n_201),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_177),
.C(n_165),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_235),
.C(n_215),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_181),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_178),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_198),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_179),
.C(n_189),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_179),
.B1(n_191),
.B2(n_185),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_243),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_225),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_240),
.A2(n_227),
.B1(n_236),
.B2(n_2),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_203),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_244),
.C(n_246),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_200),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_204),
.B1(n_197),
.B2(n_202),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_245),
.B(n_251),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_233),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_234),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_223),
.A2(n_212),
.B(n_12),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_11),
.B(n_10),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

HAxp5_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_231),
.CON(n_256),
.SN(n_256)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_246),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_261),
.C(n_262),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_18),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_54),
.C(n_18),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_249),
.C(n_243),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_239),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_264),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_238),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_255),
.C(n_257),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_272),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_0),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_0),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_274),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_0),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_4),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_255),
.C(n_261),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_283),
.C(n_268),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_287),
.Y(n_294)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_265),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_290),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_269),
.B1(n_5),
.B2(n_6),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_4),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_292),
.B(n_281),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_4),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_280),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_294),
.A2(n_287),
.B(n_288),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_296),
.A2(n_297),
.B1(n_295),
.B2(n_6),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_5),
.C(n_6),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_5),
.B(n_6),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_300),
.B(n_5),
.Y(n_301)
);

AOI221xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_7),
.B1(n_8),
.B2(n_295),
.C(n_287),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_7),
.Y(n_303)
);


endmodule