module fake_jpeg_1814_n_115 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_46),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_49),
.Y(n_52)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_40),
.B1(n_41),
.B2(n_32),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_56),
.B1(n_34),
.B2(n_37),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_58),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_45),
.B1(n_43),
.B2(n_32),
.Y(n_56)
);

OR2x4_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_63),
.Y(n_77)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_68),
.Y(n_75)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_33),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_37),
.B(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_82),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_36),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_81),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_54),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_84),
.B1(n_5),
.B2(n_6),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_83),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_16),
.C(n_31),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_14),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_61),
.B1(n_2),
.B2(n_4),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_87),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_1),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_94),
.B(n_12),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_96),
.B1(n_12),
.B2(n_18),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_5),
.B(n_6),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_7),
.B(n_8),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_9),
.B(n_10),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_73),
.B1(n_10),
.B2(n_11),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_97),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_100),
.C(n_101),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_23),
.C(n_17),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_104),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_86),
.C(n_94),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_95),
.C(n_99),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_102),
.B(n_88),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_110),
.B1(n_105),
.B2(n_96),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_108),
.C(n_98),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_98),
.B(n_27),
.Y(n_113)
);

AOI21x1_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_25),
.B(n_28),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_30),
.Y(n_115)
);


endmodule