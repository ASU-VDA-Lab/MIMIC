module real_aes_9356_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_360;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_559;
wire n_466;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_0), .A2(n_245), .B1(n_493), .B2(n_654), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_0), .A2(n_245), .B1(n_335), .B2(n_1039), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_1), .A2(n_21), .B1(n_489), .B2(n_500), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_1), .A2(n_263), .B1(n_313), .B2(n_547), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g1469 ( .A(n_2), .Y(n_1469) );
INVxp67_ASAP7_75t_SL g568 ( .A(n_3), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_3), .A2(n_26), .B1(n_594), .B2(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g904 ( .A(n_4), .Y(n_904) );
INVx1_ASAP7_75t_L g964 ( .A(n_5), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_6), .A2(n_68), .B1(n_1192), .B2(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g847 ( .A(n_7), .Y(n_847) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_8), .Y(n_295) );
INVx1_ASAP7_75t_L g447 ( .A(n_8), .Y(n_447) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_8), .B(n_316), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_8), .B(n_204), .Y(n_1434) );
INVxp67_ASAP7_75t_SL g1570 ( .A(n_9), .Y(n_1570) );
AOI22xp33_ASAP7_75t_L g1585 ( .A1(n_9), .A2(n_45), .B1(n_1586), .B2(n_1588), .Y(n_1585) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_10), .A2(n_105), .B1(n_763), .B2(n_872), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_10), .A2(n_105), .B1(n_1160), .B2(n_1161), .Y(n_1159) );
AOI22xp33_ASAP7_75t_SL g646 ( .A1(n_11), .A2(n_220), .B1(n_438), .B2(n_585), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_11), .A2(n_220), .B1(n_473), .B2(n_534), .Y(n_656) );
OAI221xp5_ASAP7_75t_SL g1412 ( .A1(n_12), .A2(n_59), .B1(n_1413), .B2(n_1418), .C(n_1420), .Y(n_1412) );
AOI221xp5_ASAP7_75t_L g1472 ( .A1(n_12), .A2(n_125), .B1(n_1473), .B2(n_1475), .C(n_1477), .Y(n_1472) );
INVx1_ASAP7_75t_L g1454 ( .A(n_13), .Y(n_1454) );
AOI221xp5_ASAP7_75t_SL g799 ( .A1(n_14), .A2(n_39), .B1(n_800), .B2(n_801), .C(n_802), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_14), .A2(n_39), .B1(n_822), .B2(n_823), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_15), .A2(n_188), .B1(n_438), .B2(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_15), .A2(n_188), .B1(n_534), .B2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_16), .A2(n_271), .B1(n_473), .B2(n_534), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_16), .A2(n_271), .B1(n_543), .B2(n_547), .Y(n_542) );
AO22x2_ASAP7_75t_L g951 ( .A1(n_17), .A2(n_952), .B1(n_1007), .B2(n_1008), .Y(n_951) );
INVx1_ASAP7_75t_L g1007 ( .A(n_17), .Y(n_1007) );
CKINVDCx5p33_ASAP7_75t_R g712 ( .A(n_18), .Y(n_712) );
INVx1_ASAP7_75t_L g1453 ( .A(n_19), .Y(n_1453) );
INVx1_ASAP7_75t_L g558 ( .A(n_20), .Y(n_558) );
INVx1_ASAP7_75t_L g754 ( .A(n_21), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g1233 ( .A1(n_22), .A2(n_76), .B1(n_1188), .B2(n_1192), .Y(n_1233) );
INVx1_ASAP7_75t_L g1544 ( .A(n_23), .Y(n_1544) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_24), .A2(n_209), .B1(n_484), .B2(n_499), .Y(n_795) );
AOI221xp5_ASAP7_75t_L g807 ( .A1(n_24), .A2(n_209), .B1(n_414), .B2(n_808), .C(n_811), .Y(n_807) );
AOI22xp33_ASAP7_75t_SL g980 ( .A1(n_25), .A2(n_276), .B1(n_423), .B2(n_981), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_25), .A2(n_276), .B1(n_390), .B2(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g567 ( .A(n_26), .Y(n_567) );
INVx1_ASAP7_75t_L g621 ( .A(n_27), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_27), .A2(n_147), .B1(n_539), .B2(n_648), .Y(n_651) );
XNOR2xp5_ASAP7_75t_L g721 ( .A(n_28), .B(n_722), .Y(n_721) );
INVxp33_ASAP7_75t_L g346 ( .A(n_29), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_29), .A2(n_239), .B1(n_450), .B2(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g364 ( .A(n_30), .Y(n_364) );
OR2x2_ASAP7_75t_L g1485 ( .A(n_30), .B(n_1468), .Y(n_1485) );
INVx1_ASAP7_75t_L g553 ( .A(n_31), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g1232 ( .A1(n_31), .A2(n_148), .B1(n_1176), .B2(n_1184), .Y(n_1232) );
OAI221xp5_ASAP7_75t_L g1426 ( .A1(n_32), .A2(n_70), .B1(n_1427), .B2(n_1435), .C(n_1440), .Y(n_1426) );
OAI22xp5_ASAP7_75t_L g1486 ( .A1(n_32), .A2(n_70), .B1(n_1487), .B2(n_1491), .Y(n_1486) );
INVx1_ASAP7_75t_L g1127 ( .A(n_33), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_33), .A2(n_132), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
INVx1_ASAP7_75t_L g1069 ( .A(n_34), .Y(n_1069) );
AOI22xp33_ASAP7_75t_SL g1083 ( .A1(n_34), .A2(n_226), .B1(n_539), .B2(n_1084), .Y(n_1083) );
BUFx2_ASAP7_75t_L g357 ( .A(n_35), .Y(n_357) );
BUFx2_ASAP7_75t_L g410 ( .A(n_35), .Y(n_410) );
INVx1_ASAP7_75t_L g445 ( .A(n_35), .Y(n_445) );
OR2x2_ASAP7_75t_L g1433 ( .A(n_35), .B(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1120 ( .A(n_36), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_36), .A2(n_110), .B1(n_504), .B2(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1224 ( .A(n_37), .Y(n_1224) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_38), .A2(n_127), .B1(n_473), .B2(n_914), .Y(n_1036) );
INVxp67_ASAP7_75t_L g1047 ( .A(n_38), .Y(n_1047) );
INVx1_ASAP7_75t_L g1133 ( .A(n_40), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_40), .A2(n_47), .B1(n_872), .B2(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g765 ( .A(n_41), .Y(n_765) );
AO22x2_ASAP7_75t_L g1110 ( .A1(n_42), .A2(n_1111), .B1(n_1112), .B2(n_1163), .Y(n_1110) );
INVx1_ASAP7_75t_L g1163 ( .A(n_42), .Y(n_1163) );
INVx1_ASAP7_75t_L g388 ( .A(n_43), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_43), .A2(n_158), .B1(n_422), .B2(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_SL g1444 ( .A(n_44), .Y(n_1444) );
AOI22xp33_ASAP7_75t_L g1502 ( .A1(n_44), .A2(n_171), .B1(n_871), .B2(n_1005), .Y(n_1502) );
INVxp67_ASAP7_75t_SL g1573 ( .A(n_45), .Y(n_1573) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_46), .A2(n_259), .B1(n_426), .B2(n_648), .Y(n_1574) );
AOI221xp5_ASAP7_75t_SL g1581 ( .A1(n_46), .A2(n_461), .B1(n_1582), .B2(n_1583), .C(n_1589), .Y(n_1581) );
INVx1_ASAP7_75t_L g1129 ( .A(n_47), .Y(n_1129) );
INVx1_ASAP7_75t_L g625 ( .A(n_48), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_48), .A2(n_255), .B1(n_416), .B2(n_438), .Y(n_650) );
OAI211xp5_ASAP7_75t_L g1542 ( .A1(n_49), .A2(n_494), .B(n_1106), .C(n_1543), .Y(n_1542) );
INVx1_ASAP7_75t_L g1563 ( .A(n_49), .Y(n_1563) );
INVx1_ASAP7_75t_L g557 ( .A(n_50), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_50), .A2(n_203), .B1(n_539), .B2(n_587), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_51), .A2(n_268), .B1(n_534), .B2(n_704), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_51), .A2(n_189), .B1(n_313), .B2(n_547), .Y(n_715) );
INVx1_ASAP7_75t_L g958 ( .A(n_52), .Y(n_958) );
INVx1_ASAP7_75t_L g939 ( .A(n_53), .Y(n_939) );
OAI211xp5_ASAP7_75t_L g943 ( .A1(n_53), .A2(n_494), .B(n_692), .C(n_944), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_54), .A2(n_117), .B1(n_1176), .B2(n_1184), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_55), .A2(n_159), .B1(n_422), .B2(n_426), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_55), .A2(n_159), .B1(n_450), .B2(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g785 ( .A(n_56), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_56), .A2(n_193), .B1(n_829), .B2(n_830), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_57), .Y(n_804) );
INVx1_ASAP7_75t_L g1119 ( .A(n_58), .Y(n_1119) );
AOI22xp33_ASAP7_75t_SL g1149 ( .A1(n_58), .A2(n_79), .B1(n_1150), .B2(n_1152), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1478 ( .A1(n_59), .A2(n_143), .B1(n_1479), .B2(n_1480), .Y(n_1478) );
CKINVDCx5p33_ASAP7_75t_R g1061 ( .A(n_60), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_61), .A2(n_66), .B1(n_865), .B2(n_866), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_61), .A2(n_66), .B1(n_414), .B2(n_800), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_62), .A2(n_246), .B1(n_452), .B2(n_878), .Y(n_1035) );
INVxp33_ASAP7_75t_L g1049 ( .A(n_62), .Y(n_1049) );
INVxp33_ASAP7_75t_SL g1445 ( .A(n_63), .Y(n_1445) );
AOI221xp5_ASAP7_75t_L g1495 ( .A1(n_63), .A2(n_229), .B1(n_1496), .B2(n_1497), .C(n_1500), .Y(n_1495) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_64), .A2(n_90), .B1(n_484), .B2(n_489), .Y(n_483) );
INVx1_ASAP7_75t_L g516 ( .A(n_64), .Y(n_516) );
INVx1_ASAP7_75t_L g685 ( .A(n_65), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_65), .A2(n_189), .B1(n_484), .B2(n_489), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g498 ( .A1(n_67), .A2(n_258), .B1(n_499), .B2(n_500), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_67), .A2(n_258), .B1(n_414), .B2(n_436), .C(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_69), .A2(n_891), .B1(n_946), .B2(n_947), .Y(n_890) );
INVx1_ASAP7_75t_L g947 ( .A(n_69), .Y(n_947) );
INVx1_ASAP7_75t_L g764 ( .A(n_71), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_72), .A2(n_131), .B1(n_1176), .B2(n_1184), .Y(n_1206) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_73), .A2(n_77), .B1(n_543), .B2(n_547), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_73), .A2(n_77), .B1(n_704), .B2(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g735 ( .A(n_74), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_75), .A2(n_248), .B1(n_414), .B2(n_417), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_75), .A2(n_248), .B1(n_455), .B2(n_458), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g1079 ( .A1(n_78), .A2(n_278), .B1(n_438), .B2(n_585), .Y(n_1079) );
AOI22xp33_ASAP7_75t_SL g1087 ( .A1(n_78), .A2(n_278), .B1(n_696), .B2(n_1088), .Y(n_1087) );
OAI222xp33_ASAP7_75t_L g1115 ( .A1(n_79), .A2(n_174), .B1(n_265), .B2(n_562), .C1(n_565), .C2(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g339 ( .A(n_80), .Y(n_339) );
INVx1_ASAP7_75t_L g643 ( .A(n_81), .Y(n_643) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_81), .A2(n_91), .B1(n_473), .B2(n_474), .Y(n_659) );
INVx1_ASAP7_75t_L g681 ( .A(n_82), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_82), .A2(n_180), .B1(n_499), .B2(n_500), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_83), .A2(n_167), .B1(n_539), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_83), .A2(n_167), .B1(n_493), .B2(n_654), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_84), .A2(n_115), .B1(n_565), .B2(n_630), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_84), .A2(n_115), .B1(n_574), .B2(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g577 ( .A(n_85), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_85), .A2(n_108), .B1(n_473), .B2(n_474), .Y(n_614) );
INVx1_ASAP7_75t_L g740 ( .A(n_86), .Y(n_740) );
OAI211xp5_ASAP7_75t_SL g768 ( .A1(n_86), .A2(n_352), .B(n_717), .C(n_769), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_87), .Y(n_781) );
INVxp33_ASAP7_75t_SL g854 ( .A(n_88), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_88), .A2(n_257), .B1(n_335), .B2(n_505), .Y(n_883) );
INVxp67_ASAP7_75t_SL g959 ( .A(n_89), .Y(n_959) );
AOI22xp33_ASAP7_75t_SL g983 ( .A1(n_89), .A2(n_212), .B1(n_504), .B2(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g541 ( .A(n_90), .Y(n_541) );
INVx1_ASAP7_75t_L g641 ( .A(n_91), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_92), .A2(n_193), .B1(n_543), .B2(n_547), .Y(n_778) );
INVx1_ASAP7_75t_L g827 ( .A(n_92), .Y(n_827) );
INVx1_ASAP7_75t_L g1022 ( .A(n_93), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_93), .A2(n_101), .B1(n_573), .B2(n_1044), .Y(n_1043) );
AO22x2_ASAP7_75t_L g1053 ( .A1(n_94), .A2(n_1054), .B1(n_1094), .B2(n_1095), .Y(n_1053) );
INVxp67_ASAP7_75t_L g1094 ( .A(n_94), .Y(n_1094) );
INVx1_ASAP7_75t_L g408 ( .A(n_95), .Y(n_408) );
INVx1_ASAP7_75t_L g1468 ( .A(n_95), .Y(n_1468) );
INVx1_ASAP7_75t_L g905 ( .A(n_96), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_97), .A2(n_175), .B1(n_871), .B2(n_874), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_97), .A2(n_175), .B1(n_808), .B2(n_843), .Y(n_880) );
INVx1_ASAP7_75t_L g961 ( .A(n_98), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_98), .A2(n_192), .B1(n_981), .B2(n_987), .Y(n_986) );
INVxp33_ASAP7_75t_SL g968 ( .A(n_99), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_99), .A2(n_202), .B1(n_1004), .B2(n_1005), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_100), .A2(n_145), .B1(n_504), .B2(n_978), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_100), .A2(n_145), .B1(n_995), .B2(n_997), .Y(n_994) );
INVx1_ASAP7_75t_L g1024 ( .A(n_101), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g1221 ( .A(n_102), .Y(n_1221) );
INVx1_ASAP7_75t_L g702 ( .A(n_103), .Y(n_702) );
OAI211xp5_ASAP7_75t_SL g716 ( .A1(n_103), .A2(n_352), .B(n_717), .C(n_719), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g1551 ( .A1(n_104), .A2(n_179), .B1(n_296), .B2(n_313), .Y(n_1551) );
INVx1_ASAP7_75t_L g1576 ( .A(n_104), .Y(n_1576) );
INVx1_ASAP7_75t_L g507 ( .A(n_106), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_107), .A2(n_197), .B1(n_562), .B2(n_565), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_107), .A2(n_197), .B1(n_573), .B2(n_574), .Y(n_572) );
INVxp67_ASAP7_75t_L g580 ( .A(n_108), .Y(n_580) );
INVx1_ASAP7_75t_L g729 ( .A(n_109), .Y(n_729) );
INVx1_ASAP7_75t_L g1123 ( .A(n_110), .Y(n_1123) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_111), .A2(n_134), .B1(n_1176), .B2(n_1184), .Y(n_1202) );
INVx1_ASAP7_75t_L g757 ( .A(n_112), .Y(n_757) );
INVx1_ASAP7_75t_L g938 ( .A(n_113), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_113), .A2(n_164), .B1(n_484), .B2(n_499), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_114), .A2(n_217), .B1(n_1176), .B2(n_1184), .Y(n_1195) );
INVx1_ASAP7_75t_L g1057 ( .A(n_116), .Y(n_1057) );
AOI22xp33_ASAP7_75t_SL g1093 ( .A1(n_116), .A2(n_240), .B1(n_473), .B2(n_474), .Y(n_1093) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_118), .A2(n_149), .B1(n_1188), .B2(n_1192), .Y(n_1187) );
XOR2xp5_ASAP7_75t_L g1535 ( .A(n_119), .B(n_1536), .Y(n_1535) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_120), .A2(n_153), .B1(n_1004), .B2(n_1140), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_120), .A2(n_153), .B1(n_1154), .B2(n_1156), .Y(n_1153) );
INVx1_ASAP7_75t_L g1212 ( .A(n_121), .Y(n_1212) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_122), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_122), .A2(n_196), .B1(n_534), .B2(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_123), .A2(n_215), .B1(n_590), .B2(n_1039), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_123), .A2(n_215), .B1(n_478), .B2(n_613), .Y(n_1086) );
INVxp33_ASAP7_75t_SL g839 ( .A(n_124), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_124), .A2(n_256), .B1(n_865), .B2(n_877), .Y(n_876) );
INVxp33_ASAP7_75t_SL g1423 ( .A(n_125), .Y(n_1423) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_126), .A2(n_166), .B1(n_866), .B2(n_907), .Y(n_906) );
INVxp67_ASAP7_75t_SL g921 ( .A(n_126), .Y(n_921) );
INVxp33_ASAP7_75t_L g1046 ( .A(n_127), .Y(n_1046) );
OAI211xp5_ASAP7_75t_L g1549 ( .A1(n_128), .A2(n_352), .B(n_1099), .C(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1577 ( .A(n_128), .Y(n_1577) );
INVx1_ASAP7_75t_L g739 ( .A(n_129), .Y(n_739) );
OAI22xp33_ASAP7_75t_SL g770 ( .A1(n_129), .A2(n_162), .B1(n_296), .B2(n_543), .Y(n_770) );
AO22x2_ASAP7_75t_L g1012 ( .A1(n_130), .A2(n_1013), .B1(n_1050), .B2(n_1051), .Y(n_1012) );
INVx1_ASAP7_75t_L g1050 ( .A(n_130), .Y(n_1050) );
INVx1_ASAP7_75t_L g1126 ( .A(n_132), .Y(n_1126) );
INVx1_ASAP7_75t_L g287 ( .A(n_133), .Y(n_287) );
INVx1_ASAP7_75t_L g640 ( .A(n_135), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_135), .A2(n_213), .B1(n_478), .B2(n_654), .Y(n_658) );
AO22x1_ASAP7_75t_SL g1209 ( .A1(n_136), .A2(n_227), .B1(n_1176), .B2(n_1184), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1546 ( .A1(n_137), .A2(n_187), .B1(n_484), .B2(n_499), .Y(n_1546) );
INVx1_ASAP7_75t_L g1555 ( .A(n_137), .Y(n_1555) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_138), .A2(n_216), .B1(n_504), .B2(n_505), .C(n_506), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_138), .A2(n_216), .B1(n_473), .B2(n_474), .Y(n_529) );
INVx1_ASAP7_75t_L g497 ( .A(n_139), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g894 ( .A1(n_140), .A2(n_352), .B(n_895), .C(n_896), .Y(n_894) );
INVx1_ASAP7_75t_L g912 ( .A(n_140), .Y(n_912) );
AO221x2_ASAP7_75t_L g1218 ( .A1(n_141), .A2(n_266), .B1(n_1204), .B2(n_1219), .C(n_1220), .Y(n_1218) );
INVx1_ASAP7_75t_L g1280 ( .A(n_142), .Y(n_1280) );
INVxp33_ASAP7_75t_SL g1421 ( .A(n_143), .Y(n_1421) );
CKINVDCx5p33_ASAP7_75t_R g1066 ( .A(n_144), .Y(n_1066) );
INVx1_ASAP7_75t_L g1026 ( .A(n_146), .Y(n_1026) );
INVx1_ASAP7_75t_L g628 ( .A(n_147), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_150), .A2(n_156), .B1(n_457), .B2(n_474), .Y(n_1030) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_150), .A2(n_156), .B1(n_438), .B2(n_585), .Y(n_1037) );
INVx1_ASAP7_75t_L g308 ( .A(n_151), .Y(n_308) );
CKINVDCx14_ASAP7_75t_R g480 ( .A(n_152), .Y(n_480) );
XOR2xp5_ASAP7_75t_L g661 ( .A(n_154), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g496 ( .A(n_155), .Y(n_496) );
INVxp33_ASAP7_75t_SL g1016 ( .A(n_157), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_157), .A2(n_169), .B1(n_335), .B2(n_648), .Y(n_1033) );
INVxp33_ASAP7_75t_L g360 ( .A(n_158), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g1196 ( .A1(n_160), .A2(n_262), .B1(n_1188), .B2(n_1192), .Y(n_1196) );
INVx1_ASAP7_75t_L g732 ( .A(n_161), .Y(n_732) );
INVx1_ASAP7_75t_L g742 ( .A(n_162), .Y(n_742) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_163), .Y(n_782) );
INVx1_ASAP7_75t_L g930 ( .A(n_164), .Y(n_930) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_165), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_165), .A2(n_210), .B1(n_435), .B2(n_436), .Y(n_434) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_166), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g803 ( .A(n_168), .Y(n_803) );
INVxp67_ASAP7_75t_SL g1019 ( .A(n_169), .Y(n_1019) );
INVxp33_ASAP7_75t_SL g1027 ( .A(n_170), .Y(n_1027) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_170), .A2(n_184), .B1(n_438), .B2(n_585), .Y(n_1032) );
INVxp67_ASAP7_75t_SL g1450 ( .A(n_171), .Y(n_1450) );
INVx1_ASAP7_75t_L g753 ( .A(n_172), .Y(n_753) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_172), .A2(n_183), .B1(n_484), .B2(n_499), .Y(n_759) );
INVx1_ASAP7_75t_L g672 ( .A(n_173), .Y(n_672) );
INVx1_ASAP7_75t_L g1130 ( .A(n_174), .Y(n_1130) );
INVx1_ASAP7_75t_L g317 ( .A(n_176), .Y(n_317) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_177), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_177), .B(n_287), .Y(n_1183) );
AND3x2_ASAP7_75t_L g1189 ( .A(n_177), .B(n_287), .C(n_1180), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_178), .A2(n_250), .B1(n_1192), .B2(n_1204), .Y(n_1207) );
OAI22xp33_ASAP7_75t_L g1541 ( .A1(n_179), .A2(n_235), .B1(n_489), .B2(n_500), .Y(n_1541) );
INVx1_ASAP7_75t_L g683 ( .A(n_180), .Y(n_683) );
INVx2_ASAP7_75t_L g300 ( .A(n_181), .Y(n_300) );
INVx1_ASAP7_75t_L g1456 ( .A(n_182), .Y(n_1456) );
INVx1_ASAP7_75t_L g756 ( .A(n_183), .Y(n_756) );
INVxp33_ASAP7_75t_SL g1017 ( .A(n_184), .Y(n_1017) );
INVx1_ASAP7_75t_L g899 ( .A(n_185), .Y(n_899) );
INVx1_ASAP7_75t_L g1214 ( .A(n_186), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1524 ( .A1(n_186), .A2(n_1525), .B1(n_1533), .B2(n_1534), .Y(n_1524) );
INVx1_ASAP7_75t_L g1562 ( .A(n_187), .Y(n_1562) );
INVx1_ASAP7_75t_L g1180 ( .A(n_190), .Y(n_1180) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_191), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_191), .A2(n_234), .B1(n_471), .B2(n_474), .Y(n_470) );
INVxp33_ASAP7_75t_SL g955 ( .A(n_192), .Y(n_955) );
INVx1_ASAP7_75t_L g1075 ( .A(n_194), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_194), .A2(n_247), .B1(n_594), .B2(n_927), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1548 ( .A1(n_195), .A2(n_269), .B1(n_543), .B2(n_547), .Y(n_1548) );
AOI22xp33_ASAP7_75t_L g1578 ( .A1(n_195), .A2(n_269), .B1(n_1496), .B2(n_1579), .Y(n_1578) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_196), .Y(n_674) );
INVx1_ASAP7_75t_L g669 ( .A(n_198), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_199), .Y(n_623) );
INVx1_ASAP7_75t_L g531 ( .A(n_200), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_201), .A2(n_280), .B1(n_296), .B2(n_313), .Y(n_893) );
INVx1_ASAP7_75t_L g910 ( .A(n_201), .Y(n_910) );
INVxp33_ASAP7_75t_SL g969 ( .A(n_202), .Y(n_969) );
INVx1_ASAP7_75t_L g560 ( .A(n_203), .Y(n_560) );
INVx1_ASAP7_75t_L g302 ( .A(n_204), .Y(n_302) );
INVx2_ASAP7_75t_L g316 ( .A(n_204), .Y(n_316) );
OAI211xp5_ASAP7_75t_L g490 ( .A1(n_205), .A2(n_491), .B(n_494), .C(n_495), .Y(n_490) );
INVx1_ASAP7_75t_L g519 ( .A(n_205), .Y(n_519) );
INVx1_ASAP7_75t_L g571 ( .A(n_206), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_206), .A2(n_267), .B1(n_478), .B2(n_613), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_207), .A2(n_243), .B1(n_587), .B2(n_590), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_207), .A2(n_243), .B1(n_602), .B2(n_603), .Y(n_601) );
XNOR2xp5_ASAP7_75t_L g617 ( .A(n_208), .B(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_210), .Y(n_382) );
INVxp67_ASAP7_75t_SL g860 ( .A(n_211), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_211), .A2(n_260), .B1(n_414), .B2(n_808), .Y(n_882) );
INVxp33_ASAP7_75t_SL g956 ( .A(n_212), .Y(n_956) );
INVx1_ASAP7_75t_L g633 ( .A(n_213), .Y(n_633) );
INVx1_ASAP7_75t_L g1060 ( .A(n_214), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_214), .A2(n_277), .B1(n_603), .B2(n_1092), .Y(n_1091) );
OAI211xp5_ASAP7_75t_L g1098 ( .A1(n_214), .A2(n_352), .B(n_1099), .C(n_1101), .Y(n_1098) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_218), .Y(n_325) );
INVx1_ASAP7_75t_L g509 ( .A(n_219), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g1122 ( .A(n_221), .Y(n_1122) );
AOI221xp5_ASAP7_75t_L g1276 ( .A1(n_222), .A2(n_223), .B1(n_1277), .B2(n_1278), .C(n_1279), .Y(n_1276) );
OAI211xp5_ASAP7_75t_L g789 ( .A1(n_224), .A2(n_494), .B(n_790), .C(n_792), .Y(n_789) );
INVx1_ASAP7_75t_L g814 ( .A(n_224), .Y(n_814) );
INVx1_ASAP7_75t_L g850 ( .A(n_225), .Y(n_850) );
INVx1_ASAP7_75t_L g1073 ( .A(n_226), .Y(n_1073) );
OAI211xp5_ASAP7_75t_L g1105 ( .A1(n_226), .A2(n_494), .B(n_1106), .C(n_1108), .Y(n_1105) );
INVx1_ASAP7_75t_L g1545 ( .A(n_228), .Y(n_1545) );
INVxp67_ASAP7_75t_SL g1447 ( .A(n_229), .Y(n_1447) );
INVx1_ASAP7_75t_L g1457 ( .A(n_230), .Y(n_1457) );
INVx1_ASAP7_75t_L g699 ( .A(n_231), .Y(n_699) );
OAI22xp33_ASAP7_75t_SL g720 ( .A1(n_231), .A2(n_268), .B1(n_296), .B2(n_543), .Y(n_720) );
INVx1_ASAP7_75t_L g842 ( .A(n_232), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_232), .A2(n_252), .B1(n_389), .B2(n_866), .Y(n_875) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_233), .Y(n_783) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_234), .Y(n_351) );
INVx1_ASAP7_75t_L g1558 ( .A(n_235), .Y(n_1558) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_236), .A2(n_253), .B1(n_489), .B2(n_500), .Y(n_794) );
INVx1_ASAP7_75t_L g812 ( .A(n_236), .Y(n_812) );
AO22x2_ASAP7_75t_L g834 ( .A1(n_237), .A2(n_835), .B1(n_836), .B2(n_884), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_237), .Y(n_835) );
INVx1_ASAP7_75t_L g897 ( .A(n_238), .Y(n_897) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_239), .Y(n_333) );
INVx1_ASAP7_75t_L g1058 ( .A(n_240), .Y(n_1058) );
INVx1_ASAP7_75t_L g1181 ( .A(n_241), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_241), .B(n_1179), .Y(n_1186) );
INVx1_ASAP7_75t_L g726 ( .A(n_242), .Y(n_726) );
INVx1_ASAP7_75t_L g965 ( .A(n_244), .Y(n_965) );
INVxp67_ASAP7_75t_SL g1042 ( .A(n_246), .Y(n_1042) );
INVx1_ASAP7_75t_L g1070 ( .A(n_247), .Y(n_1070) );
AO22x2_ASAP7_75t_L g774 ( .A1(n_249), .A2(n_775), .B1(n_776), .B2(n_832), .Y(n_774) );
INVxp67_ASAP7_75t_L g832 ( .A(n_249), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_251), .Y(n_1062) );
INVxp67_ASAP7_75t_SL g840 ( .A(n_252), .Y(n_840) );
INVx1_ASAP7_75t_L g786 ( .A(n_253), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_254), .Y(n_711) );
INVx1_ASAP7_75t_L g626 ( .A(n_255), .Y(n_626) );
INVxp33_ASAP7_75t_SL g849 ( .A(n_256), .Y(n_849) );
INVx1_ASAP7_75t_L g856 ( .A(n_257), .Y(n_856) );
INVxp67_ASAP7_75t_SL g1584 ( .A(n_259), .Y(n_1584) );
INVxp33_ASAP7_75t_SL g858 ( .A(n_260), .Y(n_858) );
INVx2_ASAP7_75t_L g299 ( .A(n_261), .Y(n_299) );
INVx1_ASAP7_75t_L g744 ( .A(n_263), .Y(n_744) );
INVxp33_ASAP7_75t_SL g974 ( .A(n_264), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_264), .A2(n_281), .B1(n_1000), .B2(n_1002), .Y(n_999) );
INVx1_ASAP7_75t_L g1131 ( .A(n_265), .Y(n_1131) );
INVxp33_ASAP7_75t_L g576 ( .A(n_267), .Y(n_576) );
INVx1_ASAP7_75t_L g846 ( .A(n_270), .Y(n_846) );
BUFx3_ASAP7_75t_L g369 ( .A(n_272), .Y(n_369) );
INVx1_ASAP7_75t_L g386 ( .A(n_272), .Y(n_386) );
BUFx3_ASAP7_75t_L g371 ( .A(n_273), .Y(n_371) );
INVx1_ASAP7_75t_L g377 ( .A(n_273), .Y(n_377) );
INVx1_ASAP7_75t_L g932 ( .A(n_274), .Y(n_932) );
OAI22xp33_ASAP7_75t_L g945 ( .A1(n_274), .A2(n_280), .B1(n_489), .B2(n_500), .Y(n_945) );
INVx1_ASAP7_75t_L g532 ( .A(n_275), .Y(n_532) );
INVx1_ASAP7_75t_L g1065 ( .A(n_277), .Y(n_1065) );
INVx1_ASAP7_75t_L g687 ( .A(n_279), .Y(n_687) );
INVx1_ASAP7_75t_L g971 ( .A(n_281), .Y(n_971) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_303), .B(n_1168), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
AND2x4_ASAP7_75t_L g1523 ( .A(n_285), .B(n_291), .Y(n_1523) );
NOR2xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_SL g1531 ( .A(n_286), .Y(n_1531) );
NAND2xp5_ASAP7_75t_L g1532 ( .A(n_286), .B(n_288), .Y(n_1532) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_288), .B(n_1531), .Y(n_1533) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x6_ASAP7_75t_L g356 ( .A(n_293), .B(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g581 ( .A(n_293), .B(n_357), .Y(n_581) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g432 ( .A(n_294), .B(n_302), .Y(n_432) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g666 ( .A(n_295), .B(n_315), .Y(n_666) );
INVx8_ASAP7_75t_L g345 ( .A(n_296), .Y(n_345) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
OR2x6_ASAP7_75t_L g313 ( .A(n_297), .B(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_297), .Y(n_508) );
INVx2_ASAP7_75t_SL g518 ( .A(n_297), .Y(n_518) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_297), .Y(n_668) );
INVx2_ASAP7_75t_SL g749 ( .A(n_297), .Y(n_749) );
INVx1_ASAP7_75t_L g937 ( .A(n_297), .Y(n_937) );
OR2x2_ASAP7_75t_L g1462 ( .A(n_297), .B(n_1433), .Y(n_1462) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx2_ASAP7_75t_L g320 ( .A(n_299), .Y(n_320) );
INVx1_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
INVx1_ASAP7_75t_L g337 ( .A(n_299), .Y(n_337) );
AND2x4_ASAP7_75t_L g350 ( .A(n_299), .B(n_338), .Y(n_350) );
AND2x2_ASAP7_75t_L g425 ( .A(n_299), .B(n_300), .Y(n_425) );
INVx1_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
INVx2_ASAP7_75t_L g338 ( .A(n_300), .Y(n_338) );
INVx1_ASAP7_75t_L g343 ( .A(n_300), .Y(n_343) );
INVx1_ASAP7_75t_L g512 ( .A(n_300), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_300), .B(n_320), .Y(n_546) );
AND2x4_ASAP7_75t_L g342 ( .A(n_301), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g574 ( .A(n_302), .B(n_328), .Y(n_574) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_302), .B(n_328), .Y(n_1044) );
OAI22xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_886), .B1(n_1166), .B2(n_1167), .Y(n_303) );
INVx1_ASAP7_75t_L g1166 ( .A(n_304), .Y(n_1166) );
XOR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_773), .Y(n_304) );
XNOR2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_549), .Y(n_305) );
XNOR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_479), .Y(n_306) );
XNOR2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_355), .B1(n_358), .B2(n_404), .C(n_411), .Y(n_309) );
NAND4xp25_ASAP7_75t_L g310 ( .A(n_311), .B(n_324), .C(n_344), .D(n_352), .Y(n_310) );
AOI22xp33_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_317), .B1(n_318), .B2(n_323), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_312), .A2(n_345), .B1(n_531), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_312), .A2(n_345), .B1(n_849), .B2(n_850), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g1064 ( .A1(n_312), .A2(n_345), .B1(n_1065), .B2(n_1066), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_312), .A2(n_345), .B1(n_1122), .B2(n_1133), .Y(n_1132) );
INVx4_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx5_ASAP7_75t_L g579 ( .A(n_313), .Y(n_579) );
AND2x4_ASAP7_75t_L g318 ( .A(n_314), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g347 ( .A(n_314), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g544 ( .A(n_314), .Y(n_544) );
AND2x4_ASAP7_75t_L g548 ( .A(n_314), .B(n_348), .Y(n_548) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g332 ( .A(n_316), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_317), .A2(n_379), .B1(n_382), .B2(n_383), .Y(n_378) );
AOI22xp33_ASAP7_75t_SL g575 ( .A1(n_318), .A2(n_345), .B1(n_576), .B2(n_577), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_318), .A2(n_345), .B1(n_640), .B2(n_641), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_318), .A2(n_548), .B1(n_839), .B2(n_840), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_318), .A2(n_347), .B1(n_968), .B2(n_969), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_318), .A2(n_347), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g1056 ( .A1(n_318), .A2(n_548), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_318), .A2(n_548), .B1(n_1126), .B2(n_1127), .Y(n_1125) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_319), .Y(n_416) );
BUFx2_ASAP7_75t_L g435 ( .A(n_319), .Y(n_435) );
BUFx2_ASAP7_75t_L g504 ( .A(n_319), .Y(n_504) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_319), .Y(n_585) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_319), .Y(n_594) );
INVx1_ASAP7_75t_L g1155 ( .A(n_319), .Y(n_1155) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g1439 ( .A(n_320), .Y(n_1439) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_333), .B2(n_334), .C1(n_339), .C2(n_340), .Y(n_324) );
AOI222xp33_ASAP7_75t_L g387 ( .A1(n_325), .A2(n_339), .B1(n_388), .B2(n_389), .C1(n_393), .C2(n_398), .Y(n_387) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_326), .A2(n_342), .B1(n_496), .B2(n_497), .C1(n_532), .C2(n_538), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_326), .A2(n_342), .B1(n_711), .B2(n_712), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_326), .A2(n_342), .B1(n_764), .B2(n_765), .Y(n_769) );
AOI222xp33_ASAP7_75t_L g780 ( .A1(n_326), .A2(n_335), .B1(n_342), .B2(n_781), .C1(n_782), .C2(n_783), .Y(n_780) );
AOI222xp33_ASAP7_75t_L g841 ( .A1(n_326), .A2(n_342), .B1(n_842), .B2(n_843), .C1(n_846), .C2(n_847), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_326), .A2(n_897), .B1(n_898), .B2(n_899), .Y(n_896) );
AOI222xp33_ASAP7_75t_L g970 ( .A1(n_326), .A2(n_340), .B1(n_964), .B2(n_965), .C1(n_971), .C2(n_972), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g1101 ( .A1(n_326), .A2(n_898), .B1(n_1061), .B2(n_1062), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1550 ( .A1(n_326), .A2(n_340), .B1(n_1544), .B2(n_1545), .Y(n_1550) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_330), .Y(n_326) );
AND2x4_ASAP7_75t_L g1063 ( .A(n_327), .B(n_330), .Y(n_1063) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g511 ( .A(n_329), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_329), .B(n_512), .Y(n_671) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g354 ( .A(n_331), .Y(n_354) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2x1p5_ASAP7_75t_L g446 ( .A(n_332), .B(n_447), .Y(n_446) );
AOI211xp5_ASAP7_75t_L g1041 ( .A1(n_334), .A2(n_353), .B(n_1042), .C(n_1043), .Y(n_1041) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_SL g441 ( .A(n_335), .Y(n_441) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g353 ( .A(n_336), .B(n_354), .Y(n_353) );
BUFx3_ASAP7_75t_L g427 ( .A(n_336), .Y(n_427) );
BUFx3_ASAP7_75t_L g539 ( .A(n_336), .Y(n_539) );
INVx1_ASAP7_75t_L g591 ( .A(n_336), .Y(n_591) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_336), .Y(n_636) );
BUFx2_ASAP7_75t_L g845 ( .A(n_336), .Y(n_845) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
AOI222xp33_ASAP7_75t_L g1059 ( .A1(n_340), .A2(n_426), .B1(n_1060), .B2(n_1061), .C1(n_1062), .C2(n_1063), .Y(n_1059) );
AOI222xp33_ASAP7_75t_L g1128 ( .A1(n_340), .A2(n_843), .B1(n_1063), .B2(n_1129), .C1(n_1130), .C2(n_1131), .Y(n_1128) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g573 ( .A(n_342), .Y(n_573) );
INVx2_ASAP7_75t_L g638 ( .A(n_342), .Y(n_638) );
INVx1_ASAP7_75t_L g1431 ( .A(n_343), .Y(n_1431) );
AOI22xp33_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_346), .B1(n_347), .B2(n_351), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_345), .A2(n_579), .B1(n_785), .B2(n_786), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_345), .A2(n_579), .B1(n_958), .B2(n_974), .Y(n_973) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_345), .A2(n_579), .B1(n_1026), .B2(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_349), .Y(n_596) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx3_ASAP7_75t_L g420 ( .A(n_350), .Y(n_420) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_350), .Y(n_438) );
INVx1_ASAP7_75t_L g1148 ( .A(n_350), .Y(n_1148) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_352), .B(n_537), .C(n_540), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g779 ( .A(n_352), .B(n_780), .C(n_784), .Y(n_779) );
NAND4xp25_ASAP7_75t_L g837 ( .A(n_352), .B(n_838), .C(n_841), .D(n_848), .Y(n_837) );
NAND4xp25_ASAP7_75t_SL g966 ( .A(n_352), .B(n_967), .C(n_970), .D(n_973), .Y(n_966) );
NAND4xp25_ASAP7_75t_L g1055 ( .A(n_352), .B(n_1056), .C(n_1059), .D(n_1064), .Y(n_1055) );
NAND4xp25_ASAP7_75t_SL g1124 ( .A(n_352), .B(n_1125), .C(n_1128), .D(n_1132), .Y(n_1124) );
CKINVDCx11_ASAP7_75t_R g352 ( .A(n_353), .Y(n_352) );
AOI211xp5_ASAP7_75t_L g570 ( .A1(n_353), .A2(n_538), .B(n_571), .C(n_572), .Y(n_570) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_353), .A2(n_633), .B(n_634), .C(n_637), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_355), .A2(n_536), .B(n_542), .Y(n_535) );
OAI31xp33_ASAP7_75t_SL g714 ( .A1(n_355), .A2(n_715), .A3(n_716), .B(n_720), .Y(n_714) );
OAI31xp33_ASAP7_75t_SL g766 ( .A1(n_355), .A2(n_767), .A3(n_768), .B(n_770), .Y(n_766) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_355), .A2(n_778), .B(n_779), .C(n_787), .Y(n_777) );
AOI221x1_ASAP7_75t_L g836 ( .A1(n_355), .A2(n_406), .B1(n_837), .B2(n_851), .C(n_861), .Y(n_836) );
OAI31xp33_ASAP7_75t_L g892 ( .A1(n_355), .A2(n_893), .A3(n_894), .B(n_900), .Y(n_892) );
AOI221x1_ASAP7_75t_L g952 ( .A1(n_355), .A2(n_797), .B1(n_953), .B2(n_966), .C(n_975), .Y(n_952) );
AOI221x1_ASAP7_75t_L g1054 ( .A1(n_355), .A2(n_797), .B1(n_1055), .B2(n_1067), .C(n_1076), .Y(n_1054) );
OAI31xp33_ASAP7_75t_L g1096 ( .A1(n_355), .A2(n_1097), .A3(n_1098), .B(n_1102), .Y(n_1096) );
AOI221x1_ASAP7_75t_L g1112 ( .A1(n_355), .A2(n_797), .B1(n_1113), .B2(n_1124), .C(n_1134), .Y(n_1112) );
OAI31xp33_ASAP7_75t_L g1547 ( .A1(n_355), .A2(n_1548), .A3(n_1549), .B(n_1551), .Y(n_1547) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g467 ( .A(n_357), .B(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g615 ( .A(n_357), .B(n_468), .Y(n_615) );
AND2x4_ASAP7_75t_L g1464 ( .A(n_357), .B(n_1465), .Y(n_1464) );
NAND4xp25_ASAP7_75t_L g358 ( .A(n_359), .B(n_378), .C(n_387), .D(n_400), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_372), .B2(n_373), .Y(n_359) );
AOI22xp5_ASAP7_75t_SL g556 ( .A1(n_361), .A2(n_379), .B1(n_557), .B2(n_558), .Y(n_556) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_361), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_361), .A2(n_373), .B1(n_955), .B2(n_956), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_361), .A2(n_373), .B1(n_1016), .B2(n_1017), .Y(n_1015) );
AND2x4_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .Y(n_361) );
AND2x6_ASAP7_75t_L g383 ( .A(n_362), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g622 ( .A(n_362), .B(n_365), .Y(n_622) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g563 ( .A(n_363), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g375 ( .A(n_364), .Y(n_375) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_364), .Y(n_381) );
AND2x2_ASAP7_75t_L g463 ( .A(n_364), .B(n_408), .Y(n_463) );
INVx2_ASAP7_75t_L g469 ( .A(n_364), .Y(n_469) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g451 ( .A(n_366), .Y(n_451) );
INVx1_ASAP7_75t_L g602 ( .A(n_366), .Y(n_602) );
INVx2_ASAP7_75t_L g873 ( .A(n_366), .Y(n_873) );
BUFx6f_ASAP7_75t_L g993 ( .A(n_366), .Y(n_993) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_366), .Y(n_1001) );
INVx6_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g379 ( .A(n_367), .B(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g613 ( .A(n_367), .Y(n_613) );
INVx2_ASAP7_75t_L g655 ( .A(n_367), .Y(n_655) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_367), .B(n_1466), .Y(n_1465) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx1_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g376 ( .A(n_369), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g392 ( .A(n_369), .B(n_371), .Y(n_392) );
INVx1_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g385 ( .A(n_371), .B(n_386), .Y(n_385) );
CKINVDCx6p67_ASAP7_75t_R g499 ( .A(n_373), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_373), .A2(n_383), .B1(n_567), .B2(n_568), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_373), .A2(n_383), .B1(n_625), .B2(n_626), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_373), .A2(n_858), .B1(n_859), .B2(n_860), .Y(n_857) );
AOI22xp5_ASAP7_75t_SL g1068 ( .A1(n_373), .A2(n_622), .B1(n_1069), .B2(n_1070), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_373), .A2(n_622), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
AND2x6_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g402 ( .A(n_374), .Y(n_402) );
INVx1_ASAP7_75t_L g485 ( .A(n_374), .Y(n_485) );
AND2x2_ASAP7_75t_L g492 ( .A(n_374), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x6_ASAP7_75t_L g398 ( .A(n_375), .B(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_376), .Y(n_457) );
BUFx3_ASAP7_75t_L g473 ( .A(n_376), .Y(n_473) );
INVx2_ASAP7_75t_SL g607 ( .A(n_376), .Y(n_607) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_376), .Y(n_696) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_376), .Y(n_704) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_376), .Y(n_728) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_376), .Y(n_1004) );
BUFx2_ASAP7_75t_L g1496 ( .A(n_376), .Y(n_1496) );
INVx1_ASAP7_75t_L g488 ( .A(n_377), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_379), .Y(n_489) );
AOI22xp5_ASAP7_75t_SL g620 ( .A1(n_379), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_379), .A2(n_383), .B1(n_850), .B2(n_854), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_379), .A2(n_383), .B1(n_958), .B2(n_959), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_379), .A2(n_383), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_379), .A2(n_383), .B1(n_1066), .B2(n_1075), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_379), .A2(n_383), .B1(n_1122), .B2(n_1123), .Y(n_1121) );
AND2x4_ASAP7_75t_L g394 ( .A(n_380), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_SL g1023 ( .A(n_380), .B(n_395), .Y(n_1023) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx4_ASAP7_75t_L g500 ( .A(n_383), .Y(n_500) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_384), .Y(n_474) );
INVx2_ASAP7_75t_L g743 ( .A(n_384), .Y(n_743) );
INVx1_ASAP7_75t_L g1580 ( .A(n_384), .Y(n_1580) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g459 ( .A(n_385), .Y(n_459) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_385), .Y(n_534) );
INVx2_ASAP7_75t_L g869 ( .A(n_385), .Y(n_869) );
INVx1_ASAP7_75t_L g1089 ( .A(n_385), .Y(n_1089) );
INVx1_ASAP7_75t_L g487 ( .A(n_386), .Y(n_487) );
AOI222xp33_ASAP7_75t_L g855 ( .A1(n_389), .A2(n_393), .B1(n_398), .B2(n_846), .C1(n_847), .C2(n_856), .Y(n_855) );
BUFx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx4f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_391), .Y(n_478) );
INVx2_ASAP7_75t_SL g710 ( .A(n_391), .Y(n_710) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_391), .Y(n_1002) );
INVx1_ASAP7_75t_L g1021 ( .A(n_391), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1505 ( .A(n_391), .B(n_1484), .Y(n_1505) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_392), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_393), .A2(n_398), .B1(n_781), .B2(n_783), .Y(n_792) );
AOI222xp33_ASAP7_75t_L g960 ( .A1(n_393), .A2(n_398), .B1(n_961), .B2(n_962), .C1(n_964), .C2(n_965), .Y(n_960) );
AOI222xp33_ASAP7_75t_L g1071 ( .A1(n_393), .A2(n_398), .B1(n_1061), .B2(n_1062), .C1(n_1072), .C2(n_1073), .Y(n_1071) );
BUFx4f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_394), .A2(n_398), .B1(n_496), .B2(n_497), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_394), .A2(n_398), .B1(n_897), .B2(n_899), .Y(n_944) );
AOI22xp33_ASAP7_75t_SL g1108 ( .A1(n_394), .A2(n_398), .B1(n_1061), .B2(n_1062), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1543 ( .A1(n_394), .A2(n_398), .B1(n_1544), .B2(n_1545), .Y(n_1543) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g564 ( .A(n_396), .Y(n_564) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g1490 ( .A(n_397), .Y(n_1490) );
INVx3_ASAP7_75t_L g565 ( .A(n_398), .Y(n_565) );
AOI222xp33_ASAP7_75t_L g708 ( .A1(n_398), .A2(n_563), .B1(n_687), .B2(n_709), .C1(n_711), .C2(n_712), .Y(n_708) );
AOI222xp33_ASAP7_75t_L g762 ( .A1(n_398), .A2(n_563), .B1(n_757), .B2(n_763), .C1(n_764), .C2(n_765), .Y(n_762) );
AOI222xp33_ASAP7_75t_L g1018 ( .A1(n_398), .A2(n_1019), .B1(n_1020), .B2(n_1022), .C1(n_1023), .C2(n_1024), .Y(n_1018) );
BUFx3_ASAP7_75t_L g1493 ( .A(n_399), .Y(n_1493) );
NAND4xp25_ASAP7_75t_L g555 ( .A(n_400), .B(n_556), .C(n_559), .D(n_566), .Y(n_555) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_400), .B(n_620), .C(n_624), .D(n_627), .Y(n_619) );
BUFx2_ASAP7_75t_L g852 ( .A(n_400), .Y(n_852) );
NAND4xp25_ASAP7_75t_L g1067 ( .A(n_400), .B(n_1068), .C(n_1071), .D(n_1074), .Y(n_1067) );
INVx5_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
CKINVDCx8_ASAP7_75t_R g494 ( .A(n_401), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g1114 ( .A(n_401), .B(n_1115), .Y(n_1114) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g453 ( .A(n_403), .Y(n_453) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_403), .Y(n_493) );
INVx1_ASAP7_75t_L g604 ( .A(n_403), .Y(n_604) );
BUFx6f_ASAP7_75t_L g1499 ( .A(n_403), .Y(n_1499) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_406), .Y(n_797) );
AND2x4_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
AND2x4_ASAP7_75t_L g501 ( .A(n_407), .B(n_409), .Y(n_501) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g468 ( .A(n_408), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g1518 ( .A(n_409), .Y(n_1518) );
BUFx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g431 ( .A(n_410), .Y(n_431) );
OR2x6_ASAP7_75t_L g665 ( .A(n_410), .B(n_666), .Y(n_665) );
NAND4xp25_ASAP7_75t_L g411 ( .A(n_412), .B(n_433), .C(n_448), .D(n_464), .Y(n_411) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_421), .C(n_428), .Y(n_412) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_416), .B(n_1416), .Y(n_1419) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g682 ( .A(n_419), .Y(n_682) );
BUFx3_ASAP7_75t_L g800 ( .A(n_419), .Y(n_800) );
AND2x4_ASAP7_75t_L g1422 ( .A(n_419), .B(n_1416), .Y(n_1422) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g679 ( .A(n_420), .Y(n_679) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_420), .Y(n_928) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g989 ( .A(n_424), .Y(n_989) );
INVx2_ASAP7_75t_SL g1151 ( .A(n_424), .Y(n_1151) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_425), .Y(n_589) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g1162 ( .A(n_427), .Y(n_1162) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_428), .A2(n_799), .B1(n_807), .B2(n_817), .C(n_819), .Y(n_798) );
AOI33xp33_ASAP7_75t_L g879 ( .A1(n_428), .A2(n_817), .A3(n_880), .B1(n_881), .B2(n_882), .B3(n_883), .Y(n_879) );
NAND3xp33_ASAP7_75t_L g976 ( .A(n_428), .B(n_977), .C(n_980), .Y(n_976) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g513 ( .A(n_430), .Y(n_513) );
NAND3xp33_ASAP7_75t_L g583 ( .A(n_430), .B(n_584), .C(n_586), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_430), .B(n_646), .C(n_647), .Y(n_645) );
AOI33xp33_ASAP7_75t_L g1034 ( .A1(n_430), .A2(n_615), .A3(n_1035), .B1(n_1036), .B2(n_1037), .B3(n_1038), .Y(n_1034) );
NAND3xp33_ASAP7_75t_L g1078 ( .A(n_430), .B(n_1079), .C(n_1080), .Y(n_1078) );
AOI33xp33_ASAP7_75t_L g1143 ( .A1(n_430), .A2(n_442), .A3(n_1144), .B1(n_1149), .B2(n_1153), .B3(n_1159), .Y(n_1143) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
OR2x6_ASAP7_75t_L g461 ( .A(n_431), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g522 ( .A(n_431), .B(n_462), .Y(n_522) );
AND2x2_ASAP7_75t_L g598 ( .A(n_431), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g609 ( .A(n_431), .B(n_610), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_439), .C(n_442), .Y(n_433) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_435), .Y(n_801) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g505 ( .A(n_438), .Y(n_505) );
INVx2_ASAP7_75t_SL g979 ( .A(n_438), .Y(n_979) );
INVx4_ASAP7_75t_L g985 ( .A(n_438), .Y(n_985) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
CKINVDCx8_ASAP7_75t_R g818 ( .A(n_442), .Y(n_818) );
NAND3xp33_ASAP7_75t_L g982 ( .A(n_442), .B(n_983), .C(n_986), .Y(n_982) );
INVx5_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx6_ASAP7_75t_L g520 ( .A(n_443), .Y(n_520) );
OR2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g1416 ( .A(n_445), .B(n_1417), .Y(n_1416) );
INVx2_ASAP7_75t_L g599 ( .A(n_446), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_454), .C(n_460), .Y(n_448) );
BUFx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_451), .Y(n_829) );
INVx1_ASAP7_75t_L g963 ( .A(n_452), .Y(n_963) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g763 ( .A(n_453), .Y(n_763) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_456), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g822 ( .A(n_457), .Y(n_822) );
AND2x4_ASAP7_75t_L g1483 ( .A(n_457), .B(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g1480 ( .A(n_459), .Y(n_1480) );
NAND3xp33_ASAP7_75t_L g990 ( .A(n_460), .B(n_991), .C(n_994), .Y(n_990) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_SL g819 ( .A1(n_461), .A2(n_466), .B1(n_820), .B2(n_824), .Y(n_819) );
INVx2_ASAP7_75t_L g863 ( .A(n_461), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_461), .A2(n_903), .B1(n_908), .B2(n_915), .Y(n_902) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g610 ( .A(n_463), .Y(n_610) );
BUFx3_ASAP7_75t_L g1501 ( .A(n_463), .Y(n_1501) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_470), .C(n_475), .Y(n_464) );
AOI33xp33_ASAP7_75t_L g862 ( .A1(n_465), .A2(n_863), .A3(n_864), .B1(n_870), .B2(n_875), .B3(n_876), .Y(n_862) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g521 ( .A1(n_466), .A2(n_522), .B1(n_523), .B2(n_530), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g689 ( .A1(n_466), .A2(n_609), .B1(n_690), .B2(n_697), .Y(n_689) );
INVx4_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx4f_ASAP7_75t_L g916 ( .A(n_467), .Y(n_916) );
BUFx4f_ASAP7_75t_L g1006 ( .A(n_467), .Y(n_1006) );
CKINVDCx5p33_ASAP7_75t_R g1477 ( .A(n_468), .Y(n_1477) );
AND2x4_ASAP7_75t_L g1466 ( .A(n_469), .B(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_478), .Y(n_874) );
XNOR2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
NAND3x1_ASAP7_75t_SL g481 ( .A(n_482), .B(n_502), .C(n_535), .Y(n_481) );
OAI31xp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_490), .A3(n_498), .B(n_501), .Y(n_482) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx2_ASAP7_75t_L g525 ( .A(n_486), .Y(n_525) );
INVx1_ASAP7_75t_L g734 ( .A(n_486), .Y(n_734) );
BUFx2_ASAP7_75t_L g909 ( .A(n_486), .Y(n_909) );
OR2x2_ASAP7_75t_L g1512 ( .A(n_486), .B(n_1485), .Y(n_1512) );
INVx1_ASAP7_75t_L g1590 ( .A(n_486), .Y(n_1590) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
AND2x2_ASAP7_75t_L g528 ( .A(n_487), .B(n_488), .Y(n_528) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_492), .A2(n_560), .B(n_561), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_492), .A2(n_628), .B(n_629), .Y(n_627) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_493), .Y(n_1072) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_494), .B(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_494), .B(n_762), .Y(n_761) );
NAND4xp25_ASAP7_75t_L g1014 ( .A(n_494), .B(n_1015), .C(n_1018), .D(n_1025), .Y(n_1014) );
AOI211xp5_ASAP7_75t_L g554 ( .A1(n_501), .A2(n_555), .B(n_569), .C(n_582), .Y(n_554) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_501), .A2(n_619), .B(n_631), .C(n_644), .Y(n_618) );
OAI31xp33_ASAP7_75t_SL g705 ( .A1(n_501), .A2(n_706), .A3(n_707), .B(n_713), .Y(n_705) );
OAI31xp33_ASAP7_75t_L g758 ( .A1(n_501), .A2(n_759), .A3(n_760), .B(n_761), .Y(n_758) );
OAI31xp33_ASAP7_75t_SL g941 ( .A1(n_501), .A2(n_942), .A3(n_943), .B(n_945), .Y(n_941) );
AOI211x1_ASAP7_75t_L g1013 ( .A1(n_501), .A2(n_1014), .B(n_1028), .C(n_1040), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_513), .B1(n_514), .B2(n_520), .C(n_521), .Y(n_502) );
INVx1_ASAP7_75t_L g813 ( .A(n_505), .Y(n_813) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_509), .B2(n_510), .Y(n_506) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_507), .A2(n_509), .B1(n_524), .B2(n_526), .C(n_529), .Y(n_523) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_508), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
OAI22xp33_ASAP7_75t_SL g515 ( .A1(n_510), .A2(n_516), .B1(n_517), .B2(n_519), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g755 ( .A1(n_510), .A2(n_748), .B1(n_756), .B2(n_757), .Y(n_755) );
BUFx2_ASAP7_75t_L g895 ( .A(n_510), .Y(n_895) );
INVx1_ASAP7_75t_L g1100 ( .A(n_510), .Y(n_1100) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g686 ( .A(n_511), .Y(n_686) );
BUFx2_ASAP7_75t_L g718 ( .A(n_511), .Y(n_718) );
OAI22xp5_ASAP7_75t_SL g802 ( .A1(n_517), .A2(n_803), .B1(n_804), .B2(n_805), .Y(n_802) );
OAI22xp33_ASAP7_75t_L g1443 ( .A1(n_517), .A2(n_816), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
OAI22xp33_ASAP7_75t_L g1455 ( .A1(n_517), .A2(n_816), .B1(n_1456), .B2(n_1457), .Y(n_1455) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g940 ( .A(n_520), .Y(n_940) );
INVx2_ASAP7_75t_L g1565 ( .A(n_520), .Y(n_1565) );
OAI33xp33_ASAP7_75t_L g724 ( .A1(n_522), .A2(n_725), .A3(n_731), .B1(n_738), .B2(n_741), .B3(n_745), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_524), .A2(n_526), .B1(n_531), .B2(n_532), .C(n_533), .Y(n_530) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_524), .A2(n_790), .B1(n_904), .B2(n_905), .C(n_906), .Y(n_903) );
OAI221xp5_ASAP7_75t_L g1575 ( .A1(n_524), .A2(n_790), .B1(n_1576), .B2(n_1577), .C(n_1578), .Y(n_1575) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g691 ( .A(n_525), .Y(n_691) );
INVx2_ASAP7_75t_L g698 ( .A(n_525), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g820 ( .A1(n_526), .A2(n_698), .B1(n_803), .B2(n_804), .C(n_821), .Y(n_820) );
OAI221xp5_ASAP7_75t_L g824 ( .A1(n_526), .A2(n_782), .B1(n_825), .B2(n_827), .C(n_828), .Y(n_824) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g791 ( .A(n_527), .Y(n_791) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g694 ( .A(n_528), .Y(n_694) );
BUFx2_ASAP7_75t_L g701 ( .A(n_528), .Y(n_701) );
BUFx4f_ASAP7_75t_L g737 ( .A(n_528), .Y(n_737) );
INVx1_ASAP7_75t_L g1107 ( .A(n_528), .Y(n_1107) );
INVx1_ASAP7_75t_L g730 ( .A(n_534), .Y(n_730) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_534), .Y(n_823) );
INVx1_ASAP7_75t_L g831 ( .A(n_534), .Y(n_831) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x6_ASAP7_75t_L g1425 ( .A(n_539), .B(n_1416), .Y(n_1425) );
NAND2x1p5_ASAP7_75t_L g1441 ( .A(n_539), .B(n_1432), .Y(n_1441) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g1569 ( .A(n_545), .Y(n_1569) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g676 ( .A(n_546), .Y(n_676) );
INVx1_ASAP7_75t_L g924 ( .A(n_546), .Y(n_924) );
INVx5_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_548), .A2(n_558), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_548), .A2(n_579), .B1(n_623), .B2(n_643), .Y(n_642) );
XOR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_660), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B1(n_616), .B2(n_617), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
XNOR2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g630 ( .A(n_563), .Y(n_630) );
AOI31xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_575), .A3(n_578), .B(n_581), .Y(n_569) );
AOI31xp33_ASAP7_75t_L g631 ( .A1(n_581), .A2(n_632), .A3(n_639), .B(n_642), .Y(n_631) );
AOI31xp33_ASAP7_75t_L g1040 ( .A1(n_581), .A2(n_1041), .A3(n_1045), .B(n_1048), .Y(n_1040) );
NAND4xp25_ASAP7_75t_L g582 ( .A(n_583), .B(n_592), .C(n_600), .D(n_611), .Y(n_582) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g648 ( .A(n_588), .Y(n_648) );
INVx2_ASAP7_75t_SL g1039 ( .A(n_588), .Y(n_1039) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx6f_ASAP7_75t_L g810 ( .A(n_589), .Y(n_810) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_589), .Y(n_1084) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_597), .C(n_598), .Y(n_592) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_598), .B(n_650), .C(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g688 ( .A(n_598), .Y(n_688) );
AOI33xp33_ASAP7_75t_L g1029 ( .A1(n_598), .A2(n_608), .A3(n_1030), .B1(n_1031), .B2(n_1032), .B3(n_1033), .Y(n_1029) );
NAND3xp33_ASAP7_75t_L g1081 ( .A(n_598), .B(n_1082), .C(n_1083), .Y(n_1081) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_605), .C(n_608), .Y(n_600) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g907 ( .A(n_607), .Y(n_907) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_608), .B(n_653), .C(n_656), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g1085 ( .A(n_608), .B(n_1086), .C(n_1087), .Y(n_1085) );
AOI33xp33_ASAP7_75t_L g1135 ( .A1(n_608), .A2(n_916), .A3(n_1136), .B1(n_1138), .B2(n_1141), .B3(n_1142), .Y(n_1135) );
INVx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .C(n_615), .Y(n_611) );
HB1xp67_ASAP7_75t_L g1582 ( .A(n_613), .Y(n_1582) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_615), .B(n_658), .C(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g745 ( .A(n_615), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g1090 ( .A(n_615), .B(n_1091), .C(n_1093), .Y(n_1090) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g1152 ( .A(n_636), .Y(n_1152) );
INVx1_ASAP7_75t_L g898 ( .A(n_638), .Y(n_898) );
NAND4xp25_ASAP7_75t_L g644 ( .A(n_645), .B(n_649), .C(n_652), .D(n_657), .Y(n_644) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g878 ( .A(n_655), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_721), .B1(n_771), .B2(n_772), .Y(n_660) );
INVx1_ASAP7_75t_L g771 ( .A(n_661), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_705), .C(n_714), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_689), .Y(n_663) );
OAI33xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .A3(n_673), .B1(n_680), .B2(n_684), .B3(n_688), .Y(n_664) );
OAI33xp33_ASAP7_75t_L g746 ( .A1(n_665), .A2(n_688), .A3(n_747), .B1(n_750), .B2(n_751), .B3(n_755), .Y(n_746) );
OAI33xp33_ASAP7_75t_L g917 ( .A1(n_665), .A2(n_918), .A3(n_920), .B1(n_929), .B2(n_935), .B3(n_940), .Y(n_917) );
OAI33xp33_ASAP7_75t_L g1442 ( .A1(n_665), .A2(n_1443), .A3(n_1446), .B1(n_1452), .B2(n_1455), .B3(n_1458), .Y(n_1442) );
OAI22xp5_ASAP7_75t_L g1566 ( .A1(n_665), .A2(n_915), .B1(n_1567), .B2(n_1575), .Y(n_1566) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_670), .B2(n_672), .Y(n_667) );
OAI22xp33_ASAP7_75t_L g918 ( .A1(n_668), .A2(n_904), .B1(n_905), .B2(n_919), .Y(n_918) );
OAI22xp33_ASAP7_75t_SL g1561 ( .A1(n_668), .A2(n_1562), .B1(n_1563), .B2(n_1564), .Y(n_1561) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_669), .A2(n_672), .B1(n_691), .B2(n_692), .C(n_695), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_670), .A2(n_732), .B1(n_735), .B2(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g806 ( .A(n_670), .Y(n_806) );
BUFx3_ASAP7_75t_L g816 ( .A(n_670), .Y(n_816) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI22xp33_ASAP7_75t_SL g673 ( .A1(n_674), .A2(n_675), .B1(n_677), .B2(n_678), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_675), .A2(n_681), .B1(n_682), .B2(n_683), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_675), .A2(n_682), .B1(n_726), .B2(n_729), .Y(n_750) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g752 ( .A(n_676), .Y(n_752) );
INVx1_ASAP7_75t_L g1557 ( .A(n_676), .Y(n_1557) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_682), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_686), .A2(n_936), .B1(n_938), .B2(n_939), .Y(n_935) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx2_ASAP7_75t_L g911 ( .A(n_694), .Y(n_911) );
BUFx3_ASAP7_75t_L g826 ( .A(n_696), .Y(n_826) );
BUFx2_ASAP7_75t_L g865 ( .A(n_696), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_700), .B2(n_702), .C(n_703), .Y(n_697) );
INVx2_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g996 ( .A(n_704), .Y(n_996) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g1137 ( .A(n_710), .Y(n_1137) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g919 ( .A(n_718), .Y(n_919) );
INVx2_ASAP7_75t_L g1564 ( .A(n_718), .Y(n_1564) );
INVx1_ASAP7_75t_L g772 ( .A(n_721), .Y(n_772) );
NAND3xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_758), .C(n_766), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_746), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_729), .B2(n_730), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
BUFx4f_ASAP7_75t_L g1139 ( .A(n_728), .Y(n_1139) );
BUFx2_ASAP7_75t_L g1479 ( .A(n_728), .Y(n_1479) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_735), .B2(n_736), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_733), .A2(n_736), .B1(n_739), .B2(n_740), .Y(n_738) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g997 ( .A(n_743), .Y(n_997) );
INVx1_ASAP7_75t_L g1005 ( .A(n_743), .Y(n_1005) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g1474 ( .A(n_763), .Y(n_1474) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_833), .B1(n_834), .B2(n_885), .Y(n_773) );
INVx1_ASAP7_75t_L g885 ( .A(n_774), .Y(n_885) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_798), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_793), .B(n_796), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI21xp33_ASAP7_75t_SL g1583 ( .A1(n_790), .A2(n_1584), .B(n_1585), .Y(n_1583) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
OAI31xp33_ASAP7_75t_L g1103 ( .A1(n_797), .A2(n_1104), .A3(n_1105), .B(n_1109), .Y(n_1103) );
OAI31xp33_ASAP7_75t_L g1540 ( .A1(n_797), .A2(n_1541), .A3(n_1542), .B(n_1546), .Y(n_1540) );
CKINVDCx5p33_ASAP7_75t_R g1451 ( .A(n_800), .Y(n_1451) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
OAI22xp33_ASAP7_75t_SL g811 ( .A1(n_812), .A2(n_813), .B1(n_814), .B2(n_815), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g1452 ( .A1(n_813), .A2(n_1448), .B1(n_1453), .B2(n_1454), .Y(n_1452) );
BUFx3_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g1458 ( .A(n_817), .Y(n_1458) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx2_ASAP7_75t_SL g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g884 ( .A(n_836), .Y(n_884) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g972 ( .A(n_844), .Y(n_972) );
INVx1_ASAP7_75t_L g981 ( .A(n_844), .Y(n_981) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND4xp25_ASAP7_75t_SL g851 ( .A(n_852), .B(n_853), .C(n_855), .D(n_857), .Y(n_851) );
NAND4xp25_ASAP7_75t_L g953 ( .A(n_852), .B(n_954), .C(n_957), .D(n_960), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_879), .Y(n_861) );
INVx2_ASAP7_75t_SL g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g1140 ( .A(n_867), .Y(n_1140) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
BUFx2_ASAP7_75t_L g914 ( .A(n_868), .Y(n_914) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
OR2x2_ASAP7_75t_L g1514 ( .A(n_869), .B(n_1485), .Y(n_1514) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
BUFx6f_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
BUFx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVxp67_ASAP7_75t_SL g1167 ( .A(n_886), .Y(n_1167) );
XNOR2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_1009), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_948), .B2(n_949), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
HB1xp67_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g946 ( .A(n_891), .Y(n_946) );
NAND3xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_901), .C(n_941), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_917), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_910), .B1(n_911), .B2(n_912), .C(n_913), .Y(n_908) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_916), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_921), .A2(n_922), .B1(n_925), .B2(n_926), .Y(n_920) );
INVx2_ASAP7_75t_SL g922 ( .A(n_923), .Y(n_922) );
INVx2_ASAP7_75t_L g931 ( .A(n_923), .Y(n_931) );
BUFx3_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g1449 ( .A(n_924), .Y(n_1449) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx3_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g934 ( .A(n_928), .Y(n_934) );
INVx2_ASAP7_75t_L g1560 ( .A(n_928), .Y(n_1560) );
INVx2_ASAP7_75t_L g1572 ( .A(n_928), .Y(n_1572) );
OAI22xp5_ASAP7_75t_SL g929 ( .A1(n_930), .A2(n_931), .B1(n_932), .B2(n_933), .Y(n_929) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx2_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g1008 ( .A(n_952), .Y(n_1008) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
NAND4xp25_ASAP7_75t_L g975 ( .A(n_976), .B(n_982), .C(n_990), .D(n_998), .Y(n_975) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx2_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
BUFx2_ASAP7_75t_L g1160 ( .A(n_989), .Y(n_1160) );
AND2x4_ASAP7_75t_L g1415 ( .A(n_989), .B(n_1416), .Y(n_1415) );
INVx4_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g1092 ( .A(n_993), .Y(n_1092) );
INVx2_ASAP7_75t_L g1476 ( .A(n_993), .Y(n_1476) );
INVx2_ASAP7_75t_SL g995 ( .A(n_996), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g998 ( .A(n_999), .B(n_1003), .C(n_1006), .Y(n_998) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
XNOR2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1052), .Y(n_1010) );
INVx2_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1013), .Y(n_1051) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1034), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1110), .B1(n_1164), .B2(n_1165), .Y(n_1052) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1053), .Y(n_1164) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1056), .Y(n_1102) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1064), .Y(n_1097) );
INVxp67_ASAP7_75t_L g1104 ( .A(n_1068), .Y(n_1104) );
INVxp67_ASAP7_75t_L g1109 ( .A(n_1074), .Y(n_1109) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
NAND3xp33_ASAP7_75t_L g1095 ( .A(n_1077), .B(n_1096), .C(n_1103), .Y(n_1095) );
AND4x1_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1081), .C(n_1085), .D(n_1090), .Y(n_1077) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1107), .Y(n_1117) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1110), .Y(n_1165) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
NAND3xp33_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1118), .C(n_1121), .Y(n_1113) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1143), .Y(n_1134) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1148), .Y(n_1158) );
BUFx2_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
OAI22xp33_ASAP7_75t_L g1279 ( .A1(n_1163), .A2(n_1280), .B1(n_1281), .B2(n_1282), .Y(n_1279) );
OAI221xp5_ASAP7_75t_L g1168 ( .A1(n_1169), .A2(n_1407), .B1(n_1408), .B2(n_1519), .C(n_1524), .Y(n_1168) );
NOR2x1_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1347), .Y(n_1169) );
NAND4xp25_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1284), .C(n_1311), .D(n_1324), .Y(n_1170) );
A2O1A1Ixp33_ASAP7_75t_L g1171 ( .A1(n_1172), .A2(n_1197), .B(n_1227), .C(n_1273), .Y(n_1171) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1172), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1172), .B(n_1261), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1172), .B(n_1231), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1172), .B(n_1335), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1193), .Y(n_1172) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1173), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1173), .B(n_1194), .Y(n_1269) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1174), .B(n_1194), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1174), .B(n_1288), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1187), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1182), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
OR2x2_ASAP7_75t_L g1223 ( .A(n_1178), .B(n_1183), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1181), .Y(n_1178) );
HB1xp67_ASAP7_75t_L g1530 ( .A(n_1179), .Y(n_1530) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1181), .Y(n_1191) );
AND2x4_ASAP7_75t_L g1184 ( .A(n_1182), .B(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1183), .B(n_1186), .Y(n_1226) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
AND2x4_ASAP7_75t_L g1192 ( .A(n_1189), .B(n_1191), .Y(n_1192) );
AND2x4_ASAP7_75t_L g1204 ( .A(n_1189), .B(n_1190), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g1528 ( .A(n_1190), .Y(n_1528) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1192), .Y(n_1213) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1194), .Y(n_1230) );
INVxp67_ASAP7_75t_SL g1288 ( .A(n_1194), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1194), .B(n_1231), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1196), .Y(n_1194) );
NOR2xp33_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1215), .Y(n_1197) );
OAI221xp5_ASAP7_75t_L g1397 ( .A1(n_1198), .A2(n_1398), .B1(n_1403), .B2(n_1404), .C(n_1405), .Y(n_1397) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1208), .Y(n_1198) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1199), .Y(n_1268) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1199), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1205), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1200), .B(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1201), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1201), .B(n_1205), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1201), .B(n_1208), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1201), .B(n_1237), .Y(n_1300) );
BUFx6f_ASAP7_75t_L g1312 ( .A(n_1201), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1203), .Y(n_1201) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1204), .Y(n_1211) );
BUFx3_ASAP7_75t_L g1277 ( .A(n_1204), .Y(n_1277) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1205), .Y(n_1237) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1205), .Y(n_1251) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1205), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1205), .B(n_1240), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1205), .B(n_1217), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1207), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1208), .B(n_1236), .Y(n_1235) );
CKINVDCx6p67_ASAP7_75t_R g1240 ( .A(n_1208), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1208), .B(n_1246), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1208), .B(n_1241), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1208), .B(n_1241), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1208), .B(n_1250), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1208), .B(n_1275), .Y(n_1403) );
OR2x6_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1210), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1209), .B(n_1210), .Y(n_1265) );
OAI22xp5_ASAP7_75t_SL g1210 ( .A1(n_1211), .A2(n_1212), .B1(n_1213), .B2(n_1214), .Y(n_1210) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1213), .Y(n_1219) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1213), .Y(n_1278) );
XNOR2xp5_ASAP7_75t_L g1409 ( .A(n_1214), .B(n_1410), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1215), .B(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1216), .B(n_1260), .Y(n_1292) );
NOR2xp33_ASAP7_75t_L g1399 ( .A(n_1216), .B(n_1400), .Y(n_1399) );
BUFx3_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx2_ASAP7_75t_SL g1247 ( .A(n_1217), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1217), .B(n_1257), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1272 ( .A(n_1217), .B(n_1237), .Y(n_1272) );
BUFx2_ASAP7_75t_L g1320 ( .A(n_1217), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1217), .B(n_1231), .Y(n_1335) );
INVx2_ASAP7_75t_SL g1217 ( .A(n_1218), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1218), .B(n_1237), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1218), .B(n_1261), .Y(n_1289) );
OAI22xp33_ASAP7_75t_L g1220 ( .A1(n_1221), .A2(n_1222), .B1(n_1224), .B2(n_1225), .Y(n_1220) );
BUFx3_ASAP7_75t_L g1281 ( .A(n_1222), .Y(n_1281) );
BUFx6f_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
HB1xp67_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1226), .Y(n_1283) );
OAI211xp5_ASAP7_75t_L g1227 ( .A1(n_1228), .A2(n_1234), .B(n_1238), .C(n_1267), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1231), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1230), .B(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1230), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1387 ( .A(n_1230), .B(n_1231), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1231), .B(n_1243), .Y(n_1242) );
CKINVDCx5p33_ASAP7_75t_R g1261 ( .A(n_1231), .Y(n_1261) );
HB1xp67_ASAP7_75t_L g1314 ( .A(n_1231), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1231), .B(n_1252), .Y(n_1326) );
NOR2xp33_ASAP7_75t_L g1342 ( .A(n_1231), .B(n_1253), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1231), .B(n_1287), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1231), .B(n_1253), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1374 ( .A(n_1231), .B(n_1375), .Y(n_1374) );
AND2x4_ASAP7_75t_SL g1231 ( .A(n_1232), .B(n_1233), .Y(n_1231) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
AOI221xp5_ASAP7_75t_L g1360 ( .A1(n_1235), .A2(n_1287), .B1(n_1361), .B2(n_1362), .C(n_1363), .Y(n_1360) );
NAND3xp33_ASAP7_75t_L g1307 ( .A(n_1236), .B(n_1308), .C(n_1309), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_1236), .A2(n_1251), .B1(n_1351), .B2(n_1389), .C(n_1392), .Y(n_1388) );
AOI211xp5_ASAP7_75t_L g1238 ( .A1(n_1239), .A2(n_1242), .B(n_1244), .C(n_1262), .Y(n_1238) );
AOI331xp33_ASAP7_75t_L g1311 ( .A1(n_1239), .A2(n_1273), .A3(n_1286), .B1(n_1312), .B2(n_1313), .B3(n_1318), .C1(n_1321), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1241), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1240), .B(n_1300), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1240), .B(n_1274), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1241), .B(n_1274), .Y(n_1294) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1241), .Y(n_1337) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1242), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1242), .B(n_1319), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1243), .B(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1243), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1243), .B(n_1272), .Y(n_1271) );
OAI321xp33_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1248), .A3(n_1252), .B1(n_1254), .B2(n_1255), .C(n_1258), .Y(n_1244) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1245), .Y(n_1308) );
INVxp67_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1247), .B(n_1326), .Y(n_1325) );
NOR2xp33_ASAP7_75t_L g1354 ( .A(n_1247), .B(n_1355), .Y(n_1354) );
HB1xp67_ASAP7_75t_L g1358 ( .A(n_1247), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1247), .B(n_1269), .Y(n_1391) );
O2A1O1Ixp33_ASAP7_75t_SL g1301 ( .A1(n_1248), .A2(n_1273), .B(n_1302), .C(n_1304), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1248), .B(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1249), .Y(n_1330) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1250), .B(n_1286), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1250), .B(n_1334), .Y(n_1333) );
INVx3_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_1251), .B(n_1290), .Y(n_1328) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
AOI222xp33_ASAP7_75t_L g1398 ( .A1(n_1253), .A2(n_1259), .B1(n_1312), .B2(n_1399), .C1(n_1401), .C2(n_1402), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1257), .B(n_1353), .Y(n_1352) );
OAI221xp5_ASAP7_75t_SL g1383 ( .A1(n_1257), .A2(n_1384), .B1(n_1386), .B2(n_1387), .C(n_1388), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1259), .B(n_1320), .Y(n_1394) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1259), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1261), .B(n_1287), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1261), .B(n_1269), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1261), .B(n_1354), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1390 ( .A(n_1261), .B(n_1391), .Y(n_1390) );
NOR2xp33_ASAP7_75t_L g1392 ( .A(n_1261), .B(n_1393), .Y(n_1392) );
NOR3xp33_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1265), .C(n_1266), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
A2O1A1Ixp33_ASAP7_75t_L g1267 ( .A1(n_1265), .A2(n_1268), .B(n_1269), .C(n_1270), .Y(n_1267) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_1265), .B(n_1322), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1266), .B(n_1317), .Y(n_1316) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1266), .B(n_1367), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1269), .B(n_1289), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1269), .B(n_1335), .Y(n_1385) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1272), .B(n_1323), .Y(n_1322) );
INVx3_ASAP7_75t_L g1381 ( .A(n_1273), .Y(n_1381) );
A2O1A1Ixp33_ASAP7_75t_L g1405 ( .A1(n_1273), .A2(n_1330), .B(n_1336), .C(n_1406), .Y(n_1405) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1336 ( .A(n_1276), .B(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1278), .Y(n_1407) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
AOI221xp5_ASAP7_75t_L g1284 ( .A1(n_1285), .A2(n_1290), .B1(n_1291), .B2(n_1293), .C(n_1295), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1289), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1287), .B(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1287), .Y(n_1355) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1289), .Y(n_1367) );
AOI21xp5_ASAP7_75t_L g1369 ( .A1(n_1290), .A2(n_1370), .B(n_1376), .Y(n_1369) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
OAI221xp5_ASAP7_75t_L g1295 ( .A1(n_1296), .A2(n_1298), .B1(n_1301), .B2(n_1305), .C(n_1307), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1296), .B(n_1339), .Y(n_1361) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1300), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1300), .B(n_1320), .Y(n_1386) );
CKINVDCx5p33_ASAP7_75t_R g1302 ( .A(n_1303), .Y(n_1302) );
AOI211xp5_ASAP7_75t_L g1348 ( .A1(n_1304), .A2(n_1349), .B(n_1352), .C(n_1356), .Y(n_1348) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
NOR2xp33_ASAP7_75t_L g1378 ( .A(n_1310), .B(n_1379), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1312), .B(n_1378), .Y(n_1377) );
NOR2xp33_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1315), .Y(n_1313) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1319), .B(n_1374), .Y(n_1402) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1320), .B(n_1337), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1320), .B(n_1374), .Y(n_1373) );
AOI221xp5_ASAP7_75t_L g1324 ( .A1(n_1325), .A2(n_1327), .B1(n_1329), .B2(n_1336), .C(n_1338), .Y(n_1324) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
OAI21xp33_ASAP7_75t_L g1329 ( .A1(n_1330), .A2(n_1331), .B(n_1333), .Y(n_1329) );
OAI21xp33_ASAP7_75t_L g1370 ( .A1(n_1330), .A2(n_1371), .B(n_1373), .Y(n_1370) );
AOI21xp33_ASAP7_75t_SL g1356 ( .A1(n_1331), .A2(n_1357), .B(n_1359), .Y(n_1356) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
AOI21xp5_ASAP7_75t_L g1338 ( .A1(n_1339), .A2(n_1340), .B(n_1343), .Y(n_1338) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
HB1xp67_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
A2O1A1Ixp33_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1360), .B(n_1380), .C(n_1382), .Y(n_1347) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1351), .B(n_1358), .Y(n_1357) );
A2O1A1Ixp33_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1366), .B(n_1368), .C(n_1369), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
NOR2xp33_ASAP7_75t_L g1384 ( .A(n_1365), .B(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
AOI21xp33_ASAP7_75t_SL g1382 ( .A1(n_1383), .A2(n_1395), .B(n_1397), .Y(n_1382) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVxp67_ASAP7_75t_L g1404 ( .A(n_1402), .Y(n_1404) );
HB1xp67_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1459), .Y(n_1410) );
NOR3xp33_ASAP7_75t_SL g1411 ( .A(n_1412), .B(n_1426), .C(n_1442), .Y(n_1411) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
BUFx2_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1422), .B1(n_1423), .B2(n_1424), .Y(n_1420) );
BUFx2_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
INVx2_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
NAND2x1_ASAP7_75t_SL g1429 ( .A(n_1430), .B(n_1432), .Y(n_1429) );
INVx2_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
NAND2x1p5_ASAP7_75t_L g1437 ( .A(n_1432), .B(n_1438), .Y(n_1437) );
INVx3_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
HB1xp67_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
BUFx4f_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
BUFx2_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
OAI22xp5_ASAP7_75t_L g1446 ( .A1(n_1447), .A2(n_1448), .B1(n_1450), .B2(n_1451), .Y(n_1446) );
BUFx2_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
AOI221xp5_ASAP7_75t_SL g1471 ( .A1(n_1453), .A2(n_1472), .B1(n_1478), .B2(n_1481), .C(n_1486), .Y(n_1471) );
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_1454), .A2(n_1456), .B1(n_1511), .B2(n_1513), .Y(n_1510) );
AOI221xp5_ASAP7_75t_L g1494 ( .A1(n_1457), .A2(n_1495), .B1(n_1502), .B2(n_1503), .C(n_1506), .Y(n_1494) );
AOI21xp5_ASAP7_75t_L g1459 ( .A1(n_1460), .A2(n_1469), .B(n_1470), .Y(n_1459) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
AND2x4_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1463), .Y(n_1461) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
AND2x4_ASAP7_75t_L g1488 ( .A(n_1466), .B(n_1489), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1466), .B(n_1493), .Y(n_1492) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1466), .Y(n_1509) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
AOI31xp33_ASAP7_75t_L g1470 ( .A1(n_1471), .A2(n_1494), .A3(n_1510), .B(n_1515), .Y(n_1470) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
HB1xp67_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
INVx2_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx2_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1490), .Y(n_1587) );
INVx3_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1493), .Y(n_1588) );
HB1xp67_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
BUFx6f_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
AND2x4_ASAP7_75t_L g1507 ( .A(n_1499), .B(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_1504), .Y(n_1503) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
HB1xp67_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_SL g1508 ( .A(n_1509), .Y(n_1508) );
INVx6_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
INVx4_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_SL g1515 ( .A(n_1516), .Y(n_1515) );
INVx5_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
BUFx8_ASAP7_75t_SL g1517 ( .A(n_1518), .Y(n_1517) );
CKINVDCx5p33_ASAP7_75t_R g1519 ( .A(n_1520), .Y(n_1519) );
BUFx2_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
HB1xp67_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
A2O1A1Ixp33_ASAP7_75t_L g1526 ( .A1(n_1527), .A2(n_1529), .B(n_1531), .C(n_1532), .Y(n_1526) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVxp33_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
HB1xp67_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
NAND3xp33_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1547), .C(n_1552), .Y(n_1539) );
NOR3xp33_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1566), .C(n_1581), .Y(n_1552) );
NOR3xp33_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1561), .C(n_1565), .Y(n_1553) );
OAI22xp5_ASAP7_75t_L g1554 ( .A1(n_1555), .A2(n_1556), .B1(n_1558), .B2(n_1559), .Y(n_1554) );
BUFx2_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
OAI221xp5_ASAP7_75t_L g1567 ( .A1(n_1568), .A2(n_1570), .B1(n_1571), .B2(n_1573), .C(n_1574), .Y(n_1567) );
INVx2_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
INVx2_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
endmodule