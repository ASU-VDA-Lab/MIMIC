module fake_jpeg_13040_n_668 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_668);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_668;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_1),
.B(n_2),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_61),
.B(n_77),
.Y(n_186)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_19),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_65),
.B(n_80),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_57),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_70),
.Y(n_214)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_71),
.Y(n_201)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_74),
.B(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_78),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_26),
.B(n_19),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_83),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_84),
.Y(n_206)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_85),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_87),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_89),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_41),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_95),
.Y(n_160)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_92),
.Y(n_202)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_93),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_18),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_94),
.B(n_15),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_R g216 ( 
.A(n_98),
.Y(n_216)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_100),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_103),
.Y(n_213)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_105),
.B(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_107),
.Y(n_218)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_108),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_28),
.B(n_16),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_127),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_22),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_113),
.B(n_114),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_22),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_116),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_117),
.Y(n_183)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_120),
.B(n_33),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_22),
.Y(n_122)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_125),
.Y(n_225)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_22),
.B(n_16),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_45),
.Y(n_128)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_22),
.Y(n_129)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_47),
.Y(n_131)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_139),
.Y(n_249)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_149),
.B(n_159),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_61),
.B(n_30),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_71),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_162),
.B(n_163),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_72),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_106),
.B(n_24),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_166),
.B(n_168),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_120),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_167),
.B(n_179),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_102),
.B(n_30),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_170),
.Y(n_252)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_173),
.Y(n_256)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_175),
.Y(n_289)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_177),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_110),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_116),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_180),
.B(n_184),
.Y(n_237)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

CKINVDCx12_ASAP7_75t_R g189 ( 
.A(n_77),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_189),
.Y(n_302)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_190),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_79),
.B(n_45),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_198),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_115),
.B(n_24),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_193),
.B(n_194),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_126),
.B(n_59),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_70),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_69),
.B(n_45),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_130),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_205),
.B1(n_209),
.B2(n_222),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_62),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_208),
.B(n_219),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_82),
.A2(n_33),
.B1(n_36),
.B2(n_44),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_128),
.B(n_59),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_64),
.A2(n_40),
.B1(n_46),
.B2(n_42),
.Y(n_222)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_115),
.B(n_40),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_224),
.B(n_131),
.Y(n_278)
);

OR2x2_ASAP7_75t_SL g226 ( 
.A(n_109),
.B(n_13),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_226),
.B(n_2),
.Y(n_286)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

INVx3_ASAP7_75t_SL g355 ( 
.A(n_228),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_85),
.B1(n_100),
.B2(n_84),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_229),
.A2(n_255),
.B1(n_264),
.B2(n_295),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_186),
.B(n_121),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_230),
.B(n_250),
.Y(n_365)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_153),
.Y(n_231)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_231),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_125),
.B1(n_83),
.B2(n_97),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_236),
.A2(n_248),
.B1(n_158),
.B2(n_212),
.Y(n_336)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_239),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_160),
.B(n_44),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_240),
.B(n_243),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_145),
.B(n_117),
.C(n_119),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_241),
.B(n_258),
.C(n_260),
.Y(n_349)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_155),
.Y(n_242)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_242),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_169),
.B(n_46),
.Y(n_243)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_142),
.Y(n_246)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_246),
.Y(n_315)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_155),
.Y(n_247)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_205),
.A2(n_75),
.B1(n_66),
.B2(n_68),
.Y(n_248)
);

OA22x2_ASAP7_75t_L g344 ( 
.A1(n_248),
.A2(n_206),
.B1(n_203),
.B2(n_221),
.Y(n_344)
);

AND2x2_ASAP7_75t_SL g250 ( 
.A(n_211),
.B(n_63),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_195),
.B(n_39),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_251),
.B(n_262),
.Y(n_363)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_197),
.Y(n_254)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_254),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_138),
.A2(n_209),
.B1(n_101),
.B2(n_96),
.Y(n_255)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_154),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_257),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_174),
.B(n_202),
.C(n_218),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_133),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_78),
.C(n_90),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_144),
.B(n_35),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_261),
.B(n_269),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_134),
.B(n_42),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_132),
.A2(n_89),
.B1(n_35),
.B2(n_39),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_176),
.A2(n_104),
.B1(n_103),
.B2(n_60),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_265),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_154),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_198),
.B(n_63),
.C(n_73),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_268),
.B(n_288),
.C(n_300),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_152),
.B(n_16),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_172),
.B(n_14),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_273),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_14),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_161),
.Y(n_274)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_14),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_275),
.B(n_276),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_156),
.B(n_13),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_150),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_277),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_185),
.Y(n_324)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_164),
.Y(n_279)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_199),
.Y(n_280)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_214),
.Y(n_281)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_214),
.Y(n_282)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_176),
.A2(n_52),
.B1(n_3),
.B2(n_4),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

INVx11_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_284),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_285),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_286),
.B(n_293),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_191),
.A2(n_171),
.B1(n_213),
.B2(n_133),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_287),
.A2(n_303),
.B1(n_183),
.B2(n_141),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_192),
.B(n_157),
.C(n_165),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_135),
.B(n_207),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_294),
.Y(n_337)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_182),
.Y(n_292)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_292),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_147),
.B(n_3),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_148),
.B(n_4),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_148),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g296 ( 
.A(n_223),
.Y(n_296)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_161),
.Y(n_297)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_135),
.B(n_6),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_306),
.Y(n_341)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_155),
.Y(n_299)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_299),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_191),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_187),
.Y(n_301)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_213),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_164),
.Y(n_304)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_147),
.Y(n_305)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

OR2x2_ASAP7_75t_SL g306 ( 
.A(n_139),
.B(n_12),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_132),
.A2(n_12),
.B1(n_188),
.B2(n_212),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_158),
.B1(n_188),
.B2(n_221),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_232),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_318),
.B(n_342),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_230),
.B(n_201),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_319),
.B(n_368),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_324),
.B(n_329),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_227),
.B(n_143),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_253),
.B(n_140),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_330),
.B(n_350),
.Y(n_413)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_234),
.Y(n_334)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_334),
.Y(n_394)
);

AND2x4_ASAP7_75t_SL g335 ( 
.A(n_230),
.B(n_151),
.Y(n_335)
);

OR2x4_ASAP7_75t_L g407 ( 
.A(n_335),
.B(n_279),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_336),
.A2(n_344),
.B1(n_328),
.B2(n_368),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_338),
.A2(n_236),
.B1(n_248),
.B2(n_203),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_237),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_344),
.A2(n_206),
.B1(n_178),
.B2(n_215),
.Y(n_411)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_291),
.Y(n_346)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_346),
.Y(n_395)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_235),
.Y(n_348)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_348),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_258),
.B(n_225),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_271),
.B(n_220),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_359),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_272),
.B(n_200),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_235),
.Y(n_360)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_360),
.Y(n_415)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_233),
.Y(n_364)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_246),
.Y(n_366)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_245),
.B(n_183),
.C(n_141),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_294),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_370),
.B(n_386),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_288),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_371),
.B(n_256),
.C(n_252),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_325),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_372),
.B(n_376),
.Y(n_428)
);

O2A1O1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_328),
.A2(n_250),
.B(n_245),
.C(n_244),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_373),
.A2(n_401),
.B(n_407),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_365),
.A2(n_245),
.B(n_268),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_374),
.A2(n_392),
.B(n_259),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_347),
.Y(n_375)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_375),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_335),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_377),
.A2(n_409),
.B1(n_411),
.B2(n_355),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_381),
.A2(n_410),
.B1(n_280),
.B2(n_345),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_333),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_382),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_340),
.A2(n_267),
.B1(n_239),
.B2(n_277),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_365),
.B(n_341),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_289),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_261),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_340),
.A2(n_267),
.B1(n_249),
.B2(n_263),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_389),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_337),
.B(n_260),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_391),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_250),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_254),
.B(n_300),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_311),
.B(n_249),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_393),
.B(n_408),
.Y(n_425)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_326),
.Y(n_397)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_397),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_335),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_398),
.B(n_414),
.Y(n_456)
);

INVx8_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_400),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_361),
.A2(n_286),
.B(n_306),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_402),
.Y(n_430)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_403),
.Y(n_436)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_352),
.Y(n_404)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_404),
.Y(n_440)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_363),
.B(n_327),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_331),
.A2(n_319),
.B1(n_338),
.B2(n_344),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_344),
.A2(n_248),
.B1(n_241),
.B2(n_136),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_323),
.B(n_249),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_412),
.B(n_302),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_316),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_312),
.A2(n_308),
.B1(n_292),
.B2(n_247),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_416),
.A2(n_281),
.B1(n_282),
.B2(n_285),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_332),
.Y(n_417)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_409),
.A2(n_355),
.B1(n_358),
.B2(n_297),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_418),
.A2(n_437),
.B1(n_444),
.B2(n_447),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_419),
.B(n_383),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_426),
.B(n_442),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_432),
.B(n_383),
.C(n_385),
.Y(n_480)
);

A2O1A1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_386),
.A2(n_313),
.B(n_285),
.C(n_284),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_435),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_373),
.A2(n_339),
.B(n_353),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_434),
.A2(n_407),
.B(n_374),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_390),
.B(n_314),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_410),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_387),
.B(n_339),
.Y(n_442)
);

AOI22x1_ASAP7_75t_SL g443 ( 
.A1(n_381),
.A2(n_353),
.B1(n_369),
.B2(n_308),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_443),
.A2(n_406),
.B(n_392),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_370),
.A2(n_136),
.B1(n_137),
.B2(n_215),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_377),
.A2(n_352),
.B1(n_345),
.B2(n_257),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_391),
.A2(n_137),
.B1(n_178),
.B2(n_274),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_451),
.Y(n_464)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_399),
.Y(n_449)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_399),
.Y(n_450)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_450),
.Y(n_470)
);

OAI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_406),
.A2(n_321),
.B1(n_310),
.B2(n_356),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_452),
.Y(n_491)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_415),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_455),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_380),
.Y(n_455)
);

INVx13_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_458),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_459),
.A2(n_418),
.B1(n_434),
.B2(n_420),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_435),
.B(n_413),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_460),
.B(n_465),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_462),
.A2(n_438),
.B1(n_439),
.B2(n_457),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_455),
.B(n_394),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_378),
.Y(n_466)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_466),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_428),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_467),
.B(n_471),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_427),
.B(n_396),
.Y(n_468)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_468),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_449),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_473),
.B(n_479),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_396),
.Y(n_474)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_474),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_450),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_476),
.B(n_483),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_477),
.A2(n_423),
.B(n_420),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_431),
.B(n_395),
.Y(n_478)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_478),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_431),
.B(n_371),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_479),
.B(n_480),
.C(n_482),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_425),
.B(n_394),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_481),
.B(n_484),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_419),
.B(n_401),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_452),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_395),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_448),
.B(n_454),
.Y(n_485)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_485),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_456),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_486),
.B(n_489),
.Y(n_518)
);

INVx11_ASAP7_75t_L g488 ( 
.A(n_443),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_488),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_445),
.B(n_379),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_442),
.B(n_379),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_492),
.B(n_441),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_445),
.B(n_417),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_493),
.B(n_494),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_433),
.B(n_382),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_467),
.B(n_426),
.Y(n_495)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_495),
.B(n_499),
.C(n_502),
.Y(n_554)
);

AO21x1_ASAP7_75t_L g560 ( 
.A1(n_496),
.A2(n_501),
.B(n_503),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_432),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_463),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_500),
.B(n_529),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_309),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_309),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_505),
.B(n_522),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_459),
.A2(n_457),
.B1(n_439),
.B2(n_436),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_510),
.A2(n_462),
.B1(n_475),
.B2(n_472),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_513),
.B(n_468),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_461),
.A2(n_422),
.B1(n_429),
.B2(n_436),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_515),
.A2(n_519),
.B1(n_485),
.B2(n_474),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_473),
.B(n_440),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_516),
.B(n_528),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_461),
.A2(n_472),
.B1(n_494),
.B2(n_488),
.Y(n_519)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_521),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_466),
.B(n_440),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_480),
.B(n_441),
.C(n_321),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_524),
.B(n_477),
.C(n_489),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_460),
.B(n_403),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_525),
.B(n_526),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_465),
.B(n_405),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_493),
.B(n_478),
.Y(n_527)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_527),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_482),
.B(n_429),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_463),
.Y(n_529)
);

OA21x2_ASAP7_75t_L g530 ( 
.A1(n_488),
.A2(n_453),
.B(n_422),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_530),
.B(n_512),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_531),
.A2(n_530),
.B1(n_512),
.B2(n_514),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_533),
.B(n_536),
.C(n_559),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_534),
.B(n_546),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_459),
.C(n_484),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_508),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_537),
.B(n_545),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_498),
.Y(n_540)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_540),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_506),
.B(n_459),
.Y(n_541)
);

MAJx2_ASAP7_75t_L g581 ( 
.A(n_541),
.B(n_553),
.C(n_555),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_542),
.A2(n_557),
.B1(n_496),
.B2(n_520),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_481),
.Y(n_544)
);

CKINVDCx14_ASAP7_75t_R g571 ( 
.A(n_544),
.Y(n_571)
);

XOR2x2_ASAP7_75t_L g545 ( 
.A(n_513),
.B(n_464),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_506),
.B(n_492),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_508),
.Y(n_547)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_547),
.Y(n_564)
);

AO21x1_ASAP7_75t_L g584 ( 
.A1(n_548),
.A2(n_511),
.B(n_514),
.Y(n_584)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_498),
.Y(n_549)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_549),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_507),
.A2(n_500),
.B1(n_529),
.B2(n_509),
.Y(n_550)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_550),
.Y(n_579)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_518),
.Y(n_552)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_552),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_528),
.B(n_491),
.Y(n_553)
);

MAJx2_ASAP7_75t_L g555 ( 
.A(n_516),
.B(n_464),
.C(n_470),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_518),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_556),
.B(n_558),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_519),
.A2(n_520),
.B1(n_530),
.B2(n_503),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_504),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_501),
.B(n_491),
.C(n_469),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_523),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_561),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_515),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_566),
.B(n_577),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_567),
.A2(n_471),
.B1(n_497),
.B2(n_453),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_535),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_569),
.B(n_572),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_570),
.A2(n_557),
.B1(n_542),
.B2(n_560),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_541),
.B(n_533),
.C(n_543),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_521),
.C(n_507),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_573),
.B(n_586),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_548),
.A2(n_523),
.B(n_510),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_576),
.A2(n_583),
.B(n_458),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_545),
.B(n_536),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_560),
.A2(n_487),
.B(n_517),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_580),
.A2(n_583),
.B(n_575),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_553),
.B(n_527),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_582),
.B(n_555),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_535),
.A2(n_504),
.B(n_517),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_584),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_511),
.C(n_469),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_586),
.Y(n_587)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_587),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_589),
.A2(n_581),
.B1(n_582),
.B2(n_563),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_590),
.B(n_604),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_575),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_591),
.B(n_596),
.Y(n_617)
);

A2O1A1O1Ixp25_ASAP7_75t_L g592 ( 
.A1(n_562),
.A2(n_539),
.B(n_532),
.C(n_534),
.D(n_554),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_592),
.B(n_573),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_571),
.A2(n_538),
.B1(n_540),
.B2(n_483),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_594),
.A2(n_606),
.B1(n_568),
.B2(n_574),
.Y(n_608)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_584),
.Y(n_595)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_595),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_565),
.B(n_551),
.C(n_470),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_565),
.B(n_497),
.C(n_476),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_597),
.B(n_604),
.C(n_588),
.Y(n_620)
);

BUFx12_ASAP7_75t_L g598 ( 
.A(n_576),
.Y(n_598)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_598),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_599),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_601),
.A2(n_607),
.B1(n_598),
.B2(n_596),
.Y(n_625)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_564),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_602),
.B(n_603),
.Y(n_613)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_578),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_566),
.B(n_430),
.Y(n_604)
);

OAI321xp33_ASAP7_75t_L g606 ( 
.A1(n_579),
.A2(n_421),
.A3(n_430),
.B1(n_458),
.B2(n_400),
.C(n_397),
.Y(n_606)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_608),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_593),
.A2(n_585),
.B1(n_570),
.B2(n_580),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_609),
.A2(n_612),
.B1(n_616),
.B2(n_343),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_588),
.B(n_572),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_598),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_593),
.A2(n_574),
.B1(n_567),
.B2(n_577),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_619),
.B(n_620),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_600),
.A2(n_581),
.B(n_563),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_622),
.B(n_285),
.C(n_389),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_597),
.B(n_421),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_623),
.B(n_624),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_599),
.A2(n_375),
.B1(n_402),
.B2(n_404),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_SL g639 ( 
.A1(n_625),
.A2(n_618),
.B1(n_611),
.B2(n_619),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_617),
.B(n_605),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g646 ( 
.A(n_628),
.B(n_632),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_613),
.B(n_592),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_629),
.B(n_631),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_614),
.B(n_590),
.C(n_601),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_610),
.B(n_310),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_633),
.B(n_634),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_621),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_635),
.A2(n_639),
.B1(n_351),
.B2(n_322),
.Y(n_645)
);

NAND2x1_ASAP7_75t_L g647 ( 
.A(n_636),
.B(n_238),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_623),
.B(n_343),
.C(n_356),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_637),
.B(n_615),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_612),
.A2(n_322),
.B(n_320),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_638),
.A2(n_351),
.B(n_242),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_631),
.B(n_620),
.C(n_625),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_640),
.B(n_641),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_630),
.A2(n_618),
.B1(n_624),
.B2(n_615),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_642),
.A2(n_645),
.B1(n_357),
.B2(n_301),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_643),
.A2(n_647),
.B(n_299),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_626),
.B(n_317),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_644),
.B(n_637),
.C(n_627),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_634),
.B(n_639),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g657 ( 
.A(n_650),
.B(n_296),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_651),
.B(n_652),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_640),
.B(n_636),
.C(n_266),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_653),
.B(n_655),
.C(n_656),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_648),
.B(n_317),
.C(n_315),
.Y(n_655)
);

O2A1O1Ixp33_ASAP7_75t_SL g660 ( 
.A1(n_657),
.A2(n_649),
.B(n_647),
.C(n_238),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_654),
.B(n_642),
.C(n_644),
.Y(n_659)
);

MAJx2_ASAP7_75t_L g663 ( 
.A(n_659),
.B(n_654),
.C(n_661),
.Y(n_663)
);

AOI322xp5_ASAP7_75t_L g662 ( 
.A1(n_660),
.A2(n_296),
.A3(n_646),
.B1(n_304),
.B2(n_196),
.C1(n_357),
.C2(n_187),
.Y(n_662)
);

NAND4xp25_ASAP7_75t_SL g664 ( 
.A(n_662),
.B(n_663),
.C(n_201),
.D(n_228),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_664),
.A2(n_658),
.B(n_305),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_665),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_666),
.B(n_315),
.C(n_231),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_667),
.B(n_151),
.Y(n_668)
);


endmodule