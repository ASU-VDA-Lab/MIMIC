module fake_jpeg_25888_n_194 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_50),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_49),
.B1(n_17),
.B2(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_51),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_17),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_65),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_27),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_26),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_21),
.B1(n_3),
.B2(n_6),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_22),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_28),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_28),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_22),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_23),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_37),
.B(n_16),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_81),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_84),
.Y(n_108)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_36),
.B1(n_34),
.B2(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_34),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_34),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_61),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_92),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_21),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_16),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_10),
.B(n_5),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.Y(n_114)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_60),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_55),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_112),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_81),
.C(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_80),
.B(n_14),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_71),
.B1(n_73),
.B2(n_61),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_118),
.B(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_90),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_99),
.B1(n_82),
.B2(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_9),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_3),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_3),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_85),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_98),
.B(n_101),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

AO21x2_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_83),
.B(n_102),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_134),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_118),
.B1(n_122),
.B2(n_115),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_100),
.B(n_81),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_110),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_131),
.C(n_137),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_83),
.Y(n_141)
);

NOR4xp25_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_94),
.C(n_100),
.D(n_64),
.Y(n_158)
);

XNOR2x2_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_86),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_144),
.B(n_108),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_147),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_108),
.A3(n_113),
.B1(n_111),
.B2(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_150),
.B1(n_155),
.B2(n_158),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_113),
.B(n_111),
.C(n_120),
.D(n_123),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_135),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_106),
.B(n_124),
.C(n_116),
.D(n_121),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_139),
.C(n_127),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_152),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_129),
.B1(n_141),
.B2(n_128),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_160),
.B(n_166),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_134),
.C(n_136),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_129),
.B1(n_130),
.B2(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_169),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_150),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_129),
.B1(n_136),
.B2(n_140),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_149),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_172),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_161),
.B(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_162),
.B(n_169),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_183),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_180),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_145),
.B1(n_164),
.B2(n_71),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_163),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_177),
.C(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_187),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_171),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_183),
.A3(n_172),
.B1(n_180),
.B2(n_171),
.C1(n_138),
.C2(n_5),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_6),
.A3(n_7),
.B1(n_13),
.B2(n_73),
.C1(n_103),
.C2(n_96),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_189),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_190),
.C(n_96),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_191),
.Y(n_194)
);


endmodule