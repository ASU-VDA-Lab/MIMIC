module fake_jpeg_25061_n_34 (n_3, n_2, n_1, n_0, n_4, n_5, n_34);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_5),
.Y(n_6)
);

INVx6_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

OAI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_12),
.B(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_14),
.B(n_15),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_7),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_6),
.C(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_17),
.B(n_8),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_7),
.B1(n_11),
.B2(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_11),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_19),
.B1(n_13),
.B2(n_8),
.Y(n_26)
);

AO221x1_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.C(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

AOI221xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.C(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_10),
.B1(n_3),
.B2(n_0),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_26),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.C(n_3),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_29),
.C(n_4),
.Y(n_32)
);

MAJx2_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_10),
.C(n_31),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_10),
.Y(n_34)
);


endmodule