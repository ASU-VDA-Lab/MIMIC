module fake_jpeg_1030_n_538 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_538);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_417;
wire n_362;
wire n_142;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_12),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_57),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_52),
.Y(n_108)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_53),
.Y(n_112)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_12),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_59),
.Y(n_149)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_16),
.B(n_12),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_0),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_75),
.Y(n_127)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_0),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_95),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_88),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_27),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_25),
.Y(n_129)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_15),
.Y(n_93)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_43),
.B(n_1),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_32),
.B1(n_45),
.B2(n_47),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_115),
.A2(n_147),
.B1(n_153),
.B2(n_78),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_51),
.A2(n_45),
.B1(n_17),
.B2(n_47),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_116),
.B(n_129),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_26),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_152),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_50),
.A2(n_25),
.B1(n_27),
.B2(n_37),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_134),
.A2(n_44),
.B1(n_23),
.B2(n_18),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_73),
.A2(n_20),
.B1(n_44),
.B2(n_40),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_18),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_86),
.A2(n_20),
.B1(n_44),
.B2(n_40),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_168),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_44),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_88),
.C(n_37),
.Y(n_186)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_26),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_123),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g256 ( 
.A(n_170),
.B(n_186),
.C(n_196),
.Y(n_256)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_21),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_180),
.Y(n_226)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_24),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_119),
.A2(n_24),
.B(n_42),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_183),
.Y(n_234)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_124),
.A2(n_103),
.B1(n_63),
.B2(n_59),
.Y(n_183)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_106),
.B(n_42),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_134),
.A2(n_129),
.B1(n_116),
.B2(n_115),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_191),
.A2(n_121),
.B1(n_138),
.B2(n_117),
.Y(n_221)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_195),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_194),
.A2(n_166),
.B1(n_162),
.B2(n_17),
.Y(n_243)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_131),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_114),
.B(n_76),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_197),
.B(n_125),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_216),
.B1(n_184),
.B2(n_23),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_131),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_199),
.B(n_202),
.Y(n_241)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

BUFx24_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_79),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_205),
.B(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_109),
.B(n_31),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_165),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_207),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_65),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_213),
.Y(n_246)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_108),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_212),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_165),
.A2(n_83),
.B1(n_55),
.B2(n_84),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_110),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_116),
.A2(n_74),
.B1(n_94),
.B2(n_93),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_113),
.B(n_31),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_218),
.Y(n_249)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_112),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_184),
.A2(n_147),
.B1(n_153),
.B2(n_71),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_220),
.A2(n_224),
.B1(n_250),
.B2(n_254),
.Y(n_266)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_221),
.A2(n_205),
.B(n_231),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_118),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_252),
.C(n_201),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_187),
.B(n_141),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_255),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_136),
.B1(n_207),
.B2(n_179),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_133),
.B1(n_130),
.B2(n_160),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_210),
.B1(n_171),
.B2(n_175),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_184),
.A2(n_169),
.B1(n_148),
.B2(n_133),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g251 ( 
.A(n_203),
.B(n_167),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_180),
.B(n_112),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_183),
.A2(n_169),
.B1(n_148),
.B2(n_135),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_176),
.B(n_181),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_274),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_263),
.A2(n_222),
.B1(n_225),
.B2(n_239),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_217),
.B(n_201),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_264),
.A2(n_272),
.B(n_256),
.Y(n_309)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_265),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_190),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_276),
.C(n_261),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_235),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_275),
.Y(n_307)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_224),
.A2(n_223),
.B1(n_234),
.B2(n_220),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_271),
.B1(n_282),
.B2(n_240),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_250),
.A2(n_198),
.B1(n_193),
.B2(n_202),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_200),
.B(n_212),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_230),
.B1(n_249),
.B2(n_245),
.Y(n_273)
);

OA22x2_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_252),
.B1(n_158),
.B2(n_143),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_249),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_235),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_188),
.C(n_172),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_279),
.B(n_281),
.Y(n_300)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_251),
.A2(n_158),
.B1(n_143),
.B2(n_149),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_280),
.A2(n_222),
.B1(n_225),
.B2(n_227),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_SL g281 ( 
.A(n_241),
.B(n_205),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_238),
.A2(n_189),
.B1(n_206),
.B2(n_215),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_243),
.A2(n_185),
.B1(n_136),
.B2(n_208),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_235),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_286),
.Y(n_315)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

OAI22x1_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_221),
.B1(n_243),
.B2(n_251),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_264),
.B(n_284),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_282),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_302),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_296),
.A2(n_299),
.B1(n_304),
.B2(n_310),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_297),
.B(n_276),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_266),
.A2(n_243),
.B1(n_226),
.B2(n_149),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_260),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_266),
.A2(n_226),
.B1(n_135),
.B2(n_246),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_240),
.C(n_242),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_262),
.C(n_269),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_306),
.A2(n_309),
.B(n_311),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_265),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_273),
.A2(n_246),
.B1(n_242),
.B2(n_130),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_262),
.A2(n_255),
.B(n_233),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_277),
.Y(n_312)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_274),
.B(n_244),
.Y(n_316)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_267),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_311),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_261),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_321),
.C(n_335),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_323),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_303),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_325),
.B(n_330),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_312),
.A2(n_283),
.B1(n_259),
.B2(n_271),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_327),
.A2(n_346),
.B1(n_289),
.B2(n_310),
.Y(n_380)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_329),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_315),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_317),
.Y(n_333)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_318),
.A2(n_275),
.B(n_285),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_334),
.B(n_313),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_292),
.B(n_276),
.C(n_257),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_299),
.A2(n_263),
.B1(n_257),
.B2(n_268),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_336),
.A2(n_339),
.B1(n_347),
.B2(n_293),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_341),
.C(n_345),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_299),
.A2(n_280),
.B1(n_287),
.B2(n_286),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_292),
.B(n_281),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_305),
.B(n_219),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_342),
.B(n_302),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_317),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_343),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_315),
.Y(n_344)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_173),
.C(n_174),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_295),
.A2(n_279),
.B1(n_160),
.B2(n_219),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_304),
.A2(n_253),
.B1(n_178),
.B2(n_195),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g349 ( 
.A1(n_307),
.A2(n_314),
.A3(n_313),
.B1(n_316),
.B2(n_296),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_349),
.B(n_307),
.Y(n_351)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_293),
.Y(n_350)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_351),
.A2(n_362),
.B(n_331),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_367),
.C(n_373),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_333),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_359),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_320),
.B(n_311),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_378),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_314),
.Y(n_358)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_324),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_360),
.A2(n_365),
.B1(n_374),
.B2(n_376),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_343),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_363),
.Y(n_398)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_330),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_337),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_304),
.Y(n_366)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_301),
.C(n_309),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_301),
.C(n_300),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_337),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_310),
.Y(n_375)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_334),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_327),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_377),
.A2(n_351),
.B(n_322),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_335),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_380),
.A2(n_322),
.B1(n_332),
.B2(n_328),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_340),
.B(n_298),
.Y(n_381)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_381),
.Y(n_394)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_356),
.B(n_321),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_399),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_345),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_393),
.Y(n_413)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_371),
.Y(n_387)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_387),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_388),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_348),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_395),
.A2(n_401),
.B1(n_358),
.B2(n_369),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_379),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_298),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_348),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_331),
.C(n_323),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_400),
.B(n_402),
.C(n_403),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_332),
.C(n_300),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_301),
.C(n_336),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_301),
.C(n_328),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_407),
.C(n_410),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_301),
.C(n_289),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_379),
.Y(n_408)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_374),
.A2(n_294),
.B(n_326),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_409),
.A2(n_370),
.B(n_376),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_339),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_346),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_411),
.B(n_380),
.C(n_377),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_393),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_384),
.A2(n_360),
.B1(n_370),
.B2(n_375),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_416),
.A2(n_434),
.B1(n_436),
.B2(n_383),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_398),
.B(n_357),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_426),
.Y(n_441)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_418),
.Y(n_448)
);

FAx1_ASAP7_75t_SL g419 ( 
.A(n_390),
.B(n_381),
.CI(n_368),
.CON(n_419),
.SN(n_419)
);

FAx1_ASAP7_75t_SL g443 ( 
.A(n_419),
.B(n_402),
.CI(n_390),
.CON(n_443),
.SN(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_421),
.A2(n_397),
.B1(n_395),
.B2(n_407),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_394),
.A2(n_355),
.B1(n_357),
.B2(n_369),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_423),
.A2(n_431),
.B1(n_410),
.B2(n_391),
.Y(n_440)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_389),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_428),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_371),
.C(n_291),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_382),
.C(n_372),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_430),
.Y(n_453)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_406),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_401),
.A2(n_288),
.B1(n_347),
.B2(n_372),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_397),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_433),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_361),
.C(n_352),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_404),
.A2(n_352),
.B1(n_306),
.B2(n_213),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_385),
.B(n_253),
.C(n_306),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_435),
.B(n_399),
.C(n_403),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_411),
.A2(n_290),
.B1(n_178),
.B2(n_192),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_437),
.A2(n_444),
.B1(n_445),
.B2(n_458),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_442),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_412),
.Y(n_466)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_440),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_400),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_446),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_422),
.A2(n_405),
.B1(n_290),
.B2(n_89),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_433),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_447),
.B(n_449),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_290),
.Y(n_449)
);

INVx11_ASAP7_75t_L g450 ( 
.A(n_419),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_450),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_422),
.A2(n_211),
.B1(n_182),
.B2(n_218),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_452),
.B(n_454),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_413),
.B(n_156),
.C(n_142),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_416),
.A2(n_214),
.B1(n_209),
.B2(n_87),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_431),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_420),
.B(n_236),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_SL g470 ( 
.A(n_456),
.B(n_435),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_434),
.A2(n_258),
.B1(n_236),
.B2(n_96),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_448),
.A2(n_418),
.B(n_428),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_460),
.A2(n_461),
.B(n_463),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_450),
.A2(n_457),
.B(n_440),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_446),
.A2(n_423),
.B(n_415),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_414),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_469),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_466),
.B(n_468),
.Y(n_491)
);

AOI21x1_ASAP7_75t_SL g467 ( 
.A1(n_453),
.A2(n_419),
.B(n_436),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_467),
.A2(n_470),
.B(n_2),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_451),
.A2(n_412),
.B(n_420),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_414),
.C(n_424),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_454),
.C(n_456),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_443),
.A2(n_236),
.B1(n_258),
.B2(n_96),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_473),
.A2(n_97),
.B1(n_3),
.B2(n_4),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_449),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_475),
.B(n_458),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_438),
.B(n_236),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_2),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_461),
.A2(n_443),
.B(n_445),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_479),
.A2(n_489),
.B(n_463),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_480),
.B(n_487),
.Y(n_500)
);

NOR2x1_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_447),
.Y(n_482)
);

NOR2x1_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_478),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_474),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_493),
.Y(n_498)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_484),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_485),
.A2(n_464),
.B1(n_477),
.B2(n_462),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_97),
.C(n_3),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_11),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_488),
.B(n_5),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_467),
.A2(n_2),
.B(n_4),
.Y(n_489)
);

INVx11_ASAP7_75t_L g490 ( 
.A(n_476),
.Y(n_490)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_490),
.Y(n_503)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_492),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_459),
.B(n_4),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_7),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_464),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_5),
.Y(n_507)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_502),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_501),
.A2(n_510),
.B(n_493),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_481),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_481),
.B(n_465),
.C(n_459),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_505),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_491),
.B(n_473),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_506),
.B(n_480),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_495),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_5),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_508),
.A2(n_485),
.B(n_484),
.Y(n_514)
);

A2O1A1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_497),
.A2(n_486),
.B(n_479),
.C(n_489),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_511),
.A2(n_518),
.B(n_519),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_486),
.C(n_492),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_513),
.B(n_514),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_515),
.A2(n_516),
.B(n_517),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_501),
.A2(n_494),
.B(n_487),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_496),
.A2(n_503),
.B(n_500),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_520),
.A2(n_503),
.B(n_498),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_522),
.A2(n_528),
.B(n_507),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_499),
.C(n_498),
.Y(n_524)
);

OA21x2_ASAP7_75t_L g529 ( 
.A1(n_524),
.A2(n_511),
.B(n_509),
.Y(n_529)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_521),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_526),
.B(n_8),
.C(n_9),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_521),
.Y(n_528)
);

NOR3xp33_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_531),
.C(n_527),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_530),
.A2(n_532),
.B(n_525),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_10),
.C(n_8),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_533),
.A2(n_534),
.B(n_535),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_529),
.A2(n_8),
.B(n_9),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_9),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_10),
.Y(n_538)
);


endmodule