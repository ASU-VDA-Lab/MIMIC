module fake_jpeg_16352_n_258 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_46),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_24),
.CON(n_47),
.SN(n_47)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_0),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_35),
.Y(n_71)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_56),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_21),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_25),
.B1(n_33),
.B2(n_24),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_59),
.B1(n_29),
.B2(n_33),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_43),
.B1(n_45),
.B2(n_18),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_28),
.B1(n_20),
.B2(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_67),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_90),
.B(n_27),
.C(n_23),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_41),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_85),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_26),
.B1(n_34),
.B2(n_43),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_92),
.B1(n_94),
.B2(n_36),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_83),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_41),
.B(n_45),
.C(n_40),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_87),
.B1(n_38),
.B2(n_23),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_41),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_21),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_45),
.B(n_40),
.C(n_39),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_93),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_35),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_94),
.Y(n_116)
);

AOI31xp33_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_32),
.A3(n_26),
.B(n_18),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_29),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_98),
.Y(n_123)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_62),
.B1(n_51),
.B2(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_104),
.A2(n_114),
.B1(n_119),
.B2(n_127),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_2),
.C(n_4),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_48),
.C(n_38),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_112),
.C(n_96),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_43),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_84),
.B(n_73),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_38),
.C(n_39),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_87),
.B1(n_71),
.B2(n_80),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_27),
.B1(n_23),
.B2(n_36),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_112),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_36),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_30),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_30),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_100),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_81),
.A2(n_30),
.B1(n_17),
.B2(n_16),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_147),
.Y(n_161)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_104),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_84),
.B1(n_99),
.B2(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_145),
.B(n_111),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_95),
.B(n_80),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_91),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_153),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_17),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_156),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_76),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_13),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_160),
.A2(n_157),
.B1(n_148),
.B2(n_144),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_109),
.C(n_118),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_173),
.C(n_177),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_110),
.B(n_119),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_145),
.B(n_138),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_182),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_108),
.C(n_107),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_181),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_115),
.C(n_127),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_76),
.C(n_96),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_179),
.C(n_151),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_76),
.C(n_9),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_105),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_139),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_188),
.C(n_173),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_160),
.B(n_175),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_189),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_143),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_161),
.B(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_197),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_151),
.A3(n_157),
.B1(n_137),
.B2(n_138),
.Y(n_197)
);

OR2x6_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_141),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_200),
.Y(n_217)
);

OAI322xp33_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_132),
.A3(n_143),
.B1(n_150),
.B2(n_152),
.C1(n_12),
.C2(n_11),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_158),
.A3(n_159),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_9),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_160),
.A2(n_132),
.B(n_133),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_203),
.Y(n_218)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_162),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_207),
.C(n_208),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_198),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_177),
.C(n_176),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_200),
.B(n_198),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_172),
.C(n_167),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_184),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_221),
.B(n_224),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_229),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_231),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_191),
.B1(n_197),
.B2(n_175),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_228),
.A2(n_193),
.B(n_207),
.C(n_11),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_210),
.C(n_215),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_202),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_236),
.C(n_6),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_205),
.C(n_208),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_180),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_238),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_226),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_234),
.A2(n_230),
.B(n_228),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_240),
.A2(n_226),
.B(n_225),
.Y(n_244)
);

NAND4xp25_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_229),
.C(n_10),
.D(n_12),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.C(n_235),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_6),
.Y(n_247)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_238),
.C(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_250),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_243),
.C(n_237),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_252),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_249),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_254),
.A2(n_253),
.B(n_252),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_254),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_255),
.Y(n_258)
);


endmodule