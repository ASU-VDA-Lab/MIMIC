module real_jpeg_2759_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_1),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_1),
.A2(n_42),
.B1(n_58),
.B2(n_59),
.Y(n_91)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_25),
.B1(n_36),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_3),
.A2(n_30),
.B1(n_53),
.B2(n_70),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_3),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_3),
.A2(n_39),
.B1(n_41),
.B2(n_53),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_4),
.B(n_126),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_4),
.B(n_57),
.C(n_59),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_56),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_41),
.C(n_88),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_4),
.A2(n_34),
.B1(n_58),
.B2(n_59),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_4),
.B(n_45),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_4),
.B(n_92),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_25),
.B1(n_34),
.B2(n_36),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_5),
.A2(n_39),
.B1(n_41),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_5),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_25),
.B1(n_36),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_7),
.A2(n_30),
.B1(n_65),
.B2(n_70),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_7),
.A2(n_39),
.B1(n_41),
.B2(n_65),
.Y(n_170)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_9),
.A2(n_39),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_9),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_117)
);

BUFx16f_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_12),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_12),
.A2(n_25),
.B1(n_36),
.B2(n_85),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_12),
.A2(n_39),
.B1(n_41),
.B2(n_85),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_14),
.A2(n_30),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_14),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_14),
.A2(n_25),
.B1(n_36),
.B2(n_69),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_69),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_14),
.A2(n_39),
.B1(n_41),
.B2(n_69),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_15),
.A2(n_39),
.B1(n_41),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_20),
.B(n_106),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_93),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_21),
.B(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_22),
.B(n_50),
.C(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_23),
.A2(n_24),
.B1(n_37),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.A3(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_24)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_25),
.A2(n_36),
.B1(n_57),
.B2(n_61),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_71)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_70),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_30),
.A2(n_33),
.B(n_34),
.C(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_34),
.A2(n_80),
.B(n_181),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_36),
.B(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_37),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_38),
.A2(n_43),
.B1(n_44),
.B2(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_39),
.A2(n_41),
.B1(n_88),
.B2(n_89),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_41),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_43),
.A2(n_44),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_43),
.B(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_43),
.A2(n_179),
.B(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_43),
.A2(n_44),
.B1(n_179),
.B2(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_44),
.A2(n_150),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_44),
.B(n_170),
.Y(n_181)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_47),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_45),
.A2(n_169),
.B(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_66),
.B2(n_77),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B(n_63),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_54),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_54),
.A2(n_63),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_55),
.B(n_64),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

AO22x2_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_59),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_59),
.B(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B(n_72),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_75),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_93),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_83),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_86),
.A2(n_159),
.B(n_161),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_86),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_90),
.A2(n_96),
.B(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_90),
.A2(n_160),
.B1(n_187),
.B2(n_195),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_92),
.B(n_97),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_103),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_94),
.B(n_103),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_98),
.A2(n_99),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_105),
.B(n_130),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_131),
.B2(n_132),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_151),
.B(n_231),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_137),
.B(n_139),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_145),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_145),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.C(n_149),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_173),
.B(n_230),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_171),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_154),
.B(n_171),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_163),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_155),
.B(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_163),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_225),
.B(n_229),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_215),
.B(n_224),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_197),
.B(n_214),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_190),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_190),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_182),
.B1(n_188),
.B2(n_189),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_185),
.C(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_208),
.B(n_213),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_203),
.B(n_207),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_206),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_211),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_217),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_221),
.C(n_222),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_228),
.Y(n_229)
);


endmodule