module real_aes_135_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_0), .B(n_122), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_1), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_2), .A2(n_116), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_3), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_4), .B(n_133), .Y(n_161) );
INVx1_ASAP7_75t_L g121 ( .A(n_5), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_6), .B(n_133), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_7), .B(n_157), .Y(n_563) );
INVx1_ASAP7_75t_L g480 ( .A(n_8), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_9), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_10), .Y(n_496) );
NAND2xp33_ASAP7_75t_L g233 ( .A(n_11), .B(n_131), .Y(n_233) );
INVx2_ASAP7_75t_L g113 ( .A(n_12), .Y(n_113) );
AOI221x1_ASAP7_75t_L g115 ( .A1(n_13), .A2(n_25), .B1(n_116), .B2(n_122), .C(n_129), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_14), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_15), .B(n_122), .Y(n_229) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_16), .A2(n_227), .B(n_228), .Y(n_226) );
INVx1_ASAP7_75t_L g571 ( .A(n_17), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_18), .B(n_111), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_19), .B(n_133), .Y(n_215) );
AO21x1_ASAP7_75t_L g155 ( .A1(n_20), .A2(n_122), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g423 ( .A(n_21), .Y(n_423) );
INVx1_ASAP7_75t_L g569 ( .A(n_22), .Y(n_569) );
INVx1_ASAP7_75t_SL g534 ( .A(n_23), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_24), .B(n_123), .Y(n_555) );
NAND2x1_ASAP7_75t_L g143 ( .A(n_26), .B(n_133), .Y(n_143) );
AOI33xp33_ASAP7_75t_L g508 ( .A1(n_27), .A2(n_54), .A3(n_462), .B1(n_467), .B2(n_509), .B3(n_510), .Y(n_508) );
NAND2x1_ASAP7_75t_L g189 ( .A(n_28), .B(n_131), .Y(n_189) );
INVx1_ASAP7_75t_L g489 ( .A(n_29), .Y(n_489) );
OR2x2_ASAP7_75t_L g114 ( .A(n_30), .B(n_86), .Y(n_114) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_30), .A2(n_86), .B(n_113), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_31), .B(n_470), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_32), .B(n_131), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_33), .A2(n_91), .B1(n_768), .B2(n_769), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_33), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_34), .B(n_133), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_35), .B(n_131), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_36), .A2(n_116), .B(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g117 ( .A(n_37), .B(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g128 ( .A(n_37), .B(n_121), .Y(n_128) );
INVx1_ASAP7_75t_L g461 ( .A(n_37), .Y(n_461) );
OR2x6_ASAP7_75t_L g421 ( .A(n_38), .B(n_422), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_39), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_40), .A2(n_51), .B1(n_412), .B2(n_413), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_40), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_41), .B(n_122), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_42), .B(n_470), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_43), .A2(n_148), .B1(n_157), .B2(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_44), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_45), .B(n_123), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_46), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_47), .B(n_131), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_48), .B(n_227), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_49), .B(n_123), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_50), .A2(n_116), .B(n_188), .Y(n_187) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_51), .A2(n_101), .B1(n_430), .B2(n_437), .C1(n_776), .C2(n_782), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_51), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_52), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_53), .B(n_131), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_55), .B(n_123), .Y(n_520) );
INVx1_ASAP7_75t_L g120 ( .A(n_56), .Y(n_120) );
INVx1_ASAP7_75t_L g125 ( .A(n_56), .Y(n_125) );
AND2x2_ASAP7_75t_L g521 ( .A(n_57), .B(n_111), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_58), .A2(n_74), .B1(n_459), .B2(n_470), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_59), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_60), .B(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_61), .B(n_148), .Y(n_498) );
AOI21xp5_ASAP7_75t_SL g458 ( .A1(n_62), .A2(n_459), .B(n_464), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_63), .A2(n_116), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g566 ( .A(n_64), .Y(n_566) );
AO21x1_ASAP7_75t_L g158 ( .A1(n_65), .A2(n_116), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_66), .B(n_122), .Y(n_179) );
INVx1_ASAP7_75t_L g519 ( .A(n_67), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_68), .B(n_122), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_69), .A2(n_459), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g172 ( .A(n_70), .B(n_112), .Y(n_172) );
INVx1_ASAP7_75t_L g118 ( .A(n_71), .Y(n_118) );
INVx1_ASAP7_75t_L g127 ( .A(n_71), .Y(n_127) );
AND2x2_ASAP7_75t_L g193 ( .A(n_72), .B(n_147), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_73), .B(n_470), .Y(n_511) );
AND2x2_ASAP7_75t_L g536 ( .A(n_75), .B(n_147), .Y(n_536) );
INVx1_ASAP7_75t_L g567 ( .A(n_76), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_77), .A2(n_459), .B(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_SL g770 ( .A1(n_78), .A2(n_767), .B1(n_771), .B2(n_774), .Y(n_770) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_79), .A2(n_459), .B(n_503), .C(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g424 ( .A(n_80), .Y(n_424) );
AND2x2_ASAP7_75t_L g177 ( .A(n_81), .B(n_147), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_82), .B(n_122), .Y(n_217) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_83), .B(n_147), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_84), .A2(n_459), .B1(n_506), .B2(n_507), .Y(n_505) );
AND2x2_ASAP7_75t_L g156 ( .A(n_85), .B(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g150 ( .A(n_87), .B(n_147), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_88), .B(n_131), .Y(n_216) );
INVx1_ASAP7_75t_L g465 ( .A(n_89), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_90), .B(n_133), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_91), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_92), .B(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_93), .A2(n_116), .B(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g512 ( .A(n_94), .B(n_147), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_95), .B(n_133), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_96), .A2(n_487), .B(n_488), .C(n_491), .Y(n_486) );
BUFx2_ASAP7_75t_L g436 ( .A(n_97), .Y(n_436) );
BUFx2_ASAP7_75t_SL g786 ( .A(n_97), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_98), .A2(n_116), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_99), .B(n_123), .Y(n_468) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_416), .B(n_425), .Y(n_102) );
OAI22xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_411), .B1(n_414), .B2(n_415), .Y(n_103) );
INVx3_ASAP7_75t_L g414 ( .A(n_104), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_104), .A2(n_448), .B1(n_772), .B2(n_773), .Y(n_771) );
NAND4xp75_ASAP7_75t_L g104 ( .A(n_105), .B(n_321), .C(n_361), .D(n_390), .Y(n_104) );
NOR2x1_ASAP7_75t_L g105 ( .A(n_106), .B(n_283), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_240), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_173), .B(n_194), .Y(n_107) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_136), .Y(n_108) );
AND2x4_ASAP7_75t_L g239 ( .A(n_109), .B(n_199), .Y(n_239) );
INVx1_ASAP7_75t_SL g292 ( .A(n_109), .Y(n_292) );
AOI21xp33_ASAP7_75t_L g327 ( .A1(n_109), .A2(n_328), .B(n_331), .Y(n_327) );
A2O1A1Ixp33_ASAP7_75t_SL g331 ( .A1(n_109), .A2(n_332), .B(n_333), .C(n_334), .Y(n_331) );
NAND2x1_ASAP7_75t_L g372 ( .A(n_109), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_109), .B(n_333), .Y(n_394) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g197 ( .A(n_110), .Y(n_197) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_110), .Y(n_271) );
OA21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_115), .B(n_135), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_111), .A2(n_179), .B(n_180), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_111), .Y(n_192) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_111), .A2(n_115), .B(n_135), .Y(n_281) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x4_ASAP7_75t_L g157 ( .A(n_113), .B(n_114), .Y(n_157) );
AND2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
BUFx3_ASAP7_75t_L g473 ( .A(n_117), .Y(n_473) );
AND2x6_ASAP7_75t_L g131 ( .A(n_118), .B(n_124), .Y(n_131) );
INVx2_ASAP7_75t_L g463 ( .A(n_118), .Y(n_463) );
AND2x4_ASAP7_75t_L g459 ( .A(n_119), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x4_ASAP7_75t_L g133 ( .A(n_120), .B(n_126), .Y(n_133) );
INVx2_ASAP7_75t_L g467 ( .A(n_120), .Y(n_467) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_121), .Y(n_472) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_128), .Y(n_122) );
INVx1_ASAP7_75t_L g490 ( .A(n_123), .Y(n_490) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx5_ASAP7_75t_L g134 ( .A(n_128), .Y(n_134) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_128), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_132), .B(n_134), .Y(n_129) );
INVxp67_ASAP7_75t_L g570 ( .A(n_131), .Y(n_570) );
INVxp67_ASAP7_75t_L g572 ( .A(n_133), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_134), .A2(n_143), .B(n_144), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_134), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_134), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_134), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_134), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_134), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_134), .A2(n_232), .B(n_233), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_134), .A2(n_465), .B(n_466), .C(n_468), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_134), .A2(n_466), .B(n_480), .C(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g506 ( .A(n_134), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_134), .A2(n_466), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_134), .A2(n_466), .B(n_534), .C(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_134), .A2(n_555), .B(n_556), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_134), .B(n_157), .Y(n_573) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_151), .Y(n_136) );
AND2x2_ASAP7_75t_L g263 ( .A(n_137), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g344 ( .A(n_137), .B(n_199), .Y(n_344) );
INVx1_ASAP7_75t_L g404 ( .A(n_137), .Y(n_404) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g248 ( .A(n_138), .B(n_164), .Y(n_248) );
AND2x2_ASAP7_75t_L g373 ( .A(n_138), .B(n_165), .Y(n_373) );
AND2x2_ASAP7_75t_L g378 ( .A(n_138), .B(n_338), .Y(n_378) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVxp67_ASAP7_75t_L g254 ( .A(n_139), .Y(n_254) );
BUFx3_ASAP7_75t_L g287 ( .A(n_139), .Y(n_287) );
AND2x2_ASAP7_75t_L g333 ( .A(n_139), .B(n_165), .Y(n_333) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_146), .B(n_150), .Y(n_139) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_140), .A2(n_146), .B(n_150), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_146), .A2(n_166), .B(n_172), .Y(n_165) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_146), .A2(n_166), .B(n_172), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_146), .A2(n_147), .B1(n_486), .B2(n_492), .Y(n_485) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_146), .A2(n_515), .B(n_521), .Y(n_514) );
AO21x2_ASAP7_75t_L g579 ( .A1(n_146), .A2(n_515), .B(n_521), .Y(n_579) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_148), .B(n_495), .Y(n_494) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx4f_ASAP7_75t_L g227 ( .A(n_149), .Y(n_227) );
AND2x2_ASAP7_75t_L g318 ( .A(n_151), .B(n_196), .Y(n_318) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_164), .Y(n_151) );
AND2x4_ASAP7_75t_L g199 ( .A(n_152), .B(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_L g310 ( .A(n_152), .B(n_294), .Y(n_310) );
AND2x2_ASAP7_75t_SL g353 ( .A(n_152), .B(n_281), .Y(n_353) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx2_ASAP7_75t_L g289 ( .A(n_153), .Y(n_289) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g250 ( .A(n_154), .Y(n_250) );
OAI21x1_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_158), .B(n_162), .Y(n_154) );
INVx1_ASAP7_75t_L g163 ( .A(n_156), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_157), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_SL g211 ( .A(n_157), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_157), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_157), .A2(n_458), .B(n_469), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_164), .B(n_250), .Y(n_253) );
AND2x2_ASAP7_75t_L g338 ( .A(n_164), .B(n_281), .Y(n_338) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g335 ( .A(n_165), .B(n_197), .Y(n_335) );
AND2x2_ASAP7_75t_L g355 ( .A(n_165), .B(n_281), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_167), .B(n_171), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_173), .B(n_244), .Y(n_273) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_173), .A2(n_367), .B1(n_368), .B2(n_369), .C(n_371), .Y(n_366) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OAI332xp33_ASAP7_75t_L g400 ( .A1(n_174), .A2(n_260), .A3(n_267), .B1(n_326), .B2(n_401), .B3(n_402), .C1(n_403), .C2(n_405), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g174 ( .A(n_175), .B(n_184), .Y(n_174) );
AND2x2_ASAP7_75t_L g205 ( .A(n_175), .B(n_185), .Y(n_205) );
AND2x2_ASAP7_75t_L g222 ( .A(n_175), .B(n_223), .Y(n_222) );
INVx4_ASAP7_75t_L g235 ( .A(n_175), .Y(n_235) );
AND2x2_ASAP7_75t_SL g295 ( .A(n_175), .B(n_236), .Y(n_295) );
INVx5_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2x1_ASAP7_75t_SL g257 ( .A(n_176), .B(n_223), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_176), .B(n_184), .Y(n_261) );
AND2x2_ASAP7_75t_L g268 ( .A(n_176), .B(n_185), .Y(n_268) );
BUFx2_ASAP7_75t_L g303 ( .A(n_176), .Y(n_303) );
AND2x2_ASAP7_75t_L g358 ( .A(n_176), .B(n_226), .Y(n_358) );
OR2x6_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
OR2x2_ASAP7_75t_L g225 ( .A(n_184), .B(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g236 ( .A(n_184), .B(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g276 ( .A(n_184), .Y(n_276) );
AND2x2_ASAP7_75t_L g346 ( .A(n_184), .B(n_245), .Y(n_346) );
AND2x2_ASAP7_75t_L g359 ( .A(n_184), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_184), .B(n_360), .Y(n_377) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_185), .Y(n_243) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_192), .B(n_193), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_191), .Y(n_186) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_192), .A2(n_530), .B(n_536), .Y(n_529) );
OAI32xp33_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_201), .A3(n_206), .B1(n_220), .B2(n_238), .Y(n_194) );
INVx2_ASAP7_75t_L g304 ( .A(n_195), .Y(n_304) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_198), .Y(n_195) );
INVx1_ASAP7_75t_L g315 ( .A(n_196), .Y(n_315) );
BUFx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x4_ASAP7_75t_L g249 ( .A(n_197), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g382 ( .A(n_197), .B(n_287), .Y(n_382) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g294 ( .A(n_200), .Y(n_294) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_205), .Y(n_202) );
INVx2_ASAP7_75t_L g282 ( .A(n_203), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_203), .B(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_SL g293 ( .A(n_204), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g370 ( .A(n_204), .Y(n_370) );
AND2x2_ASAP7_75t_L g388 ( .A(n_204), .B(n_250), .Y(n_388) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp67_ASAP7_75t_SL g332 ( .A(n_207), .B(n_261), .Y(n_332) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_208), .B(n_243), .Y(n_330) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g406 ( .A(n_209), .B(n_276), .Y(n_406) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g237 ( .A(n_210), .Y(n_237) );
INVx2_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_218), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_211), .B(n_219), .Y(n_218) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_211), .A2(n_212), .B(n_218), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_217), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_234), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_221), .B(n_280), .Y(n_365) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
AND3x2_ASAP7_75t_L g320 ( .A(n_222), .B(n_267), .C(n_276), .Y(n_320) );
AND2x2_ASAP7_75t_L g244 ( .A(n_223), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_223), .B(n_226), .Y(n_301) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g255 ( .A(n_225), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g245 ( .A(n_226), .Y(n_245) );
INVx1_ASAP7_75t_L g260 ( .A(n_226), .Y(n_260) );
BUFx3_ASAP7_75t_L g267 ( .A(n_226), .Y(n_267) );
AND2x2_ASAP7_75t_L g277 ( .A(n_226), .B(n_278), .Y(n_277) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_227), .A2(n_478), .B(n_482), .Y(n_477) );
INVx2_ASAP7_75t_SL g503 ( .A(n_227), .Y(n_503) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AND2x4_ASAP7_75t_L g286 ( .A(n_235), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_235), .B(n_245), .Y(n_329) );
AND2x2_ASAP7_75t_L g285 ( .A(n_236), .B(n_260), .Y(n_285) );
INVx2_ASAP7_75t_L g312 ( .A(n_236), .Y(n_312) );
INVx1_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
AOI211xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_246), .B(n_251), .C(n_272), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_241), .A2(n_368), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_244), .B(n_303), .Y(n_302) );
AOI211xp5_ASAP7_75t_SL g322 ( .A1(n_244), .A2(n_323), .B(n_327), .C(n_336), .Y(n_322) );
AND2x2_ASAP7_75t_L g308 ( .A(n_245), .B(n_268), .Y(n_308) );
OR2x2_ASAP7_75t_L g311 ( .A(n_245), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_248), .B(n_353), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_249), .B(n_294), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_249), .A2(n_275), .B1(n_355), .B2(n_358), .C(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g280 ( .A(n_250), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g326 ( .A(n_250), .B(n_281), .Y(n_326) );
OAI221xp5_ASAP7_75t_SL g251 ( .A1(n_252), .A2(n_255), .B1(n_258), .B2(n_262), .C(n_265), .Y(n_251) );
AND2x2_ASAP7_75t_L g397 ( .A(n_252), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g264 ( .A(n_253), .Y(n_264) );
INVx1_ASAP7_75t_L g350 ( .A(n_254), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_255), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g269 ( .A(n_257), .B(n_260), .Y(n_269) );
AND2x2_ASAP7_75t_L g345 ( .A(n_257), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g270 ( .A(n_264), .B(n_271), .Y(n_270) );
OAI21xp5_ASAP7_75t_SL g265 ( .A1(n_266), .A2(n_269), .B(n_270), .Y(n_265) );
INVx1_ASAP7_75t_L g389 ( .A(n_266), .Y(n_389) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x2_ASAP7_75t_L g368 ( .A(n_267), .B(n_295), .Y(n_368) );
AND2x2_ASAP7_75t_SL g341 ( .A(n_268), .B(n_277), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B(n_279), .Y(n_272) );
OAI22xp33_ASAP7_75t_L g309 ( .A1(n_273), .A2(n_307), .B1(n_310), .B2(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g379 ( .A(n_273), .Y(n_379) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g299 ( .A(n_276), .Y(n_299) );
INVx1_ASAP7_75t_L g360 ( .A(n_278), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_280), .B(n_282), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_280), .B(n_350), .Y(n_401) );
AND2x2_ASAP7_75t_L g369 ( .A(n_281), .B(n_370), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g362 ( .A1(n_282), .A2(n_363), .B(n_366), .C(n_374), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_305), .Y(n_283) );
AOI322xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .A3(n_288), .B1(n_290), .B2(n_295), .C1(n_296), .C2(n_304), .Y(n_284) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_286), .Y(n_402) );
AND2x2_ASAP7_75t_L g352 ( .A(n_287), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g386 ( .A(n_287), .Y(n_386) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_SL g337 ( .A(n_289), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_SL g343 ( .A(n_289), .B(n_335), .Y(n_343) );
AND2x2_ASAP7_75t_L g367 ( .A(n_289), .B(n_333), .Y(n_367) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g339 ( .A(n_293), .Y(n_339) );
NAND2xp33_ASAP7_75t_SL g296 ( .A(n_297), .B(n_302), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI221xp5_ASAP7_75t_SL g342 ( .A1(n_298), .A2(n_343), .B1(n_344), .B2(n_345), .C(n_347), .Y(n_342) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVxp67_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g409 ( .A(n_301), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_308), .B(n_309), .C(n_313), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g384 ( .A(n_308), .Y(n_384) );
INVx1_ASAP7_75t_L g316 ( .A(n_310), .Y(n_316) );
OR2x2_ASAP7_75t_L g403 ( .A(n_310), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_SL g399 ( .A(n_311), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_317), .B(n_319), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_315), .B(n_333), .Y(n_410) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_342), .Y(n_321) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_325), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
OR2x2_ASAP7_75t_L g376 ( .A(n_329), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI21xp33_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_339), .B(n_340), .Y(n_336) );
INVx2_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AOI31xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_351), .A3(n_354), .B(n_356), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_353), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_379), .B2(n_380), .C(n_383), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_387), .B2(n_389), .Y(n_383) );
CKINVDCx16_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
NOR3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_400), .C(n_407), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_392), .B(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_399), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g415 ( .A(n_411), .Y(n_415) );
OAI22x1_ASAP7_75t_L g439 ( .A1(n_414), .A2(n_440), .B1(n_444), .B2(n_447), .Y(n_439) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_417), .Y(n_428) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g781 ( .A(n_418), .Y(n_781) );
BUFx2_ASAP7_75t_L g788 ( .A(n_418), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
AND2x6_ASAP7_75t_SL g443 ( .A(n_419), .B(n_421), .Y(n_443) );
OR2x6_ASAP7_75t_SL g446 ( .A(n_419), .B(n_420), .Y(n_446) );
OR2x2_ASAP7_75t_L g775 ( .A(n_419), .B(n_421), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g425 ( .A(n_426), .B(n_429), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_SL g433 ( .A(n_434), .B(n_436), .Y(n_433) );
INVx2_ASAP7_75t_L g780 ( .A(n_434), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_434), .A2(n_784), .B(n_787), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g779 ( .A(n_436), .B(n_780), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_767), .B(n_770), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
CKINVDCx11_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
CKINVDCx6p67_ASAP7_75t_R g773 ( .A(n_441), .Y(n_773) );
INVx3_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g772 ( .A(n_445), .Y(n_772) );
CKINVDCx11_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_657), .C(n_722), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_611), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_558), .B(n_584), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_522), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_474), .Y(n_453) );
AOI21xp33_ASAP7_75t_L g658 ( .A1(n_454), .A2(n_659), .B(n_670), .Y(n_658) );
AND2x2_ASAP7_75t_SL g693 ( .A(n_454), .B(n_600), .Y(n_693) );
AND2x2_ASAP7_75t_L g708 ( .A(n_454), .B(n_709), .Y(n_708) );
OR2x6_ASAP7_75t_L g718 ( .A(n_454), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g720 ( .A(n_454), .B(n_710), .Y(n_720) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g594 ( .A(n_455), .Y(n_594) );
AND2x2_ASAP7_75t_L g607 ( .A(n_455), .B(n_608), .Y(n_607) );
INVx4_ASAP7_75t_L g626 ( .A(n_455), .Y(n_626) );
AND2x2_ASAP7_75t_L g629 ( .A(n_455), .B(n_547), .Y(n_629) );
NOR2x1_ASAP7_75t_SL g632 ( .A(n_455), .B(n_562), .Y(n_632) );
AND2x4_ASAP7_75t_L g644 ( .A(n_455), .B(n_642), .Y(n_644) );
OR2x2_ASAP7_75t_L g654 ( .A(n_455), .B(n_529), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_455), .B(n_666), .Y(n_671) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVxp67_ASAP7_75t_L g497 ( .A(n_459), .Y(n_497) );
NOR2x1p5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g510 ( .A(n_462), .Y(n_510) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x6_ASAP7_75t_L g466 ( .A(n_463), .B(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_L g487 ( .A(n_466), .Y(n_487) );
INVx2_ASAP7_75t_L g557 ( .A(n_466), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_466), .A2(n_490), .B1(n_566), .B2(n_567), .Y(n_565) );
AND2x2_ASAP7_75t_L g471 ( .A(n_467), .B(n_472), .Y(n_471) );
INVxp33_ASAP7_75t_L g509 ( .A(n_467), .Y(n_509) );
INVx1_ASAP7_75t_L g499 ( .A(n_470), .Y(n_499) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g550 ( .A(n_471), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_473), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_474), .A2(n_600), .B1(n_695), .B2(n_696), .Y(n_694) );
INVx1_ASAP7_75t_SL g738 ( .A(n_474), .Y(n_738) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_500), .Y(n_474) );
INVx2_ASAP7_75t_L g669 ( .A(n_475), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_475), .B(n_615), .Y(n_741) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_483), .Y(n_475) );
BUFx3_ASAP7_75t_L g587 ( .A(n_476), .Y(n_587) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g580 ( .A(n_477), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_477), .B(n_502), .Y(n_602) );
AND2x4_ASAP7_75t_L g619 ( .A(n_477), .B(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_L g635 ( .A(n_477), .Y(n_635) );
INVx2_ASAP7_75t_L g692 ( .A(n_477), .Y(n_692) );
AND2x2_ASAP7_75t_L g610 ( .A(n_483), .B(n_576), .Y(n_610) );
NOR2xp67_ASAP7_75t_L g656 ( .A(n_483), .B(n_579), .Y(n_656) );
AND2x2_ASAP7_75t_L g675 ( .A(n_483), .B(n_579), .Y(n_675) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g539 ( .A(n_484), .Y(n_539) );
INVx1_ASAP7_75t_L g618 ( .A(n_484), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_484), .B(n_514), .Y(n_637) );
AND2x4_ASAP7_75t_L g691 ( .A(n_484), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g650 ( .A(n_500), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_500), .B(n_708), .Y(n_707) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_513), .Y(n_500) );
AND2x2_ASAP7_75t_L g634 ( .A(n_501), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g674 ( .A(n_501), .Y(n_674) );
AND2x2_ASAP7_75t_L g679 ( .A(n_501), .B(n_579), .Y(n_679) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_502), .B(n_514), .Y(n_541) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_512), .Y(n_502) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_503), .A2(n_504), .B(n_512), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_505), .B(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g615 ( .A(n_513), .Y(n_615) );
NAND2x1p5_ASAP7_75t_L g733 ( .A(n_513), .B(n_587), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_513), .B(n_539), .Y(n_754) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_514), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
OAI21xp33_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_537), .B(n_542), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_525), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g592 ( .A(n_526), .Y(n_592) );
AND2x2_ASAP7_75t_L g606 ( .A(n_526), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g640 ( .A(n_526), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g706 ( .A(n_526), .B(n_624), .Y(n_706) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_526), .B(n_753), .C(n_754), .Y(n_752) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_527), .Y(n_583) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g599 ( .A(n_529), .Y(n_599) );
AND2x2_ASAP7_75t_L g605 ( .A(n_529), .B(n_562), .Y(n_605) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_529), .Y(n_616) );
AND2x2_ASAP7_75t_L g661 ( .A(n_529), .B(n_561), .Y(n_661) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_529), .Y(n_684) );
INVx1_ASAP7_75t_L g701 ( .A(n_529), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g743 ( .A(n_537), .Y(n_743) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_538), .B(n_614), .Y(n_715) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g577 ( .A(n_539), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AOI211x1_ASAP7_75t_L g611 ( .A1(n_543), .A2(n_612), .B(n_621), .C(n_638), .Y(n_611) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_544), .B(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g664 ( .A(n_544), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g600 ( .A(n_546), .B(n_561), .Y(n_600) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g560 ( .A(n_547), .B(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_547), .Y(n_625) );
INVx1_ASAP7_75t_L g642 ( .A(n_547), .Y(n_642) );
AND2x2_ASAP7_75t_L g710 ( .A(n_547), .B(n_562), .Y(n_710) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_553), .Y(n_547) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .C(n_552), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_574), .B(n_581), .Y(n_558) );
NOR2x1_ASAP7_75t_L g729 ( .A(n_559), .B(n_626), .Y(n_729) );
INVx2_ASAP7_75t_L g761 ( .A(n_559), .Y(n_761) );
INVx4_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g593 ( .A(n_560), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g666 ( .A(n_561), .Y(n_666) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .B(n_573), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_571), .B2(n_572), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
OR2x2_ASAP7_75t_L g668 ( .A(n_575), .B(n_669), .Y(n_668) );
NAND2x1_ASAP7_75t_SL g690 ( .A(n_575), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x4_ASAP7_75t_L g590 ( .A(n_576), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g620 ( .A(n_576), .Y(n_620) );
INVx1_ASAP7_75t_L g744 ( .A(n_577), .Y(n_744) );
AND2x2_ASAP7_75t_L g609 ( .A(n_578), .B(n_610), .Y(n_609) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx2_ASAP7_75t_L g591 ( .A(n_579), .Y(n_591) );
INVxp33_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g648 ( .A(n_583), .B(n_641), .Y(n_648) );
OAI211xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_588), .B(n_595), .C(n_603), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g672 ( .A(n_586), .B(n_673), .Y(n_672) );
NOR2xp67_ASAP7_75t_SL g677 ( .A(n_586), .B(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_587), .B(n_674), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_589), .B(n_593), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
AND2x2_ASAP7_75t_L g721 ( .A(n_590), .B(n_691), .Y(n_721) );
AOI222xp33_ASAP7_75t_L g739 ( .A1(n_593), .A2(n_740), .B1(n_742), .B2(n_745), .C1(n_746), .C2(n_749), .Y(n_739) );
INVx1_ASAP7_75t_L g703 ( .A(n_594), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_601), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_599), .Y(n_630) );
AND2x4_ASAP7_75t_SL g665 ( .A(n_599), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g719 ( .A(n_600), .Y(n_719) );
AND2x2_ASAP7_75t_L g764 ( .A(n_600), .B(n_616), .Y(n_764) );
AND2x2_ASAP7_75t_L g645 ( .A(n_601), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g758 ( .A(n_602), .B(n_637), .Y(n_758) );
OAI21xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_606), .B(n_609), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_604), .A2(n_624), .B(n_665), .Y(n_725) );
AND2x2_ASAP7_75t_L g749 ( .A(n_605), .B(n_626), .Y(n_749) );
NOR2xp33_ASAP7_75t_SL g759 ( .A(n_605), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g697 ( .A(n_608), .Y(n_697) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_608), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g732 ( .A(n_610), .Y(n_732) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_617), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g735 ( .A(n_615), .B(n_619), .Y(n_735) );
BUFx2_ASAP7_75t_L g623 ( .A(n_616), .Y(n_623) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g646 ( .A(n_618), .Y(n_646) );
INVx2_ASAP7_75t_L g652 ( .A(n_618), .Y(n_652) );
AND2x2_ASAP7_75t_L g688 ( .A(n_618), .B(n_679), .Y(n_688) );
AND2x4_ASAP7_75t_L g655 ( .A(n_619), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g695 ( .A(n_619), .B(n_652), .Y(n_695) );
AND2x2_ASAP7_75t_L g746 ( .A(n_619), .B(n_747), .Y(n_746) );
AOI31xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_627), .A3(n_631), .B(n_633), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g643 ( .A(n_623), .B(n_644), .Y(n_643) );
AND2x4_ASAP7_75t_SL g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x4_ASAP7_75t_L g641 ( .A(n_626), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_629), .A2(n_681), .B1(n_712), .B2(n_715), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_629), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g766 ( .A(n_629), .B(n_682), .Y(n_766) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g681 ( .A(n_632), .B(n_682), .Y(n_681) );
NAND2x1p5_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
AND2x2_ASAP7_75t_L g704 ( .A(n_634), .B(n_675), .Y(n_704) );
INVx1_ASAP7_75t_L g714 ( .A(n_636), .Y(n_714) );
INVx2_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_647), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B(n_645), .Y(n_639) );
INVx1_ASAP7_75t_L g737 ( .A(n_640), .Y(n_737) );
AND2x2_ASAP7_75t_L g745 ( .A(n_641), .B(n_697), .Y(n_745) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_641), .Y(n_751) );
AND2x2_ASAP7_75t_L g696 ( .A(n_644), .B(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_649), .B1(n_653), .B2(n_655), .Y(n_647) );
NOR2xp33_ASAP7_75t_SL g649 ( .A(n_650), .B(n_651), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_650), .A2(n_669), .B1(n_763), .B2(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g662 ( .A(n_655), .Y(n_662) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_685), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B(n_663), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
OAI21xp33_ASAP7_75t_L g663 ( .A1(n_661), .A2(n_664), .B(n_667), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_664), .A2(n_688), .B1(n_689), .B2(n_693), .Y(n_687) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B1(n_676), .B2(n_680), .Y(n_670) );
INVx1_ASAP7_75t_L g705 ( .A(n_673), .Y(n_705) );
NAND2x1p5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_686), .B(n_698), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_694), .Y(n_686) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
NAND2xp33_ASAP7_75t_SL g740 ( .A(n_690), .B(n_741), .Y(n_740) );
INVx3_ASAP7_75t_L g713 ( .A(n_691), .Y(n_713) );
INVx3_ASAP7_75t_L g727 ( .A(n_695), .Y(n_727) );
INVxp67_ASAP7_75t_L g756 ( .A(n_696), .Y(n_756) );
NAND4xp25_ASAP7_75t_L g698 ( .A(n_699), .B(n_707), .C(n_711), .D(n_716), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
AND2x2_ASAP7_75t_L g709 ( .A(n_701), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g757 ( .A(n_705), .Y(n_757) );
NAND2xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_714), .Y(n_712) );
OAI21xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_720), .B(n_721), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND3x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_739), .C(n_750), .Y(n_722) );
AOI221x1_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_726), .B1(n_728), .B2(n_730), .C(n_736), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp33_ASAP7_75t_SL g730 ( .A(n_731), .B(n_734), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
NAND2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI211xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B(n_755), .C(n_762), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_755) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx4f_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_781), .Y(n_777) );
INVxp67_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
CKINVDCx11_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
CKINVDCx8_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
endmodule