module fake_jpeg_14049_n_649 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_649);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_649;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_59),
.Y(n_170)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_60),
.Y(n_158)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx2_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_62),
.B(n_63),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_67),
.B(n_68),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_71),
.B(n_81),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_79),
.Y(n_164)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_80),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_85),
.Y(n_182)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_87),
.B(n_98),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_18),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_88),
.B(n_95),
.Y(n_157)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_89),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_91),
.B(n_45),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_26),
.B(n_18),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_35),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g176 ( 
.A(n_97),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_34),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_101),
.A2(n_42),
.B1(n_55),
.B2(n_54),
.Y(n_212)
);

BUFx16f_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_25),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_105),
.B(n_109),
.Y(n_192)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_51),
.Y(n_107)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_34),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_36),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_111),
.B(n_122),
.Y(n_195)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_113),
.Y(n_211)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_37),
.Y(n_119)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_48),
.Y(n_120)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_40),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_124),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_26),
.B(n_18),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_41),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_47),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_128),
.B(n_54),
.Y(n_203)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_50),
.Y(n_129)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_58),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_130),
.B(n_149),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_46),
.B1(n_22),
.B2(n_49),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_133),
.A2(n_161),
.B1(n_77),
.B2(n_99),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_80),
.B(n_58),
.C(n_56),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_143),
.B(n_4),
.C(n_5),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_113),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_62),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_152),
.B(n_155),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_101),
.Y(n_155)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_166),
.B(n_6),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_168),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_69),
.B(n_45),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_175),
.B(n_184),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_93),
.A2(n_50),
.B1(n_46),
.B2(n_22),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_177),
.A2(n_22),
.B1(n_46),
.B2(n_104),
.Y(n_229)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_178),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_179),
.B(n_181),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_38),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_102),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_129),
.B(n_38),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_193),
.B(n_205),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_107),
.A2(n_32),
.B(n_55),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_200),
.B(n_6),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_203),
.B(n_215),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_60),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_102),
.B(n_42),
.Y(n_205)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_61),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_86),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_52),
.B1(n_43),
.B2(n_32),
.Y(n_241)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_94),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_115),
.Y(n_216)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_96),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_217),
.B(n_219),
.Y(n_295)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_59),
.B(n_52),
.Y(n_219)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_65),
.Y(n_220)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_195),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_222),
.B(n_224),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_163),
.A2(n_75),
.B1(n_121),
.B2(n_73),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g325 ( 
.A1(n_223),
.A2(n_228),
.B1(n_230),
.B2(n_233),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_135),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_225),
.B(n_245),
.Y(n_314)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_227),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_229),
.A2(n_232),
.B1(n_246),
.B2(n_279),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_163),
.A2(n_72),
.B1(n_108),
.B2(n_85),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_152),
.A2(n_82),
.B1(n_70),
.B2(n_118),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_172),
.A2(n_194),
.B1(n_165),
.B2(n_173),
.Y(n_233)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_145),
.Y(n_237)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_237),
.Y(n_340)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_134),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_239),
.Y(n_359)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_139),
.Y(n_240)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_240),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_241),
.A2(n_289),
.B1(n_211),
.B2(n_137),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_187),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_157),
.A2(n_66),
.B1(n_126),
.B2(n_118),
.Y(n_246)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

INVx4_ASAP7_75t_SL g321 ( 
.A(n_249),
.Y(n_321)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_145),
.Y(n_250)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_146),
.Y(n_252)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_253),
.Y(n_350)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_255),
.Y(n_332)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_256),
.Y(n_338)
);

INVx4_ASAP7_75t_SL g257 ( 
.A(n_176),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_281),
.Y(n_300)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_142),
.Y(n_258)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_170),
.Y(n_259)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_259),
.Y(n_305)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_144),
.Y(n_260)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_160),
.Y(n_261)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_135),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_262),
.Y(n_349)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_188),
.Y(n_264)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_264),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_265),
.Y(n_347)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_268),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_159),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_269),
.B(n_274),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_172),
.A2(n_56),
.B1(n_47),
.B2(n_120),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_270),
.A2(n_272),
.B1(n_190),
.B2(n_158),
.Y(n_302)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_206),
.Y(n_271)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_271),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_194),
.A2(n_120),
.B1(n_126),
.B2(n_3),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_150),
.Y(n_273)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_164),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_132),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_275),
.B(n_278),
.Y(n_331)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_133),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_170),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_280),
.B(n_282),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_180),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_169),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_283),
.B(n_285),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g284 ( 
.A(n_131),
.B(n_130),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_284),
.B(n_292),
.Y(n_303)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_197),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_185),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_286),
.B(n_287),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_180),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_196),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_290),
.B(n_291),
.Y(n_356)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_201),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_204),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_294),
.B1(n_132),
.B2(n_168),
.Y(n_306)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_154),
.Y(n_294)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_202),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_298),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_297),
.A2(n_7),
.B(n_10),
.Y(n_339)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_189),
.Y(n_298)
);

INVx6_ASAP7_75t_SL g299 ( 
.A(n_180),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_299),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_248),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_306),
.A2(n_311),
.B1(n_312),
.B2(n_334),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_263),
.A2(n_297),
.B1(n_236),
.B2(n_230),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_307),
.B(n_315),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_309),
.B(n_320),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_247),
.A2(n_220),
.B1(n_190),
.B2(n_214),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_310),
.A2(n_336),
.B1(n_344),
.B2(n_242),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_279),
.A2(n_174),
.B1(n_136),
.B2(n_141),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_228),
.A2(n_174),
.B1(n_136),
.B2(n_141),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_267),
.B(n_214),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_284),
.A2(n_148),
.A3(n_211),
.B1(n_178),
.B2(n_209),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_226),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_277),
.B(n_292),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_319),
.B(n_339),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_295),
.B(n_210),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_231),
.B(n_151),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_329),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_151),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_232),
.A2(n_158),
.B1(n_140),
.B2(n_171),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_223),
.A2(n_198),
.B1(n_182),
.B2(n_154),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_335),
.A2(n_353),
.B1(n_239),
.B2(n_227),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_270),
.A2(n_182),
.B1(n_198),
.B2(n_140),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_243),
.B(n_147),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_342),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_254),
.B(n_138),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_272),
.A2(n_191),
.B1(n_156),
.B2(n_162),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_346),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_233),
.A2(n_162),
.B1(n_186),
.B2(n_183),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_235),
.B(n_10),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_293),
.A2(n_186),
.B1(n_153),
.B2(n_12),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_257),
.B(n_10),
.Y(n_355)
);

XNOR2x1_ASAP7_75t_SL g406 ( 
.A(n_355),
.B(n_323),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_226),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_357)
);

INVx4_ASAP7_75t_SL g386 ( 
.A(n_357),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_362),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_354),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_364),
.B(n_382),
.Y(n_416)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_365),
.Y(n_439)
);

MAJx2_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_234),
.C(n_276),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_366),
.B(n_376),
.C(n_381),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_355),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_368),
.B(n_373),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_339),
.A2(n_262),
.B(n_242),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_369),
.A2(n_380),
.B(n_388),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_327),
.A2(n_294),
.B1(n_256),
.B2(n_240),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_370),
.A2(n_371),
.B1(n_401),
.B2(n_343),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_244),
.Y(n_373)
);

INVx13_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_374),
.A2(n_377),
.B1(n_395),
.B2(n_405),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_375),
.A2(n_349),
.B1(n_358),
.B2(n_347),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_300),
.B(n_268),
.C(n_249),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_335),
.A2(n_252),
.B1(n_273),
.B2(n_265),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_320),
.B(n_244),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_379),
.B(n_387),
.Y(n_419)
);

AO22x1_ASAP7_75t_L g380 ( 
.A1(n_325),
.A2(n_266),
.B1(n_248),
.B2(n_259),
.Y(n_380)
);

MAJx2_ASAP7_75t_L g381 ( 
.A(n_300),
.B(n_238),
.C(n_266),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_348),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_316),
.B(n_253),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_398),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_300),
.B(n_251),
.C(n_280),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_399),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_330),
.B(n_275),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_327),
.A2(n_275),
.B(n_13),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_303),
.B(n_11),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_391),
.B(n_396),
.Y(n_431)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_317),
.Y(n_393)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_393),
.Y(n_423)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_301),
.Y(n_394)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

INVx13_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_355),
.Y(n_396)
);

NAND2x1_ASAP7_75t_L g397 ( 
.A(n_329),
.B(n_11),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_397),
.A2(n_404),
.B(n_331),
.Y(n_433)
);

AND2x6_ASAP7_75t_L g398 ( 
.A(n_303),
.B(n_17),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_307),
.B(n_17),
.C(n_301),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_346),
.B(n_17),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_356),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_325),
.A2(n_319),
.B1(n_302),
.B2(n_342),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

FAx1_ASAP7_75t_L g404 ( 
.A(n_353),
.B(n_326),
.CI(n_341),
.CON(n_404),
.SN(n_404)
);

INVx13_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_406),
.B(n_345),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_414),
.A2(n_403),
.B1(n_383),
.B2(n_404),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_364),
.B(n_314),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_415),
.B(n_420),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_417),
.B(n_421),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_382),
.B(n_333),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_337),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_337),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_422),
.B(n_438),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_371),
.Y(n_462)
);

XOR2x2_ASAP7_75t_L g429 ( 
.A(n_361),
.B(n_323),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_397),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_361),
.B(n_366),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_430),
.B(n_445),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_401),
.A2(n_318),
.B1(n_338),
.B2(n_347),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_432),
.A2(n_434),
.B1(n_435),
.B2(n_441),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_433),
.A2(n_385),
.B(n_406),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_370),
.A2(n_358),
.B1(n_351),
.B2(n_324),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_389),
.A2(n_351),
.B1(n_324),
.B2(n_322),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_376),
.A2(n_349),
.B1(n_305),
.B2(n_350),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_436),
.A2(n_369),
.B(n_397),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_388),
.A2(n_322),
.B1(n_308),
.B2(n_359),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_363),
.B(n_323),
.Y(n_440)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_440),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_389),
.A2(n_359),
.B1(n_308),
.B2(n_352),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_372),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_442),
.B(n_396),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_378),
.B(n_352),
.Y(n_443)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_443),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_400),
.B(n_372),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_444),
.B(n_398),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_447),
.B(n_448),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_304),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_420),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_440),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_304),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_450),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_416),
.B(n_402),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_451),
.B(n_455),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_454),
.A2(n_476),
.B(n_479),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_421),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_305),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_456),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_435),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_459),
.B(n_470),
.Y(n_495)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_424),
.Y(n_460)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_407),
.B(n_381),
.C(n_368),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_461),
.B(n_464),
.C(n_478),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_462),
.A2(n_465),
.B1(n_480),
.B2(n_429),
.Y(n_493)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_463),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_378),
.C(n_394),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_430),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_428),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_469),
.Y(n_483)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_428),
.Y(n_468)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_468),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_439),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_417),
.B(n_431),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_471),
.A2(n_436),
.B(n_438),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_472),
.B(n_433),
.Y(n_485)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_410),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_474),
.B(n_423),
.Y(n_513)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_443),
.Y(n_475)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_475),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_418),
.B(n_384),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_477),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_345),
.C(n_405),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_426),
.B(n_371),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_411),
.A2(n_404),
.B1(n_380),
.B2(n_386),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_455),
.A2(n_414),
.B1(n_411),
.B2(n_432),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_484),
.A2(n_490),
.B1(n_501),
.B2(n_512),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_500),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_487),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_458),
.B(n_409),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g535 ( 
.A(n_488),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_479),
.A2(n_426),
.B(n_429),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_SL g528 ( 
.A1(n_489),
.A2(n_476),
.B(n_463),
.C(n_468),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_477),
.A2(n_408),
.B1(n_409),
.B2(n_441),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_480),
.A2(n_465),
.B1(n_479),
.B2(n_462),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_492),
.A2(n_493),
.B1(n_478),
.B2(n_461),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_457),
.B(n_446),
.Y(n_496)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_496),
.Y(n_519)
);

AOI21xp33_ASAP7_75t_L g544 ( 
.A1(n_499),
.A2(n_510),
.B(n_367),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_473),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_446),
.A2(n_408),
.B1(n_425),
.B2(n_434),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_502),
.B(n_413),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_458),
.B(n_412),
.Y(n_503)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_503),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_457),
.B(n_475),
.Y(n_505)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_505),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_453),
.B(n_412),
.Y(n_506)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_506),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_453),
.B(n_472),
.Y(n_509)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_509),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_R g510 ( 
.A1(n_454),
.A2(n_380),
.B1(n_439),
.B2(n_386),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_459),
.A2(n_413),
.B1(n_427),
.B2(n_423),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_513),
.B(n_460),
.Y(n_527)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_473),
.Y(n_515)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_515),
.Y(n_529)
);

AOI21x1_ASAP7_75t_L g516 ( 
.A1(n_498),
.A2(n_471),
.B(n_462),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_516),
.A2(n_528),
.B(n_544),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_483),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_520),
.B(n_484),
.Y(n_550)
);

XNOR2x1_ASAP7_75t_L g569 ( 
.A(n_522),
.B(n_501),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_464),
.C(n_481),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_523),
.B(n_526),
.C(n_530),
.Y(n_547)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_510),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_524),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_492),
.A2(n_493),
.B1(n_515),
.B2(n_500),
.Y(n_525)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_525),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_481),
.C(n_466),
.Y(n_526)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_527),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_467),
.C(n_452),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_502),
.B(n_467),
.C(n_452),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_537),
.C(n_540),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_534),
.B(n_505),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_495),
.A2(n_469),
.B1(n_386),
.B2(n_437),
.Y(n_536)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_536),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_437),
.C(n_340),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_489),
.B(n_340),
.C(n_362),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_498),
.B(n_332),
.C(n_308),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_541),
.B(n_545),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_514),
.Y(n_542)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_495),
.B(n_496),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_543),
.B(n_522),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_499),
.A2(n_365),
.B(n_374),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_529),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_549),
.B(n_568),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_550),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_485),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_552),
.B(n_561),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_488),
.Y(n_554)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_554),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_517),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_555),
.B(n_558),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_530),
.B(n_507),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_535),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_559),
.B(n_543),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_523),
.B(n_534),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_519),
.Y(n_562)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_562),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_564),
.B(n_565),
.Y(n_587)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_531),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_566),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_533),
.A2(n_509),
.B1(n_511),
.B2(n_497),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_567),
.A2(n_570),
.B1(n_536),
.B2(n_512),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_520),
.B(n_491),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_541),
.C(n_525),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_533),
.A2(n_511),
.B1(n_497),
.B2(n_491),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_554),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_572),
.B(n_575),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_529),
.Y(n_573)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_573),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_551),
.A2(n_524),
.B1(n_518),
.B2(n_504),
.Y(n_574)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_574),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_557),
.B(n_507),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_576),
.A2(n_590),
.B1(n_560),
.B2(n_546),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_547),
.B(n_526),
.C(n_537),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_582),
.B(n_590),
.C(n_553),
.Y(n_594)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_583),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_563),
.A2(n_516),
.B(n_545),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_585),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g585 ( 
.A1(n_560),
.A2(n_528),
.B(n_483),
.C(n_521),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_586),
.B(n_569),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_567),
.A2(n_513),
.B1(n_494),
.B2(n_482),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_589),
.B(n_565),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_547),
.B(n_528),
.C(n_540),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_SL g616 ( 
.A(n_592),
.B(n_581),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_594),
.B(n_600),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_582),
.B(n_553),
.C(n_564),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_596),
.B(n_599),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_605),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_578),
.B(n_552),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_571),
.A2(n_556),
.B(n_568),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_578),
.B(n_548),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g620 ( 
.A(n_601),
.B(n_607),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_579),
.A2(n_570),
.B1(n_546),
.B2(n_550),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_602),
.A2(n_579),
.B1(n_577),
.B2(n_584),
.Y(n_615)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_604),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_576),
.B(n_563),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_561),
.C(n_573),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_606),
.B(n_490),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_580),
.B(n_538),
.Y(n_607)
);

INVx11_ASAP7_75t_L g610 ( 
.A(n_597),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_610),
.A2(n_585),
.B1(n_528),
.B2(n_486),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_594),
.B(n_573),
.C(n_587),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_612),
.B(n_614),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_603),
.B(n_588),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_615),
.B(n_617),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_616),
.B(n_608),
.C(n_612),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_599),
.B(n_596),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_602),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_618),
.B(n_621),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_593),
.A2(n_581),
.B(n_577),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_619),
.A2(n_595),
.B(n_482),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_617),
.B(n_605),
.Y(n_624)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_624),
.Y(n_633)
);

XNOR2x1_ASAP7_75t_L g638 ( 
.A(n_625),
.B(n_626),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_611),
.B(n_598),
.C(n_606),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_609),
.B(n_588),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_628),
.A2(n_631),
.B(n_620),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_610),
.B(n_591),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_629),
.B(n_630),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_622),
.B(n_613),
.Y(n_634)
);

AOI21x1_ASAP7_75t_L g640 ( 
.A1(n_634),
.A2(n_635),
.B(n_636),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_626),
.A2(n_608),
.B(n_619),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_627),
.B(n_616),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_637),
.B(n_623),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_639),
.B(n_641),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_632),
.Y(n_641)
);

A2O1A1O1Ixp25_ASAP7_75t_L g642 ( 
.A1(n_633),
.A2(n_638),
.B(n_630),
.C(n_595),
.D(n_592),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_642),
.B(n_486),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_644),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_643),
.B(n_640),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_494),
.C(n_395),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_359),
.C(n_332),
.Y(n_648)
);

AO21x1_ASAP7_75t_L g649 ( 
.A1(n_648),
.A2(n_392),
.B(n_393),
.Y(n_649)
);


endmodule