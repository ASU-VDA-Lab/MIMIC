module fake_aes_2000_n_1322 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1322);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1322;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_315;
wire n_1321;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_659;
wire n_432;
wire n_386;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVxp33_ASAP7_75t_SL g298 ( .A(n_133), .Y(n_298) );
INVxp33_ASAP7_75t_SL g299 ( .A(n_246), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_6), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_36), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_198), .Y(n_302) );
INVxp33_ASAP7_75t_L g303 ( .A(n_46), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_130), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_226), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_154), .Y(n_306) );
INVxp33_ASAP7_75t_L g307 ( .A(n_192), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_191), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_60), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_168), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_235), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_227), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_179), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_228), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_221), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_266), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_26), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_193), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_101), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_219), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_180), .Y(n_321) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_188), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_14), .Y(n_323) );
INVxp33_ASAP7_75t_SL g324 ( .A(n_217), .Y(n_324) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_251), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_14), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_105), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_290), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_248), .Y(n_329) );
INVxp33_ASAP7_75t_SL g330 ( .A(n_146), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_112), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_209), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_284), .Y(n_333) );
INVxp67_ASAP7_75t_SL g334 ( .A(n_166), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_136), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_280), .Y(n_336) );
INVxp33_ASAP7_75t_L g337 ( .A(n_19), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_19), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_72), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_296), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_157), .Y(n_341) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_102), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_85), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_247), .Y(n_344) );
INVxp33_ASAP7_75t_SL g345 ( .A(n_60), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_21), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_208), .Y(n_347) );
INVxp33_ASAP7_75t_SL g348 ( .A(n_205), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_176), .Y(n_349) );
INVxp33_ASAP7_75t_L g350 ( .A(n_195), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_77), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_262), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_223), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_218), .Y(n_354) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_82), .Y(n_355) );
INVxp67_ASAP7_75t_SL g356 ( .A(n_68), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_12), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_182), .Y(n_358) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_242), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_25), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_39), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_85), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_143), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_45), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_186), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_270), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_261), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_129), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_31), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_34), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_260), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_288), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_265), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_121), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_12), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_8), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_71), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_152), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_170), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_51), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_109), .Y(n_381) );
INVxp33_ASAP7_75t_L g382 ( .A(n_89), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_120), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_137), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_139), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_155), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_216), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_225), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_256), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_250), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_241), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_210), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_8), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_30), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_167), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_275), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_103), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_214), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_25), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_57), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_293), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_96), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_272), .Y(n_403) );
INVxp33_ASAP7_75t_L g404 ( .A(n_172), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_92), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_50), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_5), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_230), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_29), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_259), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_285), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_88), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_80), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_56), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_255), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_100), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_57), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_159), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_33), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_183), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_281), .Y(n_421) );
CKINVDCx14_ASAP7_75t_R g422 ( .A(n_91), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_61), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_76), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_138), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_211), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_111), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_158), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_239), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_237), .Y(n_430) );
INVxp33_ASAP7_75t_SL g431 ( .A(n_144), .Y(n_431) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_276), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_273), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_149), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_20), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_134), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_55), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_40), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_156), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_95), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_86), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_22), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_37), .B(n_201), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_61), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_113), .Y(n_445) );
OAI21x1_ASAP7_75t_L g446 ( .A1(n_402), .A2(n_93), .B(n_90), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_310), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_333), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_310), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_327), .Y(n_450) );
NOR2x1_ASAP7_75t_L g451 ( .A(n_362), .B(n_0), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_327), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_336), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_407), .B(n_0), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_407), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_336), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_340), .Y(n_457) );
AND3x2_ASAP7_75t_L g458 ( .A(n_429), .B(n_1), .C(n_2), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_340), .Y(n_459) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_362), .B(n_1), .Y(n_460) );
NAND2x1_ASAP7_75t_L g461 ( .A(n_402), .B(n_2), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_303), .B(n_337), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_341), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_326), .B(n_338), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_402), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_360), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_341), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_333), .Y(n_468) );
NOR2xp33_ASAP7_75t_SL g469 ( .A(n_391), .B(n_297), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_333), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_413), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_423), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_344), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_307), .B(n_3), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_333), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_360), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_301), .B(n_3), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_344), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_326), .B(n_4), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_472), .B(n_313), .Y(n_480) );
AND2x6_ASAP7_75t_L g481 ( .A(n_477), .B(n_347), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_465), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_477), .B(n_423), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_448), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_448), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_465), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_447), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_448), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_477), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_448), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_465), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_455), .B(n_408), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_477), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_472), .B(n_447), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_448), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_462), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_455), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_477), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_462), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_462), .B(n_422), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_471), .B(n_364), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_454), .B(n_301), .Y(n_502) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_448), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_449), .B(n_350), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_448), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_466), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_454), .B(n_376), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_448), .Y(n_508) );
INVx4_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_475), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_454), .B(n_376), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_449), .B(n_338), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_471), .B(n_382), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_450), .B(n_339), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_475), .Y(n_516) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_475), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_446), .Y(n_518) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_475), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_466), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_466), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_450), .B(n_339), .Y(n_522) );
INVx3_ASAP7_75t_L g523 ( .A(n_466), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_452), .B(n_313), .Y(n_524) );
BUFx3_ASAP7_75t_L g525 ( .A(n_446), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_446), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g527 ( .A(n_461), .B(n_443), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_494), .B(n_474), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_482), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_482), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_496), .B(n_464), .Y(n_531) );
OR2x6_ASAP7_75t_L g532 ( .A(n_509), .B(n_461), .Y(n_532) );
AOI22xp5_ASAP7_75t_SL g533 ( .A1(n_497), .A2(n_335), .B1(n_363), .B2(n_352), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_486), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_518), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_492), .Y(n_536) );
NAND3xp33_ASAP7_75t_SL g537 ( .A(n_496), .B(n_352), .C(n_335), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_512), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_518), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_502), .B(n_474), .Y(n_540) );
BUFx2_ASAP7_75t_L g541 ( .A(n_481), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_494), .B(n_474), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_504), .B(n_452), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_499), .A2(n_363), .B1(n_388), .B2(n_345), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_481), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_486), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_491), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_504), .B(n_453), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_489), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_499), .Y(n_550) );
AO22x1_ASAP7_75t_L g551 ( .A1(n_481), .A2(n_299), .B1(n_324), .B2(n_298), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_501), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_491), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_500), .B(n_453), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_489), .Y(n_555) );
INVxp67_ASAP7_75t_SL g556 ( .A(n_487), .Y(n_556) );
INVx3_ASAP7_75t_L g557 ( .A(n_489), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_500), .B(n_456), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_500), .B(n_464), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_489), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_512), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_481), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_502), .B(n_456), .Y(n_563) );
O2A1O1Ixp5_ASAP7_75t_L g564 ( .A1(n_489), .A2(n_461), .B(n_457), .C(n_459), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_502), .B(n_458), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_518), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_498), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_512), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_481), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_498), .Y(n_570) );
NOR2xp33_ASAP7_75t_R g571 ( .A(n_509), .B(n_469), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_498), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_501), .B(n_479), .Y(n_573) );
O2A1O1Ixp33_ASAP7_75t_L g574 ( .A1(n_493), .A2(n_479), .B(n_459), .C(n_463), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_498), .Y(n_575) );
AND3x2_ASAP7_75t_SL g576 ( .A(n_527), .B(n_469), .C(n_329), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_487), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_492), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_502), .B(n_457), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_487), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_512), .Y(n_581) );
BUFx6f_ASAP7_75t_SL g582 ( .A(n_509), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_492), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_501), .Y(n_584) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_480), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_481), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_481), .Y(n_587) );
AOI21x1_ASAP7_75t_L g588 ( .A1(n_520), .A2(n_467), .B(n_463), .Y(n_588) );
AO22x1_ASAP7_75t_L g589 ( .A1(n_481), .A2(n_299), .B1(n_324), .B2(n_298), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_506), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g591 ( .A(n_509), .B(n_443), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_513), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_502), .B(n_467), .Y(n_593) );
INVx2_ASAP7_75t_SL g594 ( .A(n_481), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_481), .A2(n_478), .B1(n_473), .B2(n_345), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_506), .Y(n_596) );
OR2x6_ASAP7_75t_L g597 ( .A(n_509), .B(n_451), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_507), .B(n_473), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_493), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_506), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_513), .B(n_478), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_507), .B(n_302), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_512), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_506), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_507), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_513), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_514), .Y(n_607) );
NOR2xp33_ASAP7_75t_R g608 ( .A(n_480), .B(n_388), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_507), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_507), .A2(n_309), .B1(n_393), .B2(n_346), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_506), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_523), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_511), .B(n_451), .Y(n_613) );
BUFx2_ASAP7_75t_R g614 ( .A(n_518), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_514), .Y(n_615) );
INVx5_ASAP7_75t_L g616 ( .A(n_523), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_527), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_523), .Y(n_618) );
NOR2x1p5_ASAP7_75t_SL g619 ( .A(n_520), .B(n_314), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_523), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_511), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_523), .Y(n_622) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_617), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_550), .B(n_511), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_601), .B(n_511), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_549), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_585), .B(n_511), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_535), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_552), .B(n_527), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_559), .A2(n_522), .B1(n_514), .B2(n_317), .C(n_361), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_584), .B(n_527), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_549), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_549), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_573), .B(n_540), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_556), .A2(n_526), .B(n_525), .Y(n_635) );
BUFx3_ASAP7_75t_L g636 ( .A(n_565), .Y(n_636) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_562), .B(n_514), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_592), .B(n_514), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_573), .B(n_522), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_555), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_607), .Y(n_641) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_532), .A2(n_524), .B1(n_442), .B2(n_343), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_536), .B(n_483), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_608), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_555), .Y(n_645) );
INVx4_ASAP7_75t_L g646 ( .A(n_582), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_607), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_601), .B(n_522), .Y(n_648) );
INVx4_ASAP7_75t_L g649 ( .A(n_582), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_541), .Y(n_650) );
OR2x6_ASAP7_75t_L g651 ( .A(n_544), .B(n_483), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_555), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_606), .B(n_522), .Y(n_653) );
INVxp67_ASAP7_75t_SL g654 ( .A(n_562), .Y(n_654) );
AOI22xp5_ASAP7_75t_SL g655 ( .A1(n_533), .A2(n_346), .B1(n_393), .B2(n_309), .Y(n_655) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_535), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_615), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_540), .B(n_522), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_531), .B(n_483), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_557), .Y(n_660) );
AOI21xp33_ASAP7_75t_L g661 ( .A1(n_574), .A2(n_526), .B(n_525), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_571), .Y(n_662) );
OAI21x1_ASAP7_75t_L g663 ( .A1(n_588), .A2(n_524), .B(n_488), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_606), .B(n_483), .Y(n_664) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_535), .Y(n_665) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_535), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_557), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_543), .A2(n_483), .B1(n_526), .B2(n_525), .Y(n_668) );
INVx3_ASAP7_75t_L g669 ( .A(n_557), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_565), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_578), .B(n_399), .Y(n_671) );
AND2x4_ASAP7_75t_L g672 ( .A(n_540), .B(n_460), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_613), .A2(n_525), .B1(n_526), .B2(n_460), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_583), .B(n_399), .Y(n_674) );
INVx4_ASAP7_75t_L g675 ( .A(n_582), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_577), .A2(n_521), .B(n_411), .Y(n_676) );
BUFx4f_ASAP7_75t_L g677 ( .A(n_565), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_564), .A2(n_347), .B(n_412), .C(n_411), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_613), .B(n_355), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_609), .A2(n_356), .B1(n_357), .B2(n_400), .C1(n_323), .C2(n_394), .Y(n_680) );
BUFx12f_ASAP7_75t_L g681 ( .A(n_532), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_615), .Y(n_682) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_535), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_591), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_560), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_613), .B(n_330), .Y(n_686) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_539), .Y(n_687) );
AND2x4_ASAP7_75t_L g688 ( .A(n_605), .B(n_351), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_560), .Y(n_689) );
NAND2x1p5_ASAP7_75t_L g690 ( .A(n_541), .B(n_343), .Y(n_690) );
INVx1_ASAP7_75t_SL g691 ( .A(n_621), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_560), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_599), .A2(n_445), .B(n_415), .C(n_370), .Y(n_693) );
BUFx10_ASAP7_75t_L g694 ( .A(n_532), .Y(n_694) );
BUFx3_ASAP7_75t_L g695 ( .A(n_591), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_605), .A2(n_538), .B1(n_568), .B2(n_561), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_610), .B(n_300), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_591), .B(n_406), .Y(n_698) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_537), .Y(n_699) );
INVxp67_ASAP7_75t_L g700 ( .A(n_602), .Y(n_700) );
INVx5_ASAP7_75t_L g701 ( .A(n_587), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_577), .A2(n_521), .B(n_325), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g703 ( .A1(n_554), .A2(n_348), .B1(n_431), .B2(n_330), .Y(n_703) );
BUFx4f_ASAP7_75t_L g704 ( .A(n_532), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_581), .B(n_348), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_548), .A2(n_375), .B(n_377), .C(n_369), .Y(n_706) );
BUFx2_ASAP7_75t_L g707 ( .A(n_551), .Y(n_707) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_539), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_528), .B(n_444), .Y(n_709) );
INVx5_ASAP7_75t_L g710 ( .A(n_587), .Y(n_710) );
INVx3_ASAP7_75t_L g711 ( .A(n_570), .Y(n_711) );
BUFx3_ASAP7_75t_L g712 ( .A(n_534), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_603), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_563), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_542), .A2(n_431), .B1(n_442), .B2(n_380), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_579), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_593), .Y(n_717) );
OAI33xp33_ASAP7_75t_L g718 ( .A1(n_598), .A2(n_438), .A3(n_437), .B1(n_424), .B2(n_419), .B3(n_417), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_529), .Y(n_719) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_539), .Y(n_720) );
NAND2x1_ASAP7_75t_SL g721 ( .A(n_614), .B(n_409), .Y(n_721) );
INVx3_ASAP7_75t_L g722 ( .A(n_570), .Y(n_722) );
AO22x1_ASAP7_75t_L g723 ( .A1(n_576), .A2(n_404), .B1(n_304), .B2(n_306), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_558), .B(n_414), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_529), .Y(n_725) );
INVxp67_ASAP7_75t_L g726 ( .A(n_530), .Y(n_726) );
NAND2xp33_ASAP7_75t_L g727 ( .A(n_539), .B(n_302), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_572), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_545), .Y(n_729) );
INVx3_ASAP7_75t_L g730 ( .A(n_572), .Y(n_730) );
INVx4_ASAP7_75t_L g731 ( .A(n_587), .Y(n_731) );
INVx2_ASAP7_75t_SL g732 ( .A(n_597), .Y(n_732) );
BUFx2_ASAP7_75t_L g733 ( .A(n_551), .Y(n_733) );
INVx5_ASAP7_75t_L g734 ( .A(n_545), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_597), .B(n_322), .Y(n_735) );
OR2x2_ASAP7_75t_L g736 ( .A(n_597), .B(n_304), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_530), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_595), .A2(n_441), .B1(n_435), .B2(n_360), .C(n_426), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_546), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_546), .Y(n_740) );
INVx3_ASAP7_75t_L g741 ( .A(n_575), .Y(n_741) );
BUFx12f_ASAP7_75t_L g742 ( .A(n_597), .Y(n_742) );
CKINVDCx5p33_ASAP7_75t_R g743 ( .A(n_589), .Y(n_743) );
OR2x6_ASAP7_75t_L g744 ( .A(n_589), .B(n_360), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_569), .B(n_320), .Y(n_745) );
INVxp67_ASAP7_75t_L g746 ( .A(n_534), .Y(n_746) );
O2A1O1Ixp33_ASAP7_75t_L g747 ( .A1(n_547), .A2(n_311), .B(n_312), .C(n_305), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_547), .B(n_306), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_553), .Y(n_749) );
BUFx12f_ASAP7_75t_L g750 ( .A(n_569), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_553), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_586), .B(n_308), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_586), .B(n_308), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_567), .A2(n_374), .B1(n_381), .B2(n_331), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_567), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_594), .B(n_331), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_576), .A2(n_334), .B1(n_342), .B2(n_332), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_588), .Y(n_758) );
INVx2_ASAP7_75t_SL g759 ( .A(n_616), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_594), .A2(n_374), .B1(n_387), .B2(n_381), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_619), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_627), .A2(n_566), .B1(n_539), .B2(n_576), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_634), .A2(n_435), .B1(n_441), .B2(n_360), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_634), .A2(n_441), .B1(n_435), .B2(n_566), .Y(n_764) );
BUFx12f_ASAP7_75t_L g765 ( .A(n_644), .Y(n_765) );
OR2x2_ASAP7_75t_L g766 ( .A(n_639), .B(n_387), .Y(n_766) );
O2A1O1Ixp33_ASAP7_75t_L g767 ( .A1(n_706), .A2(n_329), .B(n_349), .C(n_314), .Y(n_767) );
AND2x4_ASAP7_75t_L g768 ( .A(n_623), .B(n_619), .Y(n_768) );
BUFx2_ASAP7_75t_L g769 ( .A(n_623), .Y(n_769) );
NOR2x1_ASAP7_75t_SL g770 ( .A(n_744), .B(n_566), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_718), .A2(n_441), .B1(n_435), .B2(n_566), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_695), .B(n_616), .Y(n_772) );
INVx2_ASAP7_75t_SL g773 ( .A(n_677), .Y(n_773) );
BUFx3_ASAP7_75t_L g774 ( .A(n_677), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_671), .B(n_395), .Y(n_775) );
INVx5_ASAP7_75t_L g776 ( .A(n_744), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_627), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_718), .A2(n_441), .B1(n_435), .B2(n_566), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_648), .A2(n_590), .B1(n_600), .B2(n_596), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_648), .A2(n_590), .B1(n_600), .B2(n_596), .Y(n_780) );
AOI211xp5_ASAP7_75t_L g781 ( .A1(n_757), .A2(n_383), .B(n_432), .C(n_359), .Y(n_781) );
BUFx2_ASAP7_75t_L g782 ( .A(n_690), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_625), .A2(n_604), .B1(n_612), .B2(n_611), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_712), .Y(n_784) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_658), .Y(n_785) );
INVx6_ASAP7_75t_L g786 ( .A(n_694), .Y(n_786) );
AND2x4_ASAP7_75t_L g787 ( .A(n_732), .B(n_616), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_688), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_749), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_655), .Y(n_790) );
AND2x4_ASAP7_75t_L g791 ( .A(n_670), .B(n_616), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_751), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_631), .A2(n_580), .B1(n_611), .B2(n_604), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_742), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_688), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_726), .A2(n_580), .B1(n_395), .B2(n_425), .Y(n_796) );
NAND2x1p5_ASAP7_75t_L g797 ( .A(n_704), .B(n_616), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_719), .Y(n_798) );
O2A1O1Ixp33_ASAP7_75t_SL g799 ( .A1(n_726), .A2(n_316), .B(n_318), .C(n_315), .Y(n_799) );
CKINVDCx8_ASAP7_75t_R g800 ( .A(n_735), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_624), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_725), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_746), .A2(n_405), .B1(n_427), .B2(n_425), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_625), .Y(n_804) );
INVx1_ASAP7_75t_SL g805 ( .A(n_698), .Y(n_805) );
OAI221xp5_ASAP7_75t_L g806 ( .A1(n_715), .A2(n_620), .B1(n_618), .B2(n_612), .C(n_622), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g807 ( .A1(n_704), .A2(n_427), .B1(n_405), .B2(n_358), .Y(n_807) );
INVx1_ASAP7_75t_SL g808 ( .A(n_629), .Y(n_808) );
INVx3_ASAP7_75t_L g809 ( .A(n_637), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_737), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_651), .A2(n_620), .B1(n_622), .B2(n_618), .Y(n_811) );
INVxp33_ASAP7_75t_SL g812 ( .A(n_703), .Y(n_812) );
BUFx3_ASAP7_75t_L g813 ( .A(n_636), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_651), .A2(n_321), .B1(n_353), .B2(n_319), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_703), .A2(n_365), .B1(n_366), .B2(n_354), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_739), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_740), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_638), .B(n_367), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_674), .B(n_4), .Y(n_819) );
AOI21xp33_ASAP7_75t_L g820 ( .A1(n_743), .A2(n_389), .B(n_371), .Y(n_820) );
AND2x4_ASAP7_75t_L g821 ( .A(n_684), .B(n_368), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_746), .A2(n_378), .B1(n_379), .B2(n_373), .Y(n_822) );
OAI221xp5_ASAP7_75t_L g823 ( .A1(n_715), .A2(n_421), .B1(n_440), .B2(n_430), .C(n_439), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_659), .A2(n_386), .B1(n_390), .B2(n_385), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_641), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_659), .A2(n_396), .B1(n_397), .B2(n_392), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_728), .Y(n_827) );
AO31x2_ASAP7_75t_L g828 ( .A1(n_668), .A2(n_470), .A3(n_468), .B(n_372), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g829 ( .A1(n_651), .A2(n_358), .B1(n_418), .B2(n_328), .Y(n_829) );
AND2x4_ASAP7_75t_L g830 ( .A(n_658), .B(n_398), .Y(n_830) );
AND2x4_ASAP7_75t_L g831 ( .A(n_646), .B(n_401), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_630), .A2(n_672), .B1(n_643), .B2(n_664), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_632), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g834 ( .A1(n_661), .A2(n_488), .B(n_484), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g835 ( .A1(n_757), .A2(n_418), .B1(n_328), .B2(n_410), .Y(n_835) );
INVx2_ASAP7_75t_SL g836 ( .A(n_681), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_630), .A2(n_416), .B1(n_420), .B2(n_403), .Y(n_837) );
BUFx2_ASAP7_75t_L g838 ( .A(n_690), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_672), .A2(n_434), .B1(n_436), .B2(n_428), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_647), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_633), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_657), .Y(n_842) );
OR2x2_ASAP7_75t_L g843 ( .A(n_736), .B(n_5), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_699), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_697), .A2(n_349), .B1(n_433), .B2(n_372), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_682), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_642), .A2(n_700), .B1(n_716), .B2(n_714), .Y(n_847) );
INVx2_ASAP7_75t_SL g848 ( .A(n_694), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_709), .B(n_679), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_679), .B(n_6), .Y(n_850) );
AND2x6_ASAP7_75t_L g851 ( .A(n_628), .B(n_433), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_653), .B(n_7), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_642), .A2(n_384), .B1(n_333), .B2(n_466), .Y(n_853) );
NAND2xp5_ASAP7_75t_SL g854 ( .A(n_691), .B(n_384), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_686), .B(n_7), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_640), .Y(n_856) );
AO31x2_ASAP7_75t_L g857 ( .A1(n_668), .A2(n_468), .A3(n_470), .B(n_484), .Y(n_857) );
INVx3_ASAP7_75t_L g858 ( .A(n_637), .Y(n_858) );
BUFx2_ASAP7_75t_SL g859 ( .A(n_646), .Y(n_859) );
NOR3xp33_ASAP7_75t_L g860 ( .A(n_723), .B(n_476), .C(n_470), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_713), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_686), .B(n_9), .Y(n_862) );
INVx2_ASAP7_75t_SL g863 ( .A(n_721), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_680), .B(n_9), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_700), .A2(n_476), .B1(n_468), .B2(n_470), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_717), .B(n_10), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_691), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_735), .B(n_10), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_680), .B(n_11), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_724), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_754), .B(n_724), .Y(n_871) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_650), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_645), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_652), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_650), .Y(n_875) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_661), .A2(n_468), .B(n_484), .Y(n_876) );
INVx3_ASAP7_75t_L g877 ( .A(n_750), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_705), .B(n_11), .Y(n_878) );
OAI22xp33_ASAP7_75t_L g879 ( .A1(n_744), .A2(n_384), .B1(n_476), .B2(n_16), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_696), .A2(n_476), .B1(n_384), .B2(n_475), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_707), .A2(n_384), .B1(n_476), .B2(n_16), .Y(n_881) );
OR2x2_ASAP7_75t_L g882 ( .A(n_705), .B(n_13), .Y(n_882) );
OAI221xp5_ASAP7_75t_L g883 ( .A1(n_696), .A2(n_475), .B1(n_484), .B2(n_488), .C(n_508), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_755), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_649), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_738), .A2(n_475), .B1(n_488), .B2(n_508), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_748), .B(n_13), .Y(n_887) );
AO31x2_ASAP7_75t_L g888 ( .A1(n_758), .A2(n_508), .A3(n_485), .B(n_515), .Y(n_888) );
OAI221xp5_ASAP7_75t_L g889 ( .A1(n_738), .A2(n_508), .B1(n_485), .B2(n_515), .C(n_516), .Y(n_889) );
BUFx12f_ASAP7_75t_L g890 ( .A(n_649), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_748), .Y(n_891) );
BUFx2_ASAP7_75t_L g892 ( .A(n_675), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_693), .Y(n_893) );
INVx4_ASAP7_75t_SL g894 ( .A(n_628), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_733), .A2(n_485), .B1(n_515), .B2(n_516), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_673), .A2(n_516), .B1(n_517), .B2(n_519), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_761), .Y(n_897) );
CKINVDCx6p67_ASAP7_75t_R g898 ( .A(n_675), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_660), .A2(n_519), .B1(n_517), .B2(n_510), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_654), .A2(n_15), .B1(n_17), .B2(n_18), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_760), .B(n_15), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_654), .A2(n_17), .B1(n_18), .B2(n_20), .Y(n_902) );
INVx6_ASAP7_75t_L g903 ( .A(n_701), .Y(n_903) );
OAI22xp33_ASAP7_75t_L g904 ( .A1(n_662), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_904) );
AO221x2_ASAP7_75t_L g905 ( .A1(n_747), .A2(n_23), .B1(n_24), .B2(n_26), .C(n_27), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_673), .B(n_24), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_626), .Y(n_907) );
CKINVDCx6p67_ASAP7_75t_R g908 ( .A(n_701), .Y(n_908) );
BUFx2_ASAP7_75t_SL g909 ( .A(n_759), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_626), .Y(n_910) );
OA21x2_ASAP7_75t_L g911 ( .A1(n_876), .A2(n_663), .B(n_635), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_805), .B(n_747), .Y(n_912) );
OAI221xp5_ASAP7_75t_L g913 ( .A1(n_832), .A2(n_678), .B1(n_702), .B2(n_745), .C(n_756), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_769), .Y(n_914) );
AOI221xp5_ASAP7_75t_L g915 ( .A1(n_812), .A2(n_702), .B1(n_676), .B2(n_669), .C(n_685), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_847), .A2(n_756), .B1(n_753), .B2(n_676), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_832), .A2(n_722), .B1(n_730), .B2(n_711), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_777), .A2(n_752), .B1(n_753), .B2(n_669), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_864), .A2(n_711), .B1(n_730), .B2(n_722), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_869), .A2(n_741), .B1(n_685), .B2(n_667), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_849), .B(n_741), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_798), .Y(n_922) );
AND2x4_ASAP7_75t_L g923 ( .A(n_782), .B(n_734), .Y(n_923) );
AOI21xp33_ASAP7_75t_L g924 ( .A1(n_767), .A2(n_727), .B(n_710), .Y(n_924) );
INVx3_ASAP7_75t_L g925 ( .A(n_908), .Y(n_925) );
AOI321xp33_ASAP7_75t_L g926 ( .A1(n_781), .A2(n_689), .A3(n_692), .B1(n_635), .B2(n_30), .C(n_31), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_905), .A2(n_731), .B1(n_729), .B2(n_701), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_814), .A2(n_656), .B1(n_665), .B2(n_687), .Y(n_928) );
AOI22xp33_ASAP7_75t_SL g929 ( .A1(n_905), .A2(n_656), .B1(n_683), .B2(n_687), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_814), .A2(n_870), .B1(n_872), .B2(n_837), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_871), .A2(n_731), .B1(n_729), .B2(n_701), .Y(n_931) );
INVx3_ASAP7_75t_L g932 ( .A(n_797), .Y(n_932) );
BUFx2_ASAP7_75t_R g933 ( .A(n_794), .Y(n_933) );
INVx1_ASAP7_75t_SL g934 ( .A(n_885), .Y(n_934) );
NAND2xp5_ASAP7_75t_SL g935 ( .A(n_776), .B(n_656), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_891), .A2(n_710), .B1(n_734), .B2(n_720), .Y(n_936) );
A2O1A1Ixp33_ASAP7_75t_L g937 ( .A1(n_767), .A2(n_710), .B(n_734), .C(n_720), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_862), .A2(n_710), .B1(n_734), .B2(n_720), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_800), .B(n_708), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_835), .A2(n_708), .B1(n_687), .B2(n_683), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_815), .A2(n_708), .B1(n_683), .B2(n_666), .C(n_665), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_835), .A2(n_666), .B1(n_665), .B2(n_519), .Y(n_942) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_775), .B(n_666), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_801), .B(n_27), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_808), .B(n_28), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_872), .A2(n_28), .B1(n_29), .B2(n_32), .Y(n_946) );
AND2x4_ASAP7_75t_L g947 ( .A(n_838), .B(n_32), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_861), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_897), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_901), .A2(n_519), .B1(n_517), .B2(n_510), .Y(n_950) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_790), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_893), .A2(n_519), .B1(n_517), .B2(n_510), .Y(n_952) );
NOR2xp33_ASAP7_75t_L g953 ( .A(n_804), .B(n_35), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_819), .A2(n_519), .B1(n_517), .B2(n_510), .Y(n_954) );
INVx2_ASAP7_75t_L g955 ( .A(n_802), .Y(n_955) );
BUFx12f_ASAP7_75t_L g956 ( .A(n_765), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_855), .A2(n_519), .B1(n_517), .B2(n_510), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_816), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_821), .A2(n_519), .B1(n_517), .B2(n_510), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_821), .A2(n_517), .B1(n_510), .B2(n_505), .Y(n_960) );
AOI221xp5_ASAP7_75t_L g961 ( .A1(n_823), .A2(n_510), .B1(n_505), .B2(n_503), .C(n_495), .Y(n_961) );
BUFx4f_ASAP7_75t_SL g962 ( .A(n_890), .Y(n_962) );
OA21x2_ASAP7_75t_L g963 ( .A1(n_834), .A2(n_495), .B(n_490), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_867), .B(n_37), .Y(n_964) );
AOI21xp5_ASAP7_75t_L g965 ( .A1(n_834), .A2(n_495), .B(n_490), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_810), .Y(n_966) );
INVx5_ASAP7_75t_SL g967 ( .A(n_898), .Y(n_967) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_837), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_968) );
AOI22xp33_ASAP7_75t_SL g969 ( .A1(n_776), .A2(n_38), .B1(n_41), .B2(n_42), .Y(n_969) );
OAI221xp5_ASAP7_75t_L g970 ( .A1(n_845), .A2(n_505), .B1(n_503), .B2(n_495), .C(n_490), .Y(n_970) );
BUFx2_ASAP7_75t_L g971 ( .A(n_772), .Y(n_971) );
OAI21xp5_ASAP7_75t_SL g972 ( .A1(n_829), .A2(n_41), .B(n_42), .Y(n_972) );
OR2x6_ASAP7_75t_L g973 ( .A(n_859), .B(n_43), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_824), .A2(n_505), .B1(n_503), .B2(n_495), .C(n_490), .Y(n_974) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_776), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_975) );
OAI211xp5_ASAP7_75t_L g976 ( .A1(n_829), .A2(n_505), .B(n_503), .C(n_495), .Y(n_976) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_875), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_852), .A2(n_904), .B1(n_795), .B2(n_788), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_853), .A2(n_44), .B1(n_46), .B2(n_47), .Y(n_979) );
BUFx8_ASAP7_75t_L g980 ( .A(n_836), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_817), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_766), .B(n_47), .Y(n_982) );
BUFx6f_ASAP7_75t_L g983 ( .A(n_776), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_853), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_984) );
AOI221xp5_ASAP7_75t_L g985 ( .A1(n_826), .A2(n_505), .B1(n_503), .B2(n_490), .C(n_52), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_811), .A2(n_48), .B1(n_49), .B2(n_51), .Y(n_986) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_807), .A2(n_796), .B1(n_803), .B2(n_850), .Y(n_987) );
BUFx6f_ASAP7_75t_L g988 ( .A(n_772), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_811), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_989) );
OAI21xp5_ASAP7_75t_L g990 ( .A1(n_878), .A2(n_53), .B(n_54), .Y(n_990) );
OAI21x1_ASAP7_75t_L g991 ( .A1(n_762), .A2(n_854), .B(n_896), .Y(n_991) );
OR2x2_ASAP7_75t_L g992 ( .A(n_843), .B(n_55), .Y(n_992) );
INVx3_ASAP7_75t_L g993 ( .A(n_797), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_904), .A2(n_503), .B1(n_490), .B2(n_59), .Y(n_994) );
NOR2x1_ASAP7_75t_L g995 ( .A(n_892), .B(n_56), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_882), .A2(n_490), .B1(n_59), .B2(n_62), .Y(n_996) );
INVx2_ASAP7_75t_L g997 ( .A(n_789), .Y(n_997) );
AO21x2_ASAP7_75t_L g998 ( .A1(n_860), .A2(n_97), .B(n_94), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_839), .A2(n_58), .B1(n_62), .B2(n_63), .Y(n_999) );
OAI211xp5_ASAP7_75t_L g1000 ( .A1(n_820), .A2(n_58), .B(n_63), .C(n_64), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_830), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_1001) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_875), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1003 ( .A1(n_879), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_887), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_1004) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_770), .A2(n_69), .B1(n_70), .B2(n_71), .Y(n_1005) );
OAI221xp5_ASAP7_75t_L g1006 ( .A1(n_839), .A2(n_70), .B1(n_72), .B2(n_73), .C(n_74), .Y(n_1006) );
OAI321xp33_ASAP7_75t_L g1007 ( .A1(n_879), .A2(n_73), .A3(n_74), .B1(n_75), .B2(n_76), .C(n_77), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_792), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_825), .B(n_75), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_840), .Y(n_1010) );
OAI221xp5_ASAP7_75t_L g1011 ( .A1(n_881), .A2(n_78), .B1(n_79), .B2(n_80), .C(n_81), .Y(n_1011) );
AOI22xp5_ASAP7_75t_L g1012 ( .A1(n_807), .A2(n_78), .B1(n_79), .B2(n_81), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_842), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_846), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_860), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_793), .A2(n_83), .B1(n_84), .B2(n_86), .Y(n_1016) );
OAI21xp5_ASAP7_75t_L g1017 ( .A1(n_886), .A2(n_87), .B(n_98), .Y(n_1017) );
AOI21x1_ASAP7_75t_L g1018 ( .A1(n_768), .A2(n_196), .B(n_99), .Y(n_1018) );
INVx3_ASAP7_75t_L g1019 ( .A(n_809), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_900), .A2(n_87), .B1(n_104), .B2(n_106), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_881), .A2(n_107), .B1(n_108), .B2(n_110), .Y(n_1021) );
INVx2_ASAP7_75t_L g1022 ( .A(n_884), .Y(n_1022) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_822), .A2(n_114), .B1(n_115), .B2(n_116), .C(n_117), .Y(n_1023) );
OR2x6_ASAP7_75t_L g1024 ( .A(n_909), .B(n_118), .Y(n_1024) );
NAND3xp33_ASAP7_75t_L g1025 ( .A(n_763), .B(n_119), .C(n_122), .Y(n_1025) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_902), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_785), .A2(n_126), .B1(n_127), .B2(n_128), .Y(n_1027) );
A2O1A1Ixp33_ASAP7_75t_L g1028 ( .A1(n_866), .A2(n_906), .B(n_768), .C(n_763), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_785), .B(n_131), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_818), .A2(n_132), .B1(n_135), .B2(n_140), .C(n_141), .Y(n_1030) );
AOI221xp5_ASAP7_75t_L g1031 ( .A1(n_799), .A2(n_142), .B1(n_145), .B2(n_147), .C(n_148), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_784), .B(n_150), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_784), .A2(n_151), .B1(n_153), .B2(n_160), .Y(n_1033) );
OAI21xp33_ASAP7_75t_L g1034 ( .A1(n_771), .A2(n_161), .B(n_162), .Y(n_1034) );
OAI21x1_ASAP7_75t_L g1035 ( .A1(n_896), .A2(n_163), .B(n_164), .Y(n_1035) );
OAI211xp5_ASAP7_75t_L g1036 ( .A1(n_868), .A2(n_165), .B(n_169), .C(n_171), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_809), .B(n_173), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_831), .A2(n_174), .B1(n_175), .B2(n_177), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_833), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_827), .Y(n_1040) );
OA21x2_ASAP7_75t_L g1041 ( .A1(n_771), .A2(n_178), .B(n_181), .Y(n_1041) );
OAI211xp5_ASAP7_75t_L g1042 ( .A1(n_951), .A2(n_844), .B(n_863), .C(n_877), .Y(n_1042) );
INVx2_ASAP7_75t_L g1043 ( .A(n_963), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1044 ( .A1(n_926), .A2(n_773), .B1(n_848), .B2(n_877), .C(n_764), .Y(n_1044) );
BUFx6f_ASAP7_75t_L g1045 ( .A(n_983), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_963), .Y(n_1046) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_962), .Y(n_1047) );
BUFx2_ASAP7_75t_L g1048 ( .A(n_1024), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_948), .B(n_813), .Y(n_1049) );
OA332x1_ASAP7_75t_L g1050 ( .A1(n_999), .A2(n_865), .A3(n_880), .B1(n_831), .B2(n_828), .B3(n_857), .C1(n_778), .C2(n_786), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_978), .A2(n_778), .B1(n_780), .B2(n_779), .Y(n_1051) );
AND2x4_ASAP7_75t_L g1052 ( .A(n_932), .B(n_858), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_978), .A2(n_780), .B1(n_779), .B2(n_783), .Y(n_1053) );
AOI21xp5_ASAP7_75t_SL g1054 ( .A1(n_1024), .A2(n_851), .B(n_787), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1002), .B(n_858), .Y(n_1055) );
OAI221xp5_ASAP7_75t_L g1056 ( .A1(n_972), .A2(n_764), .B1(n_774), .B2(n_783), .C(n_886), .Y(n_1056) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_1003), .A2(n_806), .B1(n_907), .B2(n_910), .C(n_787), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_973), .A2(n_786), .B1(n_851), .B2(n_874), .Y(n_1058) );
OAI221xp5_ASAP7_75t_SL g1059 ( .A1(n_973), .A2(n_895), .B1(n_856), .B2(n_873), .C(n_841), .Y(n_1059) );
INVx2_ASAP7_75t_SL g1060 ( .A(n_962), .Y(n_1060) );
AND2x4_ASAP7_75t_L g1061 ( .A(n_932), .B(n_894), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_992), .B(n_828), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_1003), .A2(n_791), .B1(n_883), .B2(n_889), .C(n_895), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_947), .B(n_786), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_947), .B(n_791), .Y(n_1065) );
OR2x2_ASAP7_75t_L g1066 ( .A(n_922), .B(n_828), .Y(n_1066) );
OAI31xp33_ASAP7_75t_L g1067 ( .A1(n_975), .A2(n_899), .A3(n_851), .B(n_828), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_973), .A2(n_912), .B1(n_994), .B2(n_930), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_994), .A2(n_851), .B1(n_903), .B2(n_894), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_987), .A2(n_903), .B1(n_894), .B2(n_857), .Y(n_1070) );
OAI221xp5_ASAP7_75t_L g1071 ( .A1(n_951), .A2(n_903), .B1(n_857), .B2(n_888), .C(n_189), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_958), .B(n_857), .Y(n_1072) );
OA21x2_ASAP7_75t_L g1073 ( .A1(n_965), .A2(n_888), .B(n_185), .Y(n_1073) );
OAI321xp33_ASAP7_75t_L g1074 ( .A1(n_975), .A2(n_1011), .A3(n_927), .B1(n_1006), .B2(n_1012), .C(n_1021), .Y(n_1074) );
AND2x4_ASAP7_75t_L g1075 ( .A(n_993), .B(n_888), .Y(n_1075) );
NAND4xp25_ASAP7_75t_L g1076 ( .A(n_1001), .B(n_184), .C(n_187), .D(n_190), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g1077 ( .A(n_967), .Y(n_1077) );
AOI21xp5_ASAP7_75t_L g1078 ( .A1(n_976), .A2(n_888), .B(n_197), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_981), .Y(n_1079) );
AOI33xp33_ASAP7_75t_L g1080 ( .A1(n_1001), .A2(n_295), .A3(n_199), .B1(n_200), .B2(n_202), .B3(n_203), .Y(n_1080) );
BUFx3_ASAP7_75t_L g1081 ( .A(n_923), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_920), .A2(n_194), .B1(n_204), .B2(n_206), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_977), .B(n_207), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1010), .Y(n_1084) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_980), .Y(n_1085) );
OAI21xp5_ASAP7_75t_SL g1086 ( .A1(n_929), .A2(n_212), .B(n_213), .Y(n_1086) );
AND2x4_ASAP7_75t_L g1087 ( .A(n_993), .B(n_215), .Y(n_1087) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_1037), .B(n_220), .Y(n_1088) );
OAI221xp5_ASAP7_75t_SL g1089 ( .A1(n_927), .A2(n_222), .B1(n_224), .B2(n_229), .C(n_231), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_955), .B(n_232), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1014), .Y(n_1091) );
NOR2xp33_ASAP7_75t_L g1092 ( .A(n_921), .B(n_233), .Y(n_1092) );
OA21x2_ASAP7_75t_L g1093 ( .A1(n_991), .A2(n_234), .B(n_236), .Y(n_1093) );
INVxp67_ASAP7_75t_SL g1094 ( .A(n_928), .Y(n_1094) );
OAI222xp33_ASAP7_75t_L g1095 ( .A1(n_929), .A2(n_238), .B1(n_240), .B2(n_243), .C1(n_244), .C2(n_245), .Y(n_1095) );
AOI22xp33_ASAP7_75t_SL g1096 ( .A1(n_977), .A2(n_249), .B1(n_252), .B2(n_253), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_949), .Y(n_1097) );
AO21x2_ASAP7_75t_L g1098 ( .A1(n_1028), .A2(n_254), .B(n_257), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_982), .B(n_258), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_919), .A2(n_263), .B1(n_264), .B2(n_267), .Y(n_1100) );
AO21x2_ASAP7_75t_L g1101 ( .A1(n_1017), .A2(n_268), .B(n_269), .Y(n_1101) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_1007), .A2(n_271), .B1(n_274), .B2(n_277), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_919), .A2(n_278), .B1(n_279), .B2(n_282), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_920), .A2(n_283), .B1(n_286), .B2(n_287), .Y(n_1104) );
OA21x2_ASAP7_75t_L g1105 ( .A1(n_952), .A2(n_289), .B(n_291), .Y(n_1105) );
OAI211xp5_ASAP7_75t_L g1106 ( .A1(n_969), .A2(n_292), .B(n_294), .C(n_995), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_983), .Y(n_1107) );
OAI221xp5_ASAP7_75t_L g1108 ( .A1(n_1020), .A2(n_996), .B1(n_990), .B2(n_1005), .C(n_1015), .Y(n_1108) );
INVx2_ASAP7_75t_SL g1109 ( .A(n_980), .Y(n_1109) );
OR2x2_ASAP7_75t_L g1110 ( .A(n_966), .B(n_1013), .Y(n_1110) );
OAI21xp33_ASAP7_75t_L g1111 ( .A1(n_1004), .A2(n_969), .B(n_1015), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1112 ( .A1(n_968), .A2(n_946), .B1(n_986), .B2(n_989), .C(n_1016), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_917), .A2(n_913), .B1(n_914), .B2(n_953), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_917), .A2(n_964), .B1(n_996), .B2(n_915), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1022), .Y(n_1115) );
AOI22xp5_ASAP7_75t_L g1116 ( .A1(n_943), .A2(n_1000), .B1(n_918), .B2(n_945), .Y(n_1116) );
INVx2_ASAP7_75t_L g1117 ( .A(n_997), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1008), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1039), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1040), .Y(n_1120) );
AOI222xp33_ASAP7_75t_L g1121 ( .A1(n_967), .A2(n_979), .B1(n_984), .B2(n_934), .C1(n_944), .C2(n_1004), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_983), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_931), .A2(n_940), .B1(n_942), .B2(n_1021), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_971), .B(n_967), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_925), .B(n_923), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_1020), .A2(n_985), .B1(n_916), .B2(n_1009), .Y(n_1126) );
OA21x2_ASAP7_75t_L g1127 ( .A1(n_952), .A2(n_1035), .B(n_937), .Y(n_1127) );
BUFx3_ASAP7_75t_L g1128 ( .A(n_925), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_988), .B(n_1019), .Y(n_1129) );
OAI211xp5_ASAP7_75t_L g1130 ( .A1(n_1026), .A2(n_1038), .B(n_1023), .C(n_939), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_988), .B(n_1037), .Y(n_1131) );
OAI221xp5_ASAP7_75t_L g1132 ( .A1(n_1026), .A2(n_931), .B1(n_950), .B2(n_954), .C(n_938), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1032), .Y(n_1133) );
HB1xp67_ASAP7_75t_L g1134 ( .A(n_983), .Y(n_1134) );
NAND4xp25_ASAP7_75t_SL g1135 ( .A(n_1031), .B(n_1030), .C(n_933), .D(n_1027), .Y(n_1135) );
OAI222xp33_ASAP7_75t_L g1136 ( .A1(n_941), .A2(n_1033), .B1(n_1029), .B2(n_935), .C1(n_1018), .C2(n_970), .Y(n_1136) );
OAI321xp33_ASAP7_75t_L g1137 ( .A1(n_1036), .A2(n_1025), .A3(n_1034), .B1(n_957), .B2(n_936), .C(n_959), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_961), .A2(n_1041), .B1(n_960), .B2(n_974), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_998), .Y(n_1139) );
NOR2x1_ASAP7_75t_SL g1140 ( .A(n_998), .B(n_956), .Y(n_1140) );
OAI33xp33_ASAP7_75t_L g1141 ( .A1(n_924), .A2(n_904), .A3(n_1003), .B1(n_975), .B2(n_946), .B3(n_999), .Y(n_1141) );
INVx1_ASAP7_75t_SL g1142 ( .A(n_1077), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1097), .B(n_911), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1079), .Y(n_1144) );
AOI211x1_ASAP7_75t_SL g1145 ( .A1(n_1076), .A2(n_911), .B(n_1049), .C(n_1097), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_1068), .A2(n_1058), .B1(n_1108), .B2(n_1048), .Y(n_1146) );
OAI21xp5_ASAP7_75t_SL g1147 ( .A1(n_1058), .A2(n_1086), .B(n_1109), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_1068), .A2(n_1088), .B1(n_1069), .B2(n_1054), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1117), .B(n_1072), .Y(n_1149) );
OAI33xp33_ASAP7_75t_L g1150 ( .A1(n_1084), .A2(n_1091), .A3(n_1062), .B1(n_1102), .B2(n_1115), .B3(n_1119), .Y(n_1150) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1043), .Y(n_1151) );
INVx2_ASAP7_75t_SL g1152 ( .A(n_1107), .Y(n_1152) );
INVx2_ASAP7_75t_L g1153 ( .A(n_1046), .Y(n_1153) );
AO21x2_ASAP7_75t_L g1154 ( .A1(n_1139), .A2(n_1046), .B(n_1070), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1066), .Y(n_1155) );
OAI33xp33_ASAP7_75t_L g1156 ( .A1(n_1102), .A2(n_1111), .A3(n_1053), .B1(n_1110), .B2(n_1118), .B3(n_1051), .Y(n_1156) );
OAI22xp33_ASAP7_75t_L g1157 ( .A1(n_1056), .A2(n_1044), .B1(n_1085), .B2(n_1071), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1120), .Y(n_1158) );
OAI21xp33_ASAP7_75t_L g1159 ( .A1(n_1080), .A2(n_1121), .B(n_1126), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1075), .B(n_1107), .Y(n_1160) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1075), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1055), .B(n_1113), .Y(n_1162) );
NAND2xp5_ASAP7_75t_SL g1163 ( .A(n_1067), .B(n_1096), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1122), .B(n_1134), .Y(n_1164) );
OAI31xp33_ASAP7_75t_L g1165 ( .A1(n_1059), .A2(n_1130), .A3(n_1106), .B(n_1088), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1125), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1090), .Y(n_1167) );
INVx4_ASAP7_75t_L g1168 ( .A(n_1081), .Y(n_1168) );
AND2x2_ASAP7_75t_SL g1169 ( .A(n_1069), .B(n_1105), .Y(n_1169) );
INVx2_ASAP7_75t_SL g1170 ( .A(n_1045), .Y(n_1170) );
NOR3xp33_ASAP7_75t_SL g1171 ( .A(n_1135), .B(n_1141), .C(n_1095), .Y(n_1171) );
NAND2xp5_ASAP7_75t_SL g1172 ( .A(n_1096), .B(n_1080), .Y(n_1172) );
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_1141), .A2(n_1116), .B1(n_1114), .B2(n_1112), .Y(n_1173) );
INVx3_ASAP7_75t_L g1174 ( .A(n_1045), .Y(n_1174) );
OAI33xp33_ASAP7_75t_L g1175 ( .A1(n_1133), .A2(n_1123), .A3(n_1100), .B1(n_1103), .B2(n_1138), .B3(n_1129), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1065), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1073), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1113), .B(n_1064), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1114), .B(n_1131), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1094), .B(n_1045), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1045), .B(n_1083), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1094), .B(n_1126), .Y(n_1182) );
AO21x2_ASAP7_75t_L g1183 ( .A1(n_1078), .A2(n_1074), .B(n_1098), .Y(n_1183) );
OAI221xp5_ASAP7_75t_L g1184 ( .A1(n_1132), .A2(n_1089), .B1(n_1057), .B2(n_1128), .C(n_1082), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1140), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1087), .Y(n_1186) );
NOR2xp33_ASAP7_75t_L g1187 ( .A(n_1047), .B(n_1060), .Y(n_1187) );
NAND2x1_ASAP7_75t_L g1188 ( .A(n_1105), .B(n_1093), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1073), .Y(n_1189) );
AND2x4_ASAP7_75t_L g1190 ( .A(n_1061), .B(n_1087), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1124), .Y(n_1191) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1093), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1099), .B(n_1127), .Y(n_1193) );
NAND3xp33_ASAP7_75t_L g1194 ( .A(n_1092), .B(n_1104), .C(n_1063), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1127), .B(n_1052), .Y(n_1195) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1093), .Y(n_1196) );
AND2x4_ASAP7_75t_L g1197 ( .A(n_1101), .B(n_1050), .Y(n_1197) );
AND2x4_ASAP7_75t_SL g1198 ( .A(n_1136), .B(n_1105), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1199 ( .A(n_1127), .B(n_1137), .Y(n_1199) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_1068), .A2(n_978), .B1(n_1058), .B2(n_994), .Y(n_1200) );
NAND2xp5_ASAP7_75t_SL g1201 ( .A(n_1048), .B(n_929), .Y(n_1201) );
NAND4xp25_ASAP7_75t_SL g1202 ( .A(n_1042), .B(n_1077), .C(n_951), .D(n_1054), .Y(n_1202) );
AOI221xp5_ASAP7_75t_L g1203 ( .A1(n_1141), .A2(n_904), .B1(n_812), .B2(n_536), .C(n_869), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1097), .B(n_1117), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1097), .B(n_1117), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1079), .Y(n_1206) );
INVx2_ASAP7_75t_L g1207 ( .A(n_1043), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1072), .Y(n_1208) );
OAI221xp5_ASAP7_75t_L g1209 ( .A1(n_1042), .A2(n_972), .B1(n_951), .B2(n_1044), .C(n_978), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1204), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1204), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1205), .Y(n_1212) );
INVx4_ASAP7_75t_L g1213 ( .A(n_1190), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1149), .B(n_1161), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1149), .B(n_1161), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1208), .B(n_1155), .Y(n_1216) );
NOR2xp33_ASAP7_75t_L g1217 ( .A(n_1142), .B(n_1187), .Y(n_1217) );
OAI21xp5_ASAP7_75t_L g1218 ( .A1(n_1171), .A2(n_1159), .B(n_1172), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1195), .B(n_1208), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1195), .B(n_1143), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1205), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1173), .B(n_1158), .Y(n_1222) );
INVx2_ASAP7_75t_SL g1223 ( .A(n_1152), .Y(n_1223) );
AOI211xp5_ASAP7_75t_SL g1224 ( .A1(n_1157), .A2(n_1209), .B(n_1148), .C(n_1147), .Y(n_1224) );
NOR2xp33_ASAP7_75t_R g1225 ( .A(n_1202), .B(n_1190), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1155), .B(n_1182), .Y(n_1226) );
NOR3xp33_ASAP7_75t_SL g1227 ( .A(n_1146), .B(n_1184), .C(n_1163), .Y(n_1227) );
OR2x6_ASAP7_75t_L g1228 ( .A(n_1201), .B(n_1188), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1151), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1182), .B(n_1160), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1207), .Y(n_1231) );
NOR3xp33_ASAP7_75t_SL g1232 ( .A(n_1163), .B(n_1203), .C(n_1165), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1193), .B(n_1153), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1193), .B(n_1207), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1179), .B(n_1180), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1144), .B(n_1206), .Y(n_1236) );
NOR3xp33_ASAP7_75t_SL g1237 ( .A(n_1175), .B(n_1172), .C(n_1156), .Y(n_1237) );
NOR3xp33_ASAP7_75t_SL g1238 ( .A(n_1200), .B(n_1194), .C(n_1178), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1166), .B(n_1162), .Y(n_1239) );
NOR2xp33_ASAP7_75t_L g1240 ( .A(n_1191), .B(n_1176), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1164), .B(n_1197), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1197), .B(n_1179), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1197), .B(n_1154), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1154), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1154), .B(n_1169), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1169), .B(n_1180), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1167), .B(n_1186), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1181), .B(n_1177), .Y(n_1248) );
NOR3xp33_ASAP7_75t_L g1249 ( .A(n_1185), .B(n_1201), .C(n_1150), .Y(n_1249) );
AND2x4_ASAP7_75t_L g1250 ( .A(n_1174), .B(n_1198), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1199), .B(n_1168), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1189), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1236), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1216), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1239), .B(n_1145), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1216), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1222), .B(n_1170), .Y(n_1257) );
NOR2xp33_ASAP7_75t_L g1258 ( .A(n_1218), .B(n_1183), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1247), .Y(n_1259) );
NAND4xp25_ASAP7_75t_L g1260 ( .A(n_1224), .B(n_1189), .C(n_1174), .D(n_1192), .Y(n_1260) );
NAND2xp33_ASAP7_75t_R g1261 ( .A(n_1225), .B(n_1196), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1210), .B(n_1196), .Y(n_1262) );
OR2x2_ASAP7_75t_L g1263 ( .A(n_1230), .B(n_1235), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1211), .B(n_1212), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1214), .B(n_1215), .Y(n_1265) );
OR2x6_ASAP7_75t_L g1266 ( .A(n_1213), .B(n_1228), .Y(n_1266) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1226), .B(n_1240), .Y(n_1267) );
AND2x4_ASAP7_75t_L g1268 ( .A(n_1241), .B(n_1242), .Y(n_1268) );
AOI21xp5_ASAP7_75t_L g1269 ( .A1(n_1223), .A2(n_1224), .B(n_1228), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1220), .B(n_1219), .Y(n_1270) );
INVx2_ASAP7_75t_SL g1271 ( .A(n_1223), .Y(n_1271) );
NAND3x1_ASAP7_75t_L g1272 ( .A(n_1249), .B(n_1243), .C(n_1245), .Y(n_1272) );
OAI221xp5_ASAP7_75t_L g1273 ( .A1(n_1227), .A2(n_1232), .B1(n_1238), .B2(n_1237), .C(n_1217), .Y(n_1273) );
XNOR2x1_ASAP7_75t_L g1274 ( .A(n_1273), .B(n_1235), .Y(n_1274) );
XNOR2xp5_ASAP7_75t_L g1275 ( .A(n_1272), .B(n_1219), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1276 ( .A(n_1267), .B(n_1213), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1264), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1278 ( .A(n_1253), .B(n_1221), .Y(n_1278) );
AOI22xp5_ASAP7_75t_L g1279 ( .A1(n_1261), .A2(n_1246), .B1(n_1245), .B2(n_1248), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1254), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1270), .B(n_1220), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1256), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1283 ( .A(n_1259), .B(n_1251), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1265), .B(n_1243), .Y(n_1284) );
NAND2xp33_ASAP7_75t_L g1285 ( .A(n_1272), .B(n_1251), .Y(n_1285) );
OR2x2_ASAP7_75t_L g1286 ( .A(n_1263), .B(n_1234), .Y(n_1286) );
O2A1O1Ixp33_ASAP7_75t_L g1287 ( .A1(n_1258), .A2(n_1228), .B(n_1244), .C(n_1246), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1257), .Y(n_1288) );
OAI22xp5_ASAP7_75t_L g1289 ( .A1(n_1269), .A2(n_1250), .B1(n_1233), .B2(n_1229), .Y(n_1289) );
XNOR2x2_ASAP7_75t_L g1290 ( .A(n_1260), .B(n_1231), .Y(n_1290) );
INVx3_ASAP7_75t_L g1291 ( .A(n_1266), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1268), .B(n_1252), .Y(n_1292) );
BUFx2_ASAP7_75t_L g1293 ( .A(n_1271), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1262), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1255), .Y(n_1295) );
NOR2xp33_ASAP7_75t_L g1296 ( .A(n_1274), .B(n_1295), .Y(n_1296) );
AOI21xp33_ASAP7_75t_L g1297 ( .A1(n_1274), .A2(n_1285), .B(n_1287), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1288), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1283), .B(n_1294), .Y(n_1299) );
NAND2xp33_ASAP7_75t_SL g1300 ( .A(n_1275), .B(n_1261), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1286), .Y(n_1301) );
AND2x4_ASAP7_75t_L g1302 ( .A(n_1291), .B(n_1293), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1302), .B(n_1284), .Y(n_1303) );
AOI22xp5_ASAP7_75t_L g1304 ( .A1(n_1296), .A2(n_1276), .B1(n_1289), .B2(n_1291), .Y(n_1304) );
NAND4xp25_ASAP7_75t_SL g1305 ( .A(n_1297), .B(n_1279), .C(n_1290), .D(n_1292), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1302), .B(n_1284), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1298), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1307), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1304), .Y(n_1309) );
NOR3xp33_ASAP7_75t_L g1310 ( .A(n_1305), .B(n_1300), .C(n_1299), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1308), .Y(n_1311) );
AO22x2_ASAP7_75t_L g1312 ( .A1(n_1309), .A2(n_1306), .B1(n_1303), .B2(n_1301), .Y(n_1312) );
NAND3x1_ASAP7_75t_L g1313 ( .A(n_1310), .B(n_1281), .C(n_1278), .Y(n_1313) );
AND2x2_ASAP7_75t_SL g1314 ( .A(n_1311), .B(n_1308), .Y(n_1314) );
INVx2_ASAP7_75t_L g1315 ( .A(n_1312), .Y(n_1315) );
BUFx2_ASAP7_75t_L g1316 ( .A(n_1315), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1314), .Y(n_1317) );
OR2x6_ASAP7_75t_L g1318 ( .A(n_1315), .B(n_1313), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1316), .Y(n_1319) );
NOR2xp67_ASAP7_75t_L g1320 ( .A(n_1317), .B(n_1277), .Y(n_1320) );
HB1xp67_ASAP7_75t_L g1321 ( .A(n_1319), .Y(n_1321) );
AOI221xp5_ASAP7_75t_L g1322 ( .A1(n_1321), .A2(n_1318), .B1(n_1320), .B2(n_1282), .C(n_1280), .Y(n_1322) );
endmodule