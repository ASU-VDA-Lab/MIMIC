module fake_jpeg_23033_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_8),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_30),
.B(n_37),
.Y(n_54)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_4),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_2),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_3),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_27),
.C(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_17),
.B1(n_21),
.B2(n_13),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_19),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_36),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_38),
.B1(n_33),
.B2(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_13),
.B1(n_21),
.B2(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_44),
.B1(n_25),
.B2(n_32),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_28),
.A2(n_15),
.B1(n_27),
.B2(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_49),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_16),
.B1(n_18),
.B2(n_31),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_22),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_5),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_32),
.B1(n_29),
.B2(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_71),
.Y(n_82)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_5),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_75),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_43),
.B1(n_42),
.B2(n_52),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_42),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_57),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_85),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_93),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_95),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_71),
.C(n_57),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_90),
.C(n_77),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_62),
.B(n_73),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_87),
.Y(n_107)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_86),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_97),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_106),
.C(n_107),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_91),
.B(n_88),
.C(n_76),
.D(n_90),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_98),
.C(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_79),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_79),
.A3(n_86),
.B1(n_101),
.B2(n_107),
.C1(n_102),
.C2(n_77),
.Y(n_116)
);

OAI321xp33_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_103),
.A3(n_11),
.B1(n_10),
.B2(n_69),
.C(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_95),
.B1(n_78),
.B2(n_81),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_111),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_125),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_126),
.B(n_122),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_92),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_111),
.B(n_92),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_127),
.B(n_61),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_64),
.Y(n_131)
);


endmodule