module fake_jpeg_12870_n_153 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_13),
.B(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_4),
.B(n_2),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_70),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_73),
.B1(n_66),
.B2(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_1),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_3),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_67),
.C(n_48),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_6),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_6),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_83),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_65),
.B1(n_53),
.B2(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_49),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_14),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_25),
.B(n_27),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_85),
.B1(n_84),
.B2(n_65),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_96),
.B1(n_101),
.B2(n_31),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_55),
.C(n_64),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_30),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_53),
.B1(n_52),
.B2(n_47),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_63),
.B(n_47),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_17),
.B(n_18),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_63),
.B1(n_8),
.B2(n_9),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_105),
.B1(n_19),
.B2(n_20),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_10),
.CI(n_11),
.CON(n_102),
.SN(n_102)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_104),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_13),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_39),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_15),
.B1(n_16),
.B2(n_45),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_32),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_113),
.B1(n_114),
.B2(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_118),
.Y(n_131)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_122),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_125),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_95),
.C(n_102),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_97),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_129),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_133),
.B1(n_110),
.B2(n_126),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_102),
.C(n_107),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_143),
.A2(n_144),
.B(n_136),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_147),
.A2(n_136),
.B(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_148),
.B(n_149),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_131),
.C(n_139),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_140),
.A3(n_139),
.B1(n_146),
.B2(n_128),
.C1(n_137),
.C2(n_129),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_132),
.Y(n_153)
);


endmodule