module fake_jpeg_22724_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_47),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR4xp25_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_15),
.C(n_14),
.D(n_13),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_23),
.B1(n_22),
.B2(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_101)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_0),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_23),
.B1(n_22),
.B2(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_59),
.B1(n_71),
.B2(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_23),
.B1(n_31),
.B2(n_28),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_25),
.Y(n_60)
);

AO22x1_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_16),
.B1(n_29),
.B2(n_19),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_16),
.B1(n_29),
.B2(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_20),
.B1(n_18),
.B2(n_25),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_17),
.B1(n_33),
.B2(n_30),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_33),
.B(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_13),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_35),
.B1(n_26),
.B2(n_21),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_78),
.A2(n_111),
.B1(n_74),
.B2(n_77),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_84),
.B(n_51),
.Y(n_119)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_96),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_49),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_87),
.A2(n_89),
.B1(n_104),
.B2(n_74),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_103),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_98),
.B1(n_78),
.B2(n_87),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_100),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_35),
.B1(n_44),
.B2(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_46),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_33),
.B1(n_24),
.B2(n_8),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_75),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_15),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_109),
.Y(n_133)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_14),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_26),
.B1(n_14),
.B2(n_12),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_12),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_12),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_79),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_99),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_116),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_140),
.B1(n_101),
.B2(n_98),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_142),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_82),
.B(n_69),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_123),
.B(n_127),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_82),
.B(n_56),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_101),
.B1(n_108),
.B2(n_100),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_143),
.B1(n_84),
.B2(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_8),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

NAND2x1_ASAP7_75t_SL g134 ( 
.A(n_87),
.B(n_49),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_105),
.B(n_88),
.C(n_80),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_92),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_68),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_106),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_94),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_151),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_149),
.A2(n_153),
.B1(n_177),
.B2(n_137),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_157),
.B(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_159),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_90),
.B1(n_49),
.B2(n_70),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_173),
.B1(n_131),
.B2(n_137),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_81),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_156),
.A2(n_125),
.B(n_9),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_121),
.B(n_81),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_83),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_132),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_83),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_109),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_168),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_115),
.B(n_70),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_93),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_93),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_123),
.B(n_52),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_50),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_130),
.A2(n_74),
.B1(n_85),
.B2(n_72),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_128),
.B(n_48),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_134),
.B(n_143),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_77),
.B1(n_72),
.B2(n_54),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_176),
.A2(n_143),
.B1(n_134),
.B2(n_135),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_179),
.A2(n_195),
.B1(n_204),
.B2(n_173),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_136),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_205),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_136),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_194),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_164),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_120),
.C(n_124),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_191),
.C(n_201),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_120),
.C(n_124),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_198),
.B(n_180),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_149),
.A2(n_72),
.B1(n_119),
.B2(n_117),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_158),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_199),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_117),
.C(n_126),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_157),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_160),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_161),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_211),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_125),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_159),
.C(n_153),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_210),
.A2(n_146),
.B(n_178),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_156),
.B(n_91),
.CI(n_2),
.CON(n_211),
.SN(n_211)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_226),
.B1(n_236),
.B2(n_238),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_214),
.B(n_231),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_227),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_223),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_161),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_232),
.B(n_210),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_181),
.Y(n_223)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_235),
.C(n_203),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_170),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_147),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_186),
.A2(n_166),
.B(n_178),
.C(n_174),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_184),
.B1(n_197),
.B2(n_183),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_171),
.C(n_165),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_195),
.A2(n_148),
.B1(n_151),
.B2(n_162),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_172),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_237),
.B(n_239),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_180),
.A2(n_147),
.B(n_155),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_155),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_221),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_244),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_217),
.B(n_179),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_187),
.A3(n_193),
.B1(n_202),
.B2(n_197),
.C1(n_209),
.C2(n_207),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_252),
.A3(n_220),
.B1(n_231),
.B2(n_234),
.C1(n_224),
.C2(n_235),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_205),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_250),
.A2(n_251),
.B(n_236),
.Y(n_267)
);

OAI322xp33_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_146),
.A3(n_191),
.B1(n_182),
.B2(n_201),
.C1(n_211),
.C2(n_184),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_225),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_253),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_261),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_182),
.B1(n_183),
.B2(n_211),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_213),
.B1(n_219),
.B2(n_216),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_228),
.B(n_177),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_262),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_175),
.Y(n_260)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_91),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_88),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_224),
.B1(n_220),
.B2(n_234),
.Y(n_264)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_241),
.B(n_230),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_271),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_230),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_251),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_234),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_274),
.B(n_1),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g274 ( 
.A(n_244),
.B(n_234),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_240),
.A2(n_214),
.B1(n_227),
.B2(n_216),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_248),
.B1(n_249),
.B2(n_259),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_258),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_280),
.B1(n_80),
.B2(n_122),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_139),
.B1(n_122),
.B2(n_105),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_242),
.C(n_258),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_285),
.C(n_294),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_284),
.A2(n_293),
.B1(n_273),
.B2(n_271),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_257),
.C(n_262),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_288),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_246),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_264),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_292),
.B(n_274),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_9),
.B(n_139),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_122),
.C(n_2),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_281),
.C(n_276),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_1),
.C(n_3),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_301),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_282),
.A2(n_270),
.B1(n_265),
.B2(n_274),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_291),
.Y(n_311)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_267),
.B(n_277),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_300),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_284),
.A2(n_272),
.B1(n_122),
.B2(n_4),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_289),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_292),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_306),
.Y(n_316)
);

AND2x6_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_272),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_1),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_309),
.C(n_307),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_3),
.C(n_4),
.Y(n_309)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_298),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_323),
.C(n_283),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_322),
.B(n_325),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_313),
.A2(n_308),
.B(n_304),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_318),
.B(n_310),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_317),
.B(n_311),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_326),
.A2(n_327),
.B1(n_329),
.B2(n_319),
.Y(n_330)
);

AOI222xp33_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_290),
.B1(n_285),
.B2(n_309),
.C1(n_7),
.C2(n_5),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_331),
.B(n_5),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_328),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_331)
);

NOR4xp25_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_6),
.C(n_7),
.D(n_313),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_6),
.C(n_7),
.Y(n_334)
);


endmodule