module real_aes_3031_n_254 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_254);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_254;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_283;
wire n_314;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_0), .A2(n_251), .B1(n_491), .B2(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g688 ( .A(n_1), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_2), .A2(n_112), .B1(n_317), .B2(n_379), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_3), .A2(n_78), .B1(n_371), .B2(n_373), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_4), .A2(n_125), .B1(n_352), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_5), .A2(n_64), .B1(n_394), .B2(n_395), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_6), .A2(n_56), .B1(n_304), .B2(n_309), .Y(n_303) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_7), .A2(n_188), .B1(n_281), .B2(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g664 ( .A(n_7), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_8), .A2(n_163), .B1(n_442), .B2(n_472), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_9), .A2(n_82), .B1(n_329), .B2(n_365), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_10), .A2(n_27), .B1(n_316), .B2(n_321), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_11), .A2(n_12), .B1(n_352), .B2(n_354), .Y(n_351) );
XOR2x2_ASAP7_75t_L g451 ( .A(n_13), .B(n_452), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_14), .A2(n_115), .B1(n_416), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_15), .A2(n_101), .B1(n_409), .B2(n_410), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_16), .A2(n_103), .B1(n_337), .B2(n_533), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_17), .A2(n_172), .B1(n_485), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_18), .A2(n_38), .B1(n_394), .B2(n_395), .Y(n_514) );
AO22x2_ASAP7_75t_L g288 ( .A1(n_19), .A2(n_62), .B1(n_281), .B2(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_19), .B(n_663), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_20), .A2(n_59), .B1(n_317), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_21), .A2(n_197), .B1(n_381), .B2(n_382), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_22), .A2(n_152), .B1(n_427), .B2(n_429), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_23), .A2(n_36), .B1(n_344), .B2(n_347), .Y(n_343) );
AOI22xp5_ASAP7_75t_SL g539 ( .A1(n_24), .A2(n_229), .B1(n_294), .B2(n_470), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_25), .A2(n_137), .B1(n_394), .B2(n_395), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_26), .A2(n_253), .B1(n_427), .B2(n_429), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_28), .A2(n_196), .B1(n_429), .B2(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_29), .A2(n_186), .B1(n_600), .B2(n_684), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_30), .B(n_440), .Y(n_439) );
OA22x2_ASAP7_75t_L g360 ( .A1(n_31), .A2(n_361), .B1(n_362), .B2(n_389), .Y(n_360) );
INVx1_ASAP7_75t_L g389 ( .A(n_31), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_32), .A2(n_225), .B1(n_330), .B2(n_365), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g254 ( .A1(n_33), .A2(n_255), .B(n_264), .C(n_666), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_34), .A2(n_175), .B1(n_355), .B2(n_433), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_35), .A2(n_242), .B1(n_317), .B2(n_468), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_37), .A2(n_223), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_39), .A2(n_224), .B1(n_400), .B2(n_401), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_40), .B(n_388), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_41), .A2(n_176), .B1(n_367), .B2(n_486), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_42), .A2(n_238), .B1(n_294), .B2(n_684), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_43), .A2(n_245), .B1(n_409), .B2(n_410), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_44), .A2(n_170), .B1(n_642), .B2(n_643), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_45), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_46), .A2(n_205), .B1(n_382), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_47), .A2(n_67), .B1(n_700), .B2(n_701), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_48), .A2(n_168), .B1(n_457), .B2(n_459), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_49), .A2(n_202), .B1(n_600), .B2(n_601), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_50), .A2(n_158), .B1(n_397), .B2(n_398), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_51), .A2(n_57), .B1(n_384), .B2(n_386), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_52), .A2(n_110), .B1(n_384), .B2(n_442), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_53), .A2(n_243), .B1(n_317), .B2(n_322), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_54), .A2(n_72), .B1(n_304), .B2(n_309), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_55), .A2(n_116), .B1(n_317), .B2(n_379), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_58), .A2(n_63), .B1(n_337), .B2(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_60), .A2(n_147), .B1(n_459), .B2(n_581), .Y(n_580) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_61), .A2(n_65), .B1(n_240), .B2(n_633), .C1(n_634), .C2(n_635), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_66), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_68), .A2(n_226), .B1(n_608), .B2(n_609), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_69), .A2(n_198), .B1(n_329), .B2(n_331), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_70), .A2(n_199), .B1(n_397), .B2(n_398), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_71), .A2(n_92), .B1(n_375), .B2(n_376), .Y(n_374) );
AOI222xp33_ASAP7_75t_L g650 ( .A1(n_73), .A2(n_151), .B1(n_213), .B2(n_305), .C1(n_442), .C2(n_633), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_74), .A2(n_139), .B1(n_533), .B2(n_642), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_75), .A2(n_143), .B1(n_446), .B2(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g281 ( .A(n_76), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_77), .A2(n_138), .B1(n_333), .B2(n_367), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_79), .A2(n_250), .B1(n_337), .B2(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_80), .B(n_403), .Y(n_402) );
XNOR2x2_ASAP7_75t_L g390 ( .A(n_81), .B(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_83), .A2(n_236), .B1(n_371), .B2(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_84), .A2(n_217), .B1(n_400), .B2(n_401), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_85), .A2(n_150), .B1(n_406), .B2(n_407), .Y(n_524) );
OA22x2_ASAP7_75t_L g619 ( .A1(n_86), .A2(n_620), .B1(n_621), .B2(n_636), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_86), .Y(n_620) );
INVx1_ASAP7_75t_L g691 ( .A(n_87), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_88), .B(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_89), .A2(n_127), .B1(n_375), .B2(n_461), .Y(n_460) );
AO22x2_ASAP7_75t_L g589 ( .A1(n_90), .A2(n_590), .B1(n_591), .B2(n_616), .Y(n_589) );
INVx1_ASAP7_75t_L g616 ( .A(n_90), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_91), .B(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_93), .A2(n_149), .B1(n_535), .B2(n_536), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_94), .A2(n_174), .B1(n_375), .B2(n_376), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_95), .A2(n_114), .B1(n_375), .B2(n_376), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_96), .A2(n_122), .B1(n_446), .B2(n_447), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_97), .A2(n_219), .B1(n_336), .B2(n_340), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_98), .A2(n_128), .B1(n_614), .B2(n_615), .Y(n_613) );
INVx1_ASAP7_75t_SL g282 ( .A(n_99), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_99), .B(n_124), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_100), .A2(n_208), .B1(n_355), .B2(n_455), .Y(n_563) );
INVx2_ASAP7_75t_L g261 ( .A(n_102), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_104), .A2(n_159), .B1(n_493), .B2(n_611), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_105), .A2(n_189), .B1(n_457), .B2(n_536), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_106), .A2(n_145), .B1(n_317), .B2(n_322), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_107), .A2(n_220), .B1(n_367), .B2(n_368), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_108), .A2(n_118), .B1(n_382), .B2(n_446), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_109), .A2(n_244), .B1(n_468), .B2(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_111), .B(n_594), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_113), .A2(n_221), .B1(n_356), .B2(n_371), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_117), .A2(n_218), .B1(n_340), .B2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_119), .A2(n_212), .B1(n_499), .B2(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_120), .A2(n_179), .B1(n_707), .B2(n_708), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_121), .A2(n_216), .B1(n_373), .B2(n_433), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_123), .A2(n_203), .B1(n_316), .B2(n_470), .Y(n_682) );
AO22x2_ASAP7_75t_L g284 ( .A1(n_124), .A2(n_200), .B1(n_281), .B2(n_285), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_126), .A2(n_210), .B1(n_305), .B2(n_442), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_129), .B(n_388), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_130), .A2(n_191), .B1(n_489), .B2(n_583), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_131), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g500 ( .A1(n_132), .A2(n_239), .B1(n_442), .B2(n_472), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_133), .A2(n_185), .B1(n_406), .B2(n_407), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_134), .A2(n_246), .B1(n_352), .B2(n_354), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_135), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_136), .A2(n_171), .B1(n_340), .B2(n_455), .Y(n_454) );
OA22x2_ASAP7_75t_L g269 ( .A1(n_140), .A2(n_270), .B1(n_271), .B2(n_357), .Y(n_269) );
INVx1_ASAP7_75t_L g357 ( .A(n_140), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_141), .A2(n_156), .B1(n_365), .B2(n_433), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_142), .A2(n_148), .B1(n_356), .B2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_144), .A2(n_180), .B1(n_331), .B2(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g283 ( .A(n_146), .Y(n_283) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_153), .A2(n_215), .B1(n_294), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_154), .A2(n_164), .B1(n_415), .B2(n_416), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_155), .B(n_438), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_157), .A2(n_162), .B1(n_412), .B2(n_413), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_160), .A2(n_178), .B1(n_485), .B2(n_486), .Y(n_484) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_161), .B(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_165), .A2(n_248), .B1(n_406), .B2(n_407), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_166), .A2(n_230), .B1(n_412), .B2(n_413), .Y(n_520) );
XNOR2x1_ASAP7_75t_L g548 ( .A(n_167), .B(n_549), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_169), .A2(n_201), .B1(n_375), .B2(n_461), .Y(n_640) );
INVx1_ASAP7_75t_L g566 ( .A(n_173), .Y(n_566) );
AOI22xp33_ASAP7_75t_SL g498 ( .A1(n_177), .A2(n_183), .B1(n_294), .B2(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_181), .A2(n_249), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_182), .A2(n_193), .B1(n_294), .B2(n_299), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_184), .B(n_275), .Y(n_473) );
XNOR2x1_ASAP7_75t_L g481 ( .A(n_187), .B(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_190), .A2(n_207), .B1(n_398), .B2(n_512), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_192), .A2(n_231), .B1(n_349), .B2(n_427), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_194), .A2(n_252), .B1(n_466), .B2(n_468), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_195), .A2(n_209), .B1(n_415), .B2(n_678), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_204), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_206), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g660 ( .A(n_206), .Y(n_660) );
INVx1_ASAP7_75t_L g258 ( .A(n_211), .Y(n_258) );
AND2x2_ASAP7_75t_R g693 ( .A(n_211), .B(n_660), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_214), .B(n_275), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_222), .B(n_274), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_227), .A2(n_237), .B1(n_305), .B2(n_310), .Y(n_540) );
INVxp67_ASAP7_75t_L g263 ( .A(n_228), .Y(n_263) );
INVx1_ASAP7_75t_L g687 ( .A(n_232), .Y(n_687) );
XNOR2xp5_ASAP7_75t_L g695 ( .A(n_233), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g718 ( .A(n_233), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_234), .B(n_442), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_235), .A2(n_247), .B1(n_328), .B2(n_331), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_241), .B(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2x1_ASAP7_75t_R g256 ( .A(n_257), .B(n_259), .Y(n_256) );
OR2x2_ASAP7_75t_L g717 ( .A(n_257), .B(n_260), .Y(n_717) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_258), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_587), .B1(n_655), .B2(n_656), .C(n_657), .Y(n_264) );
INVx1_ASAP7_75t_L g655 ( .A(n_265), .Y(n_655) );
XOR2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_478), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B1(n_418), .B2(n_419), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AO22x2_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_358), .B1(n_359), .B2(n_417), .Y(n_268) );
INVx2_ASAP7_75t_L g417 ( .A(n_269), .Y(n_417) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_326), .Y(n_271) );
NAND4xp25_ASAP7_75t_SL g272 ( .A(n_273), .B(n_293), .C(n_303), .D(n_315), .Y(n_272) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx4_ASAP7_75t_SL g388 ( .A(n_276), .Y(n_388) );
INVx4_ASAP7_75t_SL g403 ( .A(n_276), .Y(n_403) );
INVx3_ASAP7_75t_SL g503 ( .A(n_276), .Y(n_503) );
INVx6_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_286), .Y(n_277) );
AND2x4_ASAP7_75t_L g301 ( .A(n_278), .B(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_L g323 ( .A(n_278), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g395 ( .A(n_278), .B(n_324), .Y(n_395) );
AND2x2_ASAP7_75t_L g398 ( .A(n_278), .B(n_302), .Y(n_398) );
AND2x4_ASAP7_75t_L g438 ( .A(n_278), .B(n_286), .Y(n_438) );
AND2x2_ASAP7_75t_L g513 ( .A(n_278), .B(n_302), .Y(n_513) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_284), .Y(n_278) );
INVx2_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
AND2x2_ASAP7_75t_L g307 ( .A(n_279), .B(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_279), .Y(n_314) );
OAI22x1_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B1(n_282), .B2(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g285 ( .A(n_281), .Y(n_285) );
INVx2_ASAP7_75t_L g289 ( .A(n_281), .Y(n_289) );
INVx1_ASAP7_75t_L g292 ( .A(n_281), .Y(n_292) );
AND2x2_ASAP7_75t_L g297 ( .A(n_284), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
BUFx2_ASAP7_75t_L g350 ( .A(n_284), .Y(n_350) );
AND2x4_ASAP7_75t_L g330 ( .A(n_286), .B(n_307), .Y(n_330) );
AND2x4_ASAP7_75t_L g339 ( .A(n_286), .B(n_334), .Y(n_339) );
AND2x2_ASAP7_75t_L g353 ( .A(n_286), .B(n_297), .Y(n_353) );
AND2x6_ASAP7_75t_L g406 ( .A(n_286), .B(n_297), .Y(n_406) );
AND2x2_ASAP7_75t_L g409 ( .A(n_286), .B(n_307), .Y(n_409) );
AND2x2_ASAP7_75t_L g522 ( .A(n_286), .B(n_334), .Y(n_522) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g296 ( .A(n_288), .B(n_290), .Y(n_296) );
AND2x2_ASAP7_75t_L g313 ( .A(n_288), .B(n_291), .Y(n_313) );
INVx1_ASAP7_75t_L g320 ( .A(n_288), .Y(n_320) );
INVxp67_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_320), .Y(n_319) );
BUFx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g381 ( .A(n_295), .Y(n_381) );
BUFx3_ASAP7_75t_L g446 ( .A(n_295), .Y(n_446) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_295), .Y(n_711) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g306 ( .A(n_296), .B(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g356 ( .A(n_296), .B(n_334), .Y(n_356) );
AND2x2_ASAP7_75t_L g397 ( .A(n_296), .B(n_297), .Y(n_397) );
AND2x4_ASAP7_75t_L g400 ( .A(n_296), .B(n_307), .Y(n_400) );
AND2x2_ASAP7_75t_L g416 ( .A(n_296), .B(n_334), .Y(n_416) );
AND2x2_ASAP7_75t_L g512 ( .A(n_296), .B(n_297), .Y(n_512) );
AND2x2_ASAP7_75t_L g346 ( .A(n_297), .B(n_319), .Y(n_346) );
AND2x2_ASAP7_75t_L g412 ( .A(n_297), .B(n_319), .Y(n_412) );
AND2x4_ASAP7_75t_L g334 ( .A(n_298), .B(n_308), .Y(n_334) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g382 ( .A(n_300), .Y(n_382) );
INVx2_ASAP7_75t_L g447 ( .A(n_300), .Y(n_447) );
INVx1_ASAP7_75t_L g470 ( .A(n_300), .Y(n_470) );
INVx2_ASAP7_75t_SL g499 ( .A(n_300), .Y(n_499) );
INVx2_ASAP7_75t_L g552 ( .A(n_300), .Y(n_552) );
INVx6_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_SL g686 ( .A(n_304), .Y(n_686) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g385 ( .A(n_306), .Y(n_385) );
BUFx5_ASAP7_75t_L g472 ( .A(n_306), .Y(n_472) );
AND2x2_ASAP7_75t_L g318 ( .A(n_307), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g394 ( .A(n_307), .B(n_319), .Y(n_394) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g386 ( .A(n_311), .Y(n_386) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx12f_ASAP7_75t_L g442 ( .A(n_312), .Y(n_442) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x4_ASAP7_75t_L g333 ( .A(n_313), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g349 ( .A(n_313), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_SL g401 ( .A(n_313), .B(n_314), .Y(n_401) );
AND2x4_ASAP7_75t_L g410 ( .A(n_313), .B(n_334), .Y(n_410) );
AND2x4_ASAP7_75t_L g413 ( .A(n_313), .B(n_350), .Y(n_413) );
AND2x2_ASAP7_75t_SL g635 ( .A(n_313), .B(n_314), .Y(n_635) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx3_ASAP7_75t_L g467 ( .A(n_318), .Y(n_467) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_318), .Y(n_554) );
AND2x4_ASAP7_75t_L g342 ( .A(n_319), .B(n_334), .Y(n_342) );
AND2x6_ASAP7_75t_L g407 ( .A(n_319), .B(n_334), .Y(n_407) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_320), .Y(n_325) );
BUFx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g379 ( .A(n_323), .Y(n_379) );
BUFx4f_ASAP7_75t_L g468 ( .A(n_323), .Y(n_468) );
INVx1_ASAP7_75t_L g543 ( .A(n_323), .Y(n_543) );
INVx2_ASAP7_75t_L g603 ( .A(n_323), .Y(n_603) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND4xp25_ASAP7_75t_L g326 ( .A(n_327), .B(n_335), .C(n_343), .D(n_351), .Y(n_326) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx3_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
INVx6_ASAP7_75t_L g458 ( .A(n_330), .Y(n_458) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_SL g459 ( .A(n_332), .Y(n_459) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx3_ASAP7_75t_L g365 ( .A(n_333), .Y(n_365) );
BUFx3_ASAP7_75t_L g536 ( .A(n_333), .Y(n_536) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx4_ASAP7_75t_L g415 ( .A(n_338), .Y(n_415) );
INVx3_ASAP7_75t_L g433 ( .A(n_338), .Y(n_433) );
INVx2_ASAP7_75t_SL g495 ( .A(n_338), .Y(n_495) );
INVx2_ASAP7_75t_L g606 ( .A(n_338), .Y(n_606) );
INVx3_ASAP7_75t_SL g642 ( .A(n_338), .Y(n_642) );
INVx8_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g373 ( .A(n_341), .Y(n_373) );
INVx1_ASAP7_75t_SL g489 ( .A(n_341), .Y(n_489) );
INVx2_ASAP7_75t_L g533 ( .A(n_341), .Y(n_533) );
INVx2_ASAP7_75t_L g609 ( .A(n_341), .Y(n_609) );
INVx2_ASAP7_75t_L g628 ( .A(n_341), .Y(n_628) );
INVx8_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_346), .Y(n_375) );
INVx2_ASAP7_75t_L g428 ( .A(n_346), .Y(n_428) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
INVx2_ASAP7_75t_L g429 ( .A(n_348), .Y(n_429) );
INVx5_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g461 ( .A(n_349), .Y(n_461) );
BUFx2_ASAP7_75t_L g493 ( .A(n_349), .Y(n_493) );
BUFx2_ASAP7_75t_L g701 ( .A(n_349), .Y(n_701) );
BUFx3_ASAP7_75t_L g608 ( .A(n_352), .Y(n_608) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx3_ASAP7_75t_L g372 ( .A(n_353), .Y(n_372) );
BUFx2_ASAP7_75t_L g455 ( .A(n_353), .Y(n_455) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g571 ( .A(n_355), .Y(n_571) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g369 ( .A(n_356), .Y(n_369) );
BUFx3_ASAP7_75t_L g486 ( .A(n_356), .Y(n_486) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_356), .Y(n_643) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
XNOR2x1_ASAP7_75t_L g359 ( .A(n_360), .B(n_390), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_363), .B(n_377), .Y(n_362) );
NAND4xp25_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .C(n_370), .D(n_374), .Y(n_363) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_365), .Y(n_615) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g463 ( .A(n_369), .Y(n_463) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_SL g488 ( .A(n_372), .Y(n_488) );
INVx2_ASAP7_75t_SL g583 ( .A(n_372), .Y(n_583) );
INVx3_ASAP7_75t_L g676 ( .A(n_372), .Y(n_676) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_375), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .C(n_383), .D(n_387), .Y(n_377) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g440 ( .A(n_385), .Y(n_440) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_404), .Y(n_391) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_393), .B(n_396), .C(n_399), .D(n_402), .Y(n_392) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_400), .Y(n_634) );
BUFx2_ASAP7_75t_L g594 ( .A(n_403), .Y(n_594) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .C(n_411), .D(n_414), .Y(n_404) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_415), .Y(n_581) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AO22x1_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_449), .B1(n_474), .B2(n_475), .Y(n_419) );
INVx1_ASAP7_75t_L g474 ( .A(n_420), .Y(n_474) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
XOR2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_448), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_434), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_430), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g492 ( .A(n_428), .Y(n_492) );
INVx1_ASAP7_75t_L g612 ( .A(n_428), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_443), .Y(n_434) );
OAI211xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B(n_439), .C(n_441), .Y(n_435) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g633 ( .A(n_438), .Y(n_633) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_440), .Y(n_708) );
INVx2_ASAP7_75t_L g690 ( .A(n_442), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g597 ( .A(n_446), .Y(n_597) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g477 ( .A(n_451), .Y(n_477) );
NOR2xp67_ASAP7_75t_L g452 ( .A(n_453), .B(n_464), .Y(n_452) );
NAND4xp25_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .C(n_460), .D(n_462), .Y(n_453) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g485 ( .A(n_458), .Y(n_485) );
INVx3_ASAP7_75t_L g535 ( .A(n_458), .Y(n_535) );
INVx1_ASAP7_75t_SL g614 ( .A(n_458), .Y(n_614) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .C(n_471), .D(n_473), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
XNOR2x1_ASAP7_75t_L g478 ( .A(n_479), .B(n_546), .Y(n_478) );
AO22x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_504), .B2(n_505), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_496), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .C(n_490), .D(n_494), .Y(n_483) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .C(n_500), .D(n_501), .Y(n_496) );
INVx3_ASAP7_75t_L g689 ( .A(n_502), .Y(n_689) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OA22x2_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_527), .B2(n_545), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
XOR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_526), .Y(n_507) );
NAND2x1_ASAP7_75t_SL g508 ( .A(n_509), .B(n_518), .Y(n_508) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_510), .B(n_515), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_514), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
NOR2x1_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_SL g545 ( .A(n_527), .Y(n_545) );
XNOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_544), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_537), .Y(n_528) );
NAND4xp25_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .C(n_532), .D(n_534), .Y(n_529) );
NAND4xp25_ASAP7_75t_SL g537 ( .A(n_538), .B(n_539), .C(n_540), .D(n_541), .Y(n_537) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_564), .B1(n_585), .B2(n_586), .Y(n_547) );
INVx2_ASAP7_75t_L g586 ( .A(n_548), .Y(n_586) );
NAND4xp75_ASAP7_75t_L g549 ( .A(n_550), .B(n_555), .C(n_558), .D(n_561), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
BUFx6f_ASAP7_75t_SL g600 ( .A(n_554), .Y(n_600) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g585 ( .A(n_564), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B1(n_573), .B2(n_584), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_568), .B(n_574), .C(n_579), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_579), .Y(n_573) );
NAND4xp25_ASAP7_75t_SL g574 ( .A(n_575), .B(n_576), .C(n_577), .D(n_578), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx1_ASAP7_75t_L g656 ( .A(n_587), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_589), .B1(n_617), .B2(n_654), .Y(n_587) );
INVx4_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_604), .Y(n_591) );
NAND4xp25_ASAP7_75t_SL g592 ( .A(n_593), .B(n_595), .C(n_598), .D(n_599), .Y(n_592) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g684 ( .A(n_603), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .C(n_610), .D(n_613), .Y(n_604) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g654 ( .A(n_617), .Y(n_654) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_637), .B1(n_652), .B2(n_653), .Y(n_618) );
INVx1_ASAP7_75t_L g652 ( .A(n_619), .Y(n_652) );
INVx2_ASAP7_75t_L g636 ( .A(n_621), .Y(n_636) );
NAND4xp75_ASAP7_75t_L g621 ( .A(n_622), .B(n_625), .C(n_629), .D(n_632), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_SL g653 ( .A(n_637), .Y(n_653) );
XOR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_651), .Y(n_637) );
NAND4xp75_ASAP7_75t_L g638 ( .A(n_639), .B(n_644), .C(n_647), .D(n_650), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx2_ASAP7_75t_L g679 ( .A(n_643), .Y(n_679) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_659), .B(n_662), .Y(n_714) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
OAI222xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_692), .B1(n_694), .B2(n_712), .C1(n_715), .C2(n_718), .Y(n_666) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_680), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_685), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
OAI222xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_688), .B2(n_689), .C1(n_690), .C2(n_691), .Y(n_685) );
INVx2_ASAP7_75t_L g707 ( .A(n_690), .Y(n_707) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_697), .B(n_704), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .C(n_702), .D(n_703), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .C(n_709), .D(n_710), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
CKINVDCx6p67_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_716), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
endmodule