module real_jpeg_32031_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_578;
wire n_332;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_268;
wire n_597;
wire n_42;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_0),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_0),
.Y(n_269)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_0),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_22),
.Y(n_18)
);

CKINVDCx11_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_2),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_3),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_3),
.B(n_156),
.Y(n_256)
);

NAND2x1_ASAP7_75t_L g275 ( 
.A(n_3),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_3),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_3),
.B(n_356),
.Y(n_355)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_3),
.B(n_164),
.C(n_462),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_3),
.B(n_467),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_3),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_3),
.B(n_462),
.Y(n_482)
);

NAND3xp33_ASAP7_75t_SL g545 ( 
.A(n_3),
.B(n_164),
.C(n_462),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_5),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_6),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_6),
.Y(n_464)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_6),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_7),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_7),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_7),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_SL g334 ( 
.A(n_7),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_7),
.B(n_424),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_7),
.B(n_218),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_7),
.B(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_7),
.B(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_8),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_8),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_8),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_8),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_8),
.B(n_496),
.Y(n_495)
);

BUFx2_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_9),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_9),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_9),
.B(n_104),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_9),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_9),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_9),
.B(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_9),
.B(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_10),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_11),
.Y(n_339)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_12),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_13),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_14),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_14),
.B(n_218),
.Y(n_217)
);

AOI22x1_ASAP7_75t_L g340 ( 
.A1(n_14),
.A2(n_15),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

NAND2x1_ASAP7_75t_L g265 ( 
.A(n_15),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_15),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_15),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_15),
.B(n_421),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_15),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_15),
.B(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_15),
.B(n_523),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_16),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_16),
.B(n_128),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_16),
.B(n_111),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_16),
.B(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_17),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_17),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_17),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_SL g329 ( 
.A(n_17),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_17),
.B(n_382),
.Y(n_381)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_616),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_131),
.B(n_288),
.C(n_596),
.D(n_615),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_183),
.Y(n_24)
);

OAI211xp5_ASAP7_75t_L g596 ( 
.A1(n_25),
.A2(n_597),
.B(n_600),
.C(n_602),
.Y(n_596)
);

NOR2xp67_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_115),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_90),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_27),
.B(n_90),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_56),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_28),
.B(n_56),
.C(n_90),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_46),
.C(n_51),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_29),
.B(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.C(n_42),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_30),
.A2(n_31),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_30),
.B(n_127),
.C(n_131),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_30),
.A2(n_31),
.B1(n_303),
.B2(n_416),
.Y(n_415)
);

CKINVDCx11_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_31),
.B(n_303),
.C(n_306),
.Y(n_302)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_33),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_33),
.Y(n_517)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_34),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_34),
.A2(n_178),
.B1(n_609),
.B2(n_610),
.Y(n_608)
);

NAND2x1_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_40),
.Y(n_167)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_40),
.Y(n_358)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_41),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_42),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_42),
.A2(n_63),
.B1(n_72),
.B2(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_42),
.A2(n_63),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_42),
.A2(n_63),
.B1(n_312),
.B2(n_317),
.Y(n_311)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NOR2x1_ASAP7_75t_R g107 ( 
.A(n_47),
.B(n_108),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_47),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_47),
.B(n_226),
.Y(n_234)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_54),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_55),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_55),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_78),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_58),
.B(n_78),
.C(n_613),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_62),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.C(n_72),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_63),
.B(n_312),
.C(n_318),
.Y(n_359)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_66),
.B(n_127),
.C(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_67),
.B(n_135),
.Y(n_206)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_71),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_71),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_73),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_72),
.A2(n_73),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_73),
.B(n_84),
.C(n_88),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_74),
.B(n_265),
.C(n_267),
.Y(n_264)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_75),
.Y(n_451)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_76),
.Y(n_356)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_77),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_77),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

XOR2x2_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_79),
.B(n_146),
.C(n_148),
.Y(n_179)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_83),
.B(n_212),
.C(n_216),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_83),
.A2(n_84),
.B1(n_153),
.B2(n_154),
.Y(n_610)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_84),
.B(n_260),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_SL g615 ( 
.A(n_84),
.B(n_154),
.C(n_178),
.Y(n_615)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_87),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.C(n_112),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2x1_ASAP7_75t_L g181 ( 
.A(n_92),
.B(n_182),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_95),
.B(n_113),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_103),
.C(n_107),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_96),
.A2(n_97),
.B1(n_103),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_98),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_98),
.B(n_395),
.Y(n_394)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_103),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_103),
.B(n_164),
.C(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_104),
.Y(n_305)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2x1_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_115),
.B(n_601),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_173),
.C(n_181),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_116),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_117),
.A2(n_174),
.B(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_150),
.C(n_169),
.Y(n_117)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_133),
.C(n_140),
.Y(n_118)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_119),
.Y(n_285)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_122),
.Y(n_131)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_124),
.Y(n_266)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_127),
.B(n_267),
.Y(n_379)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_132),
.B(n_206),
.Y(n_205)
);

XOR2x2_ASAP7_75t_L g458 ( 
.A(n_132),
.B(n_267),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_133),
.A2(n_134),
.B1(n_140),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_138),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_140),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_141)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_142),
.A2(n_148),
.B1(n_255),
.B2(n_256),
.Y(n_352)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_144),
.Y(n_426)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_145),
.Y(n_309)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g249 ( 
.A(n_148),
.B(n_250),
.C(n_254),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_148),
.A2(n_250),
.B(n_254),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_150),
.A2(n_151),
.B1(n_170),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_159),
.B(n_168),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_155),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_153),
.B(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_153),
.A2(n_154),
.B1(n_225),
.B2(n_234),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_154),
.A2(n_225),
.B(n_228),
.C(n_233),
.Y(n_224)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_155),
.Y(n_223)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.C(n_166),
.Y(n_159)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_160),
.A2(n_208),
.B1(n_354),
.B2(n_355),
.Y(n_404)
);

OR2x2_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_161),
.Y(n_468)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_162),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_166),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_164),
.A2(n_229),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_164),
.Y(n_245)
);

XNOR2x2_ASAP7_75t_L g481 ( 
.A(n_164),
.B(n_482),
.Y(n_481)
);

INVx8_ASAP7_75t_L g396 ( 
.A(n_165),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_172),
.A2(n_243),
.B(n_246),
.Y(n_242)
);

OAI211xp5_ASAP7_75t_L g246 ( 
.A1(n_172),
.A2(n_229),
.B(n_245),
.C(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.C(n_180),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_235),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_184),
.A2(n_598),
.B(n_599),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_L g599 ( 
.A(n_185),
.B(n_192),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B(n_190),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.C(n_201),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_199),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_221),
.C(n_224),
.Y(n_202)
);

XOR2x1_ASAP7_75t_SL g286 ( 
.A(n_203),
.B(n_287),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.C(n_210),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_205),
.B(n_211),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_207),
.B(n_570),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_208),
.B(n_354),
.C(n_357),
.Y(n_353)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_220),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_221),
.B(n_224),
.Y(n_287)
);

INVx5_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_229),
.B(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_232),
.Y(n_320)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_232),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_236),
.B(n_238),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_281),
.C(n_286),
.Y(n_238)
);

INVxp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_240),
.B(n_282),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_261),
.C(n_278),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_241),
.B(n_567),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.C(n_258),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_242),
.Y(n_368)
);

XNOR2x1_ASAP7_75t_L g417 ( 
.A(n_244),
.B(n_298),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_248),
.B(n_259),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_255),
.B(n_257),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_250),
.B(n_254),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_262),
.B(n_279),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.C(n_275),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_264),
.B(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_265),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_268),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_271),
.A2(n_272),
.B1(n_275),
.B2(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_275),
.Y(n_366)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g577 ( 
.A(n_286),
.B(n_578),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_587),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_437),
.C(n_562),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_409),
.Y(n_290)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_291),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_371),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_292),
.B(n_371),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_347),
.B2(n_370),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_293),
.B(n_581),
.C(n_582),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_322),
.C(n_326),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_295),
.B(n_373),
.Y(n_372)
);

AO21x1_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_310),
.B(n_321),
.Y(n_295)
);

NAND2xp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_302),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_297),
.B(n_302),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_299),
.B(n_507),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_299),
.B(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_303),
.Y(n_416)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_SL g414 ( 
.A(n_306),
.B(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_309),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_310),
.B(n_434),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_318),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx4f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_322),
.B(n_326),
.Y(n_373)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_340),
.B2(n_346),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_334),
.Y(n_328)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_329),
.Y(n_362)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_340),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_362),
.C(n_363),
.Y(n_361)
);

INVx3_ASAP7_75t_SL g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_342),
.B(n_477),
.Y(n_476)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_346),
.A2(n_394),
.B(n_397),
.Y(n_393)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_347),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_367),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_348),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_360),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g572 ( 
.A(n_349),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.C(n_359),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_350),
.B(n_353),
.Y(n_408)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_361),
.Y(n_573)
);

INVxp33_ASAP7_75t_L g574 ( 
.A(n_364),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_367),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.C(n_405),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_372),
.B(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_375),
.B(n_406),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_393),
.C(n_401),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_377),
.B(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.C(n_386),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_378),
.A2(n_379),
.B1(n_547),
.B2(n_548),
.Y(n_546)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_380),
.A2(n_381),
.B1(n_387),
.B2(n_388),
.Y(n_548)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_385),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_402),
.Y(n_412)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

INVxp33_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_435),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_410),
.B(n_435),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.C(n_432),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_411),
.B(n_555),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_413),
.A2(n_433),
.B1(n_556),
.B2(n_557),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_413),
.Y(n_557)
);

MAJx2_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.C(n_418),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_414),
.B(n_539),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_417),
.A2(n_418),
.B1(n_540),
.B2(n_541),
.Y(n_539)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_417),
.Y(n_541)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_418),
.Y(n_540)
);

MAJx2_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_423),
.C(n_427),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_420),
.B1(n_427),
.B2(n_428),
.Y(n_446)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_446),
.Y(n_445)
);

INVx3_ASAP7_75t_SL g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_433),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_552),
.B(n_561),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_535),
.B(n_551),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_483),
.B(n_534),
.Y(n_440)
);

NAND3xp33_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_469),
.C(n_470),
.Y(n_441)
);

AOI21xp33_ASAP7_75t_SL g534 ( 
.A1(n_442),
.A2(n_469),
.B(n_470),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_456),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_444),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_457),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_445),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_447),
.B(n_456),
.C(n_550),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_452),
.C(n_453),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_448),
.A2(n_449),
.B1(n_452),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_452),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_472),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_454),
.B(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_458),
.B(n_465),
.C(n_545),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_R g560 ( 
.A(n_458),
.B(n_465),
.C(n_545),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_461),
.B1(n_465),
.B2(n_466),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_474),
.C(n_481),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_471),
.B(n_498),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_474),
.A2(n_475),
.B1(n_481),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_476),
.A2(n_478),
.B1(n_479),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_476),
.Y(n_488)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_481),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_484),
.A2(n_500),
.B(n_533),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_497),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_485),
.B(n_497),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_489),
.C(n_495),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_486),
.A2(n_487),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_490),
.B(n_495),
.Y(n_529)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_527),
.B(n_532),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_512),
.B(n_526),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_506),
.Y(n_502)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_518),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_518),
.Y(n_526)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_521),
.B1(n_522),
.B2(n_525),
.Y(n_518)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_519),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_525),
.Y(n_531)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_531),
.Y(n_532)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_529),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_549),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_549),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_538),
.B1(n_542),
.B2(n_543),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_559),
.C(n_560),
.Y(n_558)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_546),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_546),
.Y(n_559)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_554),
.B(n_558),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_554),
.B(n_558),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_562),
.A2(n_588),
.B(n_592),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_563),
.A2(n_576),
.B1(n_579),
.B2(n_583),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_L g593 ( 
.A(n_564),
.B(n_577),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_564),
.B(n_577),
.Y(n_595)
);

OAI22x1_ASAP7_75t_L g564 ( 
.A1(n_565),
.A2(n_568),
.B1(n_571),
.B2(n_575),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_566),
.B(n_569),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_569),
.B(n_571),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_569),
.Y(n_575)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_571),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_573),
.C(n_574),
.Y(n_571)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_580),
.B(n_584),
.Y(n_594)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_585),
.B(n_586),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_589),
.A2(n_590),
.B(n_591),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_593),
.A2(n_594),
.B(n_595),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_603),
.B(n_606),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_604),
.B(n_614),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_612),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_606),
.A2(n_607),
.B1(n_608),
.B2(n_611),
.Y(n_605)
);

CKINVDCx11_ASAP7_75t_R g606 ( 
.A(n_607),
.Y(n_606)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_608),
.Y(n_611)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);


endmodule