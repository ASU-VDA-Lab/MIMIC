module fake_jpeg_9080_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_24),
.B(n_0),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_35),
.B1(n_20),
.B2(n_25),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_48),
.B1(n_46),
.B2(n_17),
.Y(n_86)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_68),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_27),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_73),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_75),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_35),
.B1(n_17),
.B2(n_27),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_85),
.B1(n_86),
.B2(n_29),
.Y(n_111)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_15),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_42),
.B1(n_35),
.B2(n_40),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_88),
.B1(n_98),
.B2(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_82),
.B(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_18),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_48),
.B1(n_46),
.B2(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_18),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_37),
.B1(n_43),
.B2(n_39),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_40),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_96),
.C(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_90),
.B(n_97),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_93),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_30),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_27),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_69),
.A2(n_43),
.B1(n_18),
.B2(n_26),
.Y(n_98)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_59),
.B1(n_65),
.B2(n_54),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_50),
.B(n_57),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_69),
.B1(n_68),
.B2(n_50),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_81),
.B1(n_74),
.B2(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_122),
.Y(n_138)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_106),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_111),
.B1(n_115),
.B2(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_109),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_19),
.B1(n_33),
.B2(n_24),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_116),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_28),
.C(n_29),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_19),
.B1(n_28),
.B2(n_36),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_120),
.A3(n_102),
.B1(n_129),
.B2(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_43),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_66),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_129),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_66),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_147),
.Y(n_164)
);

AO21x2_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_98),
.B(n_88),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_91),
.B1(n_64),
.B2(n_99),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_143),
.B1(n_151),
.B2(n_116),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_79),
.B(n_36),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_144),
.B(n_148),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_101),
.B(n_103),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_157),
.B(n_127),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_88),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_144),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_145),
.B1(n_117),
.B2(n_126),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_103),
.A2(n_98),
.B1(n_88),
.B2(n_94),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_98),
.Y(n_144)
);

INVx5_ASAP7_75t_SL g146 ( 
.A(n_124),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_146),
.A2(n_152),
.B1(n_158),
.B2(n_110),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_67),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_154),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_106),
.B1(n_117),
.B2(n_121),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_23),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_26),
.C(n_23),
.Y(n_167)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_36),
.B(n_64),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_109),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_159),
.A2(n_158),
.B(n_146),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_64),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_167),
.C(n_155),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_162),
.B(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_174),
.B1(n_176),
.B2(n_189),
.Y(n_198)
);

AOI22x1_ASAP7_75t_SL g212 ( 
.A1(n_170),
.A2(n_147),
.B1(n_95),
.B2(n_152),
.Y(n_212)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_175),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_113),
.B1(n_121),
.B2(n_126),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_131),
.A2(n_117),
.B1(n_21),
.B2(n_26),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_136),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_130),
.C(n_154),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_22),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_180),
.B(n_190),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_131),
.A2(n_21),
.B1(n_23),
.B2(n_51),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_21),
.B1(n_64),
.B2(n_51),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_184),
.B(n_147),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx6_ASAP7_75t_SL g195 ( 
.A(n_185),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_131),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_133),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_189),
.A2(n_191),
.B1(n_92),
.B2(n_110),
.Y(n_217)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_131),
.A2(n_70),
.B1(n_80),
.B2(n_93),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_137),
.B(n_149),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_192),
.A2(n_196),
.B(n_199),
.Y(n_237)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_203),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_142),
.B(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_179),
.A2(n_142),
.B(n_148),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_200),
.A2(n_208),
.B(n_30),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_205),
.C(n_183),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_164),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_132),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_135),
.B(n_143),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_173),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_171),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_218),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_170),
.B(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_22),
.Y(n_216)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_186),
.B1(n_163),
.B2(n_172),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_159),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_234),
.C(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_SL g270 ( 
.A1(n_229),
.A2(n_240),
.B(n_222),
.C(n_219),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_161),
.Y(n_230)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_232),
.B(n_196),
.Y(n_249)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_195),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_168),
.B1(n_185),
.B2(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_243),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_211),
.A2(n_95),
.B1(n_168),
.B2(n_30),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_240),
.B(n_211),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_32),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_32),
.B1(n_31),
.B2(n_2),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_199),
.A2(n_31),
.B1(n_1),
.B2(n_3),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_244),
.B(n_220),
.Y(n_257)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_248),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_0),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_247),
.Y(n_255)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_262),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_R g252 ( 
.A1(n_229),
.A2(n_212),
.B1(n_192),
.B2(n_201),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_241),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_207),
.B(n_200),
.Y(n_253)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_257),
.B(n_259),
.Y(n_283)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_220),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_266),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_202),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_263),
.A2(n_270),
.B1(n_245),
.B2(n_239),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_216),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_197),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_207),
.C(n_214),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_233),
.C(n_226),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_227),
.B1(n_217),
.B2(n_242),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_273),
.A2(n_277),
.B1(n_268),
.B2(n_263),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_232),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_282),
.C(n_284),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_228),
.B1(n_244),
.B2(n_243),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_237),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_287),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_270),
.Y(n_303)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_245),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_226),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_282),
.C(n_269),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_197),
.Y(n_287)
);

OAI22x1_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_251),
.B1(n_259),
.B2(n_253),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_270),
.B(n_278),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_298),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_258),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_297),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_255),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_251),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_250),
.C(n_268),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_292),
.C(n_290),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_294),
.B1(n_289),
.B2(n_279),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_286),
.B(n_231),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_302),
.B(n_287),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_270),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_313),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_7),
.B1(n_15),
.B2(n_13),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_299),
.A2(n_300),
.B1(n_297),
.B2(n_275),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_308),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_316),
.C(n_13),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_315),
.C(n_13),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_276),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_16),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_274),
.B(n_8),
.Y(n_315)
);

OAI21x1_ASAP7_75t_SL g316 ( 
.A1(n_295),
.A2(n_8),
.B(n_15),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_320),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_7),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_322),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_16),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_323),
.A2(n_304),
.B(n_309),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_310),
.C(n_11),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_11),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_10),
.B1(n_9),
.B2(n_3),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_332),
.A3(n_324),
.B1(n_317),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_315),
.B1(n_310),
.B2(n_311),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_330),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_1),
.B(n_4),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_10),
.B1(n_9),
.B2(n_3),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_333),
.B(n_335),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_336),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_328),
.C(n_326),
.Y(n_338)
);

AOI322xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_329),
.A3(n_334),
.B1(n_331),
.B2(n_6),
.C1(n_1),
.C2(n_5),
.Y(n_339)
);

OAI21x1_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_4),
.B(n_5),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_6),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_6),
.B(n_335),
.Y(n_342)
);


endmodule