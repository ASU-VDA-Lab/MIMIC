module real_jpeg_32142_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_0),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_0),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_0),
.A2(n_68),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

AOI22x1_ASAP7_75t_L g134 ( 
.A1(n_0),
.A2(n_68),
.B1(n_135),
.B2(n_139),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_0),
.A2(n_146),
.A3(n_151),
.B1(n_154),
.B2(n_162),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_0),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_0),
.B(n_132),
.Y(n_280)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_1),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_1),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g340 ( 
.A(n_1),
.Y(n_340)
);

CKINVDCx11_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_2),
.B(n_504),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_3),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_3),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_3),
.Y(n_480)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_6),
.A2(n_310),
.B1(n_313),
.B2(n_314),
.Y(n_309)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_6),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_6),
.A2(n_313),
.B1(n_382),
.B2(n_384),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_6),
.A2(n_313),
.B1(n_428),
.B2(n_433),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_6),
.A2(n_313),
.B1(n_471),
.B2(n_476),
.Y(n_470)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_7),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_8),
.A2(n_15),
.B(n_18),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

OAI22x1_ASAP7_75t_SL g29 ( 
.A1(n_10),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_34),
.B1(n_87),
.B2(n_91),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_34),
.B1(n_125),
.B2(n_128),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_10),
.A2(n_34),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_11),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_12),
.A2(n_343),
.B1(n_344),
.B2(n_346),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_12),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_12),
.A2(n_343),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_12),
.A2(n_343),
.B1(n_458),
.B2(n_461),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_12),
.A2(n_343),
.B1(n_486),
.B2(n_489),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_500),
.B(n_503),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_414),
.B(n_494),
.Y(n_19)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_358),
.B(n_411),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_297),
.Y(n_21)
);

OAI21x1_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_241),
.B(n_296),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_171),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_24),
.B(n_171),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_105),
.C(n_143),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_25),
.B(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_70),
.B2(n_71),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_26),
.B(n_72),
.C(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_26),
.B(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_26),
.B(n_354),
.C(n_355),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_26),
.B(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g401 ( 
.A(n_27),
.B(n_402),
.Y(n_401)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_38),
.B1(n_54),
.B2(n_64),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22x1_ASAP7_75t_L g238 ( 
.A1(n_29),
.A2(n_39),
.B1(n_65),
.B2(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_32),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_33),
.Y(n_432)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_37),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_38),
.A2(n_54),
.B(n_64),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_R g482 ( 
.A(n_38),
.B(n_425),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_39),
.B(n_65),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_39),
.A2(n_239),
.B1(n_427),
.B2(n_457),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_54),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_47),
.B2(n_50),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_48),
.Y(n_436)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_49),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_49),
.Y(n_197)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_53),
.Y(n_161)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_54),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_54),
.B(n_68),
.Y(n_266)
);

HB1xp67_ASAP7_75t_SL g425 ( 
.A(n_54),
.Y(n_425)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_57),
.Y(n_167)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_68),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_68),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_68),
.A2(n_198),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_68),
.B(n_248),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_68),
.A2(n_112),
.B(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_69),
.Y(n_463)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_81),
.B(n_104),
.Y(n_71)
);

OAI211xp5_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_82),
.B(n_85),
.C(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_73),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g223 ( 
.A(n_73),
.B(n_224),
.Y(n_223)
);

AO22x1_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_76),
.Y(n_227)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_81),
.B(n_274),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_95),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_83),
.Y(n_204)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_86),
.A2(n_96),
.B1(n_100),
.B2(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_90),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_90),
.Y(n_312)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_94),
.Y(n_259)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_94),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_95),
.A2(n_309),
.B(n_318),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_97),
.B(n_170),
.Y(n_169)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_105),
.A2(n_106),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_105),
.B(n_201),
.C(n_266),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_105),
.A2(n_143),
.B1(n_144),
.B2(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_105),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_105),
.B(n_336),
.Y(n_374)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_106),
.Y(n_294)
);

AOI22x1_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_123),
.B1(n_132),
.B2(n_133),
.Y(n_106)
);

AOI22x1_ASAP7_75t_L g261 ( 
.A1(n_107),
.A2(n_132),
.B1(n_133),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_107),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_107),
.A2(n_132),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_112),
.B(n_117),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_108),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_111),
.Y(n_383)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_111),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_112),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_114),
.Y(n_250)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_117),
.B(n_233),
.C(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_117),
.A2(n_236),
.B1(n_381),
.B2(n_388),
.Y(n_380)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_119),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_119),
.Y(n_347)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_124),
.Y(n_262)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_131),
.Y(n_387)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_134),
.Y(n_236)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_168),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_145),
.B(n_168),
.Y(n_287)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_169),
.B(n_342),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_170),
.A2(n_309),
.B1(n_337),
.B2(n_341),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_208),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_205),
.B2(n_206),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_173),
.B(n_208),
.C(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_201),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_175),
.Y(n_321)
);

AOI21x1_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_179),
.B(n_189),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_185),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_185),
.Y(n_488)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_198),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_224)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_201),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_201),
.B(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_202),
.B(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_202),
.B(n_280),
.Y(n_281)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_203),
.Y(n_318)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_206),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g268 ( 
.A(n_207),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_207),
.B(n_269),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_230),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_209),
.B(n_352),
.C(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_209),
.B(n_422),
.C(n_438),
.Y(n_450)
);

MAJx2_ASAP7_75t_L g493 ( 
.A(n_209),
.B(n_450),
.C(n_464),
.Y(n_493)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_210),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_211),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_211),
.A2(n_305),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

OA21x2_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B(n_219),
.Y(n_211)
);

OA22x2_ASAP7_75t_L g323 ( 
.A1(n_212),
.A2(n_213),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

NAND2x1p5_ASAP7_75t_L g399 ( 
.A(n_212),
.B(n_324),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_212),
.A2(n_219),
.B(n_470),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_212),
.A2(n_324),
.B1(n_470),
.B2(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_220),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_220),
.B(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_222),
.Y(n_489)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_223),
.Y(n_324)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_231),
.B(n_238),
.C(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_232),
.B(n_404),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_237),
.A2(n_238),
.B1(n_260),
.B2(n_271),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_237),
.B(n_260),
.C(n_287),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_237),
.A2(n_238),
.B1(n_323),
.B2(n_357),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g392 ( 
.A(n_238),
.B(n_356),
.C(n_393),
.Y(n_392)
);

AOI21x1_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_290),
.B(n_295),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_284),
.B(n_289),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_267),
.B(n_283),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_263),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_SL g283 ( 
.A(n_245),
.B(n_263),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_260),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_260),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_251),
.B(n_255),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_250),
.Y(n_405)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_260),
.A2(n_271),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_260),
.B(n_308),
.Y(n_352)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21x1_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_272),
.B(n_282),
.Y(n_267)
);

AOI21x1_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_279),
.B(n_281),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_326),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_299),
.B(n_301),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_319),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_304),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_330),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_330),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_319),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_332),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B(n_331),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_353),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_348),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_366),
.C(n_367),
.Y(n_365)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_348),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_353),
.Y(n_367)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_356),
.B(n_423),
.C(n_456),
.Y(n_483)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_357),
.B(n_455),
.Y(n_454)
);

NAND4xp25_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.C(n_364),
.D(n_390),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_368),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_373),
.C(n_376),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_376),
.B2(n_377),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_380),
.B2(n_389),
.Y(n_377)
);

OA21x2_ASAP7_75t_SL g441 ( 
.A1(n_378),
.A2(n_442),
.B(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_380),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_380),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_381),
.Y(n_403)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_412),
.B(n_413),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_409),
.B(n_410),
.Y(n_390)
);

NOR3xp33_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_409),
.C(n_410),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_394),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_392),
.B(n_400),
.C(n_446),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_400),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_396),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_399),
.B(n_502),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_407),
.Y(n_400)
);

HB1xp67_ASAP7_75t_SL g419 ( 
.A(n_401),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_402),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_465),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_444),
.B(n_447),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2x1p5_ASAP7_75t_L g497 ( 
.A(n_417),
.B(n_445),
.Y(n_497)
);

XOR2x2_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_441),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_420),
.B1(n_439),
.B2(n_440),
.Y(n_418)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_419),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_440),
.C(n_441),
.Y(n_448)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_423),
.B1(n_424),
.B2(n_438),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_424),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B(n_437),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_445),
.Y(n_444)
);

OAI21x1_ASAP7_75t_SL g496 ( 
.A1(n_447),
.A2(n_497),
.B(n_498),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_448),
.B(n_449),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_454),
.B2(n_464),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_454),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI221x1_ASAP7_75t_L g494 ( 
.A1(n_465),
.A2(n_467),
.B1(n_495),
.B2(n_496),
.C(n_499),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_490),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_468),
.B(n_484),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_468),
.B(n_484),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_481),
.C(n_483),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_481),
.Y(n_492)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx8_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx6_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_492),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_484),
.B(n_501),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_485),
.Y(n_502)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_493),
.Y(n_495)
);


endmodule