module real_jpeg_2198_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_288;
wire n_221;
wire n_292;
wire n_249;
wire n_215;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_195;
wire n_110;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_244;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_2),
.A2(n_27),
.B1(n_47),
.B2(n_48),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_2),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_2),
.A2(n_27),
.B1(n_58),
.B2(n_59),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_37),
.B1(n_58),
.B2(n_59),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_29),
.C(n_33),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_31),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_3),
.B(n_44),
.C(n_48),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_3),
.B(n_84),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_3),
.B(n_56),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_3),
.B(n_57),
.C(n_59),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_3),
.B(n_50),
.Y(n_227)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_40),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_6),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_6),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_106)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_9),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_15),
.B(n_291),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_11),
.B(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_52),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_12),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_286),
.B(n_289),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_73),
.B(n_285),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_70),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_18),
.B(n_70),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_64),
.C(n_66),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_19),
.B(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.C(n_53),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_20),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_20),
.A2(n_99),
.B1(n_137),
.B2(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_20),
.B(n_137),
.C(n_147),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_20),
.A2(n_99),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_22),
.A2(n_67),
.B(n_69),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_24),
.B(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_33),
.B(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_36),
.B(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_38),
.A2(n_53),
.B1(n_257),
.B2(n_274),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_38),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_38)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_39),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_41),
.A2(n_50),
.B1(n_95),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_42),
.A2(n_46),
.B(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

AOI22x1_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_46),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_48),
.B1(n_57),
.B2(n_60),
.Y(n_62)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_48),
.B(n_220),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_53),
.A2(n_257),
.B1(n_258),
.B2(n_261),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_53),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_53),
.B(n_121),
.C(n_258),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_61),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_61),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_55),
.A2(n_106),
.B(n_107),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_55),
.A2(n_61),
.B1(n_90),
.B2(n_91),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_55),
.A2(n_61),
.B(n_91),
.Y(n_163)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_56),
.A2(n_63),
.B1(n_109),
.B2(n_136),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_59),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_64),
.B(n_66),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_67),
.B(n_71),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_70),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_70),
.B(n_287),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_72),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_280),
.B(n_284),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_251),
.B(n_277),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_141),
.B(n_250),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_122),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_77),
.B(n_122),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_100),
.C(n_111),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_78),
.B(n_100),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_92),
.B2(n_93),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_94),
.C(n_99),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_88),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_81),
.A2(n_88),
.B1(n_89),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_81),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_83),
.A2(n_84),
.B1(n_116),
.B2(n_153),
.Y(n_152)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_86),
.B(n_115),
.Y(n_114)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_86),
.A2(n_115),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_88),
.A2(n_89),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_88),
.A2(n_89),
.B1(n_200),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_89),
.B(n_195),
.C(n_200),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_89),
.B(n_152),
.C(n_227),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_120),
.C(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_94),
.A2(n_98),
.B1(n_163),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_94),
.A2(n_98),
.B1(n_117),
.B2(n_118),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_94),
.B(n_117),
.C(n_234),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_96),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_110),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_105),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_110),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_103),
.B(n_116),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_110),
.A2(n_126),
.B(n_132),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_111),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_119),
.C(n_120),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_112),
.A2(n_113),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_114),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_117),
.A2(n_118),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_117),
.B(n_221),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_121),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_120),
.A2(n_121),
.B1(n_256),
.B2(n_262),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_120),
.A2(n_121),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_121),
.B(n_271),
.C(n_275),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_140),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_133),
.B2(n_134),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_125),
.B(n_133),
.C(n_140),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_130),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_131),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_137),
.B(n_139),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_171),
.C(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_137),
.A2(n_155),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_139),
.A2(n_255),
.B1(n_263),
.B2(n_264),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_139),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_245),
.B(n_249),
.Y(n_141)
);

OAI211xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_174),
.B(n_188),
.C(n_244),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_164),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_164),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_156),
.B2(n_157),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_159),
.C(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_151),
.A2(n_152),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_152),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_152),
.B(n_215),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_170),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_172),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_189),
.C(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_176),
.B(n_177),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_178),
.B(n_180),
.C(n_186),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_185),
.B2(n_186),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_206),
.B(n_243),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_194),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_237),
.B(n_242),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_231),
.B(n_236),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_223),
.B(n_230),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_217),
.B(n_222),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_214),
.B(n_216),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_229),
.Y(n_230)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_241),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_267),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_266),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_266),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_256),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_258),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_264),
.C(n_265),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_276),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_276),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_283),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);


endmodule