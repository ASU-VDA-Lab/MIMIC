module fake_netlist_1_11120_n_639 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_639);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_639;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_72), .Y(n_75) );
INVxp33_ASAP7_75t_L g76 ( .A(n_69), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_44), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_19), .Y(n_78) );
INVxp67_ASAP7_75t_L g79 ( .A(n_26), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_11), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_4), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_29), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_49), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_55), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_13), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_25), .Y(n_86) );
BUFx2_ASAP7_75t_L g87 ( .A(n_57), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_10), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_39), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_21), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_23), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_35), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_53), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_12), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_2), .Y(n_96) );
INVxp33_ASAP7_75t_SL g97 ( .A(n_3), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_0), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_17), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_52), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_40), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_22), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_58), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_5), .Y(n_104) );
INVxp33_ASAP7_75t_L g105 ( .A(n_74), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_0), .Y(n_106) );
NOR2xp67_ASAP7_75t_L g107 ( .A(n_13), .B(n_38), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_37), .Y(n_108) );
NOR2xp67_ASAP7_75t_L g109 ( .A(n_32), .B(n_59), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_54), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_6), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_7), .Y(n_112) );
BUFx10_ASAP7_75t_L g113 ( .A(n_10), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_56), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_60), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_64), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_19), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_27), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_41), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_68), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_103), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_103), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_103), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_112), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_112), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_112), .Y(n_126) );
AND2x6_ASAP7_75t_L g127 ( .A(n_83), .B(n_33), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_119), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_87), .B(n_1), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_112), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_103), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_103), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_75), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_75), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_87), .B(n_1), .Y(n_136) );
AND3x2_ASAP7_75t_L g137 ( .A(n_95), .B(n_2), .C(n_3), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_103), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_77), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_77), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_94), .B(n_4), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_104), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_98), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_82), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_82), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_86), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_91), .B(n_5), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_92), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_113), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_99), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_93), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_101), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_113), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_156), .B(n_76), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_159), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_132), .Y(n_163) );
NAND3xp33_ASAP7_75t_L g164 ( .A(n_130), .B(n_117), .C(n_80), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_143), .B(n_113), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_156), .B(n_105), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_157), .B(n_106), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_156), .B(n_78), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_157), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_159), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_159), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_160), .B(n_84), .Y(n_173) );
AND2x6_ASAP7_75t_L g174 ( .A(n_136), .B(n_114), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_132), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_156), .B(n_79), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_136), .A2(n_78), .B1(n_80), .B2(n_81), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_126), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_160), .B(n_97), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_160), .B(n_85), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_126), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_160), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_126), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_144), .B(n_120), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_126), .Y(n_186) );
AO22x2_ASAP7_75t_L g187 ( .A1(n_134), .A2(n_120), .B1(n_118), .B2(n_115), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_142), .A2(n_81), .B1(n_111), .B2(n_88), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_124), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_128), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_134), .B(n_118), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_124), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_128), .Y(n_194) );
NAND2xp33_ASAP7_75t_L g195 ( .A(n_127), .B(n_108), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_121), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_128), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_125), .Y(n_198) );
CKINVDCx8_ASAP7_75t_R g199 ( .A(n_127), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_125), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_135), .B(n_111), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_151), .A2(n_96), .B1(n_116), .B2(n_107), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_131), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_131), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_135), .B(n_140), .Y(n_206) );
BUFx4_ASAP7_75t_L g207 ( .A(n_137), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_158), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_140), .B(n_113), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_147), .A2(n_90), .B1(n_100), .B2(n_110), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_158), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_127), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_132), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_147), .B(n_115), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_139), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_149), .B(n_114), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_121), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_209), .B(n_149), .Y(n_218) );
NOR2xp33_ASAP7_75t_SL g219 ( .A(n_199), .B(n_127), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_211), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_212), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_170), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_211), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_200), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_183), .B(n_150), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_200), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_183), .B(n_150), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_166), .B(n_153), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_200), .Y(n_229) );
OR2x6_ASAP7_75t_L g230 ( .A(n_187), .B(n_153), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_168), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_203), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_164), .B(n_155), .Y(n_233) );
INVx5_ASAP7_75t_L g234 ( .A(n_174), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_174), .A2(n_127), .B1(n_154), .B2(n_152), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_203), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_203), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_178), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_174), .A2(n_127), .B1(n_154), .B2(n_152), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_168), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_169), .B(n_155), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_212), .B(n_148), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
AND2x2_ASAP7_75t_SL g244 ( .A(n_195), .B(n_101), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_182), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_182), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_166), .B(n_146), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_210), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_199), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_194), .Y(n_251) );
BUFx12f_ASAP7_75t_L g252 ( .A(n_174), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_182), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_169), .B(n_148), .Y(n_254) );
INVx4_ASAP7_75t_L g255 ( .A(n_174), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_201), .B(n_146), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_174), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_184), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_169), .B(n_145), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_195), .A2(n_145), .B(n_141), .Y(n_260) );
INVxp67_ASAP7_75t_SL g261 ( .A(n_214), .Y(n_261) );
CKINVDCx6p67_ASAP7_75t_R g262 ( .A(n_161), .Y(n_262) );
INVx5_ASAP7_75t_L g263 ( .A(n_184), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_184), .Y(n_264) );
BUFx8_ASAP7_75t_L g265 ( .A(n_207), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_190), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_190), .Y(n_267) );
NAND2x2_ASAP7_75t_L g268 ( .A(n_207), .B(n_6), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_194), .Y(n_269) );
NOR2x1_ASAP7_75t_R g270 ( .A(n_167), .B(n_141), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_180), .B(n_102), .Y(n_271) );
OR2x6_ASAP7_75t_L g272 ( .A(n_187), .B(n_129), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_198), .Y(n_273) );
INVx4_ASAP7_75t_L g274 ( .A(n_214), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_191), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_187), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g277 ( .A1(n_189), .A2(n_129), .B1(n_139), .B2(n_102), .C(n_108), .Y(n_277) );
NOR2x1_ASAP7_75t_SL g278 ( .A(n_230), .B(n_198), .Y(n_278) );
INVxp33_ASAP7_75t_L g279 ( .A(n_222), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_224), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_261), .B(n_181), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_276), .A2(n_187), .B1(n_214), .B2(n_201), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_222), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_255), .B(n_201), .Y(n_284) );
CKINVDCx16_ASAP7_75t_R g285 ( .A(n_231), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_240), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_240), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_224), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_219), .A2(n_173), .B(n_191), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_255), .B(n_177), .Y(n_291) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_260), .A2(n_110), .B(n_216), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_266), .Y(n_293) );
AOI221x1_ASAP7_75t_L g294 ( .A1(n_267), .A2(n_133), .B1(n_132), .B2(n_138), .C(n_123), .Y(n_294) );
BUFx4f_ASAP7_75t_L g295 ( .A(n_252), .Y(n_295) );
INVx6_ASAP7_75t_SL g296 ( .A(n_230), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_248), .Y(n_297) );
NOR2x1_ASAP7_75t_R g298 ( .A(n_265), .B(n_215), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_265), .Y(n_299) );
AOI21xp33_ASAP7_75t_L g300 ( .A1(n_270), .A2(n_202), .B(n_185), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_267), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_228), .B(n_206), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_273), .Y(n_303) );
OR2x6_ASAP7_75t_L g304 ( .A(n_252), .B(n_186), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_265), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_273), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_228), .B(n_215), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_276), .A2(n_193), .B1(n_204), .B2(n_176), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_250), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_230), .Y(n_310) );
NOR2xp67_ASAP7_75t_SL g311 ( .A(n_250), .B(n_127), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g312 ( .A1(n_226), .A2(n_192), .B(n_197), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_230), .A2(n_208), .B1(n_205), .B2(n_139), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_255), .Y(n_314) );
OR2x6_ASAP7_75t_L g315 ( .A(n_257), .B(n_109), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_234), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_257), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_272), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_248), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_226), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_272), .B(n_7), .Y(n_321) );
INVx1_ASAP7_75t_SL g322 ( .A(n_256), .Y(n_322) );
INVx5_ASAP7_75t_L g323 ( .A(n_257), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_297), .B(n_256), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_286), .A2(n_287), .B1(n_283), .B2(n_318), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_307), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_290), .A2(n_294), .B(n_293), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_307), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_282), .A2(n_272), .B1(n_244), .B2(n_274), .Y(n_329) );
CKINVDCx11_ASAP7_75t_R g330 ( .A(n_285), .Y(n_330) );
CKINVDCx14_ASAP7_75t_R g331 ( .A(n_299), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_318), .A2(n_272), .B1(n_244), .B2(n_274), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_319), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_296), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_323), .B(n_234), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_310), .A2(n_249), .B1(n_274), .B2(n_277), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_302), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_309), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_296), .A2(n_234), .B1(n_259), .B2(n_239), .Y(n_340) );
NAND2xp33_ASAP7_75t_L g341 ( .A(n_309), .B(n_250), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_310), .A2(n_234), .B1(n_259), .B2(n_235), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_288), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_301), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_279), .B(n_259), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_322), .B(n_218), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_284), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_313), .A2(n_234), .B1(n_225), .B2(n_227), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_288), .Y(n_349) );
CKINVDCx6p67_ASAP7_75t_R g350 ( .A(n_304), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_293), .A2(n_303), .B(n_306), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_321), .A2(n_268), .B1(n_254), .B2(n_241), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_352), .A2(n_300), .B1(n_249), .B2(n_271), .C(n_233), .Y(n_353) );
BUFx12f_ASAP7_75t_L g354 ( .A(n_330), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g355 ( .A1(n_332), .A2(n_321), .B1(n_268), .B2(n_278), .Y(n_355) );
OAI31xp33_ASAP7_75t_SL g356 ( .A1(n_352), .A2(n_291), .A3(n_312), .B(n_284), .Y(n_356) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_338), .A2(n_281), .B(n_315), .C(n_291), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_326), .A2(n_291), .B1(n_306), .B2(n_303), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_329), .A2(n_284), .B1(n_308), .B2(n_299), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_334), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_328), .A2(n_349), .B1(n_343), .B2(n_345), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_324), .A2(n_233), .B1(n_301), .B2(n_315), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_351), .A2(n_292), .B(n_278), .Y(n_363) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_337), .A2(n_305), .B1(n_315), .B2(n_304), .C(n_295), .Y(n_364) );
NAND3xp33_ASAP7_75t_L g365 ( .A(n_325), .B(n_315), .C(n_233), .Y(n_365) );
NAND3xp33_ASAP7_75t_L g366 ( .A(n_346), .B(n_294), .C(n_220), .Y(n_366) );
INVx4_ASAP7_75t_L g367 ( .A(n_350), .Y(n_367) );
AOI322xp5_ASAP7_75t_L g368 ( .A1(n_331), .A2(n_305), .A3(n_298), .B1(n_223), .B2(n_220), .C1(n_14), .C2(n_15), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_344), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g370 ( .A1(n_347), .A2(n_304), .B1(n_295), .B2(n_243), .C(n_245), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_344), .B(n_262), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_331), .A2(n_223), .B1(n_320), .B2(n_253), .C(n_232), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_350), .A2(n_292), .B1(n_320), .B2(n_304), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_327), .A2(n_292), .B(n_280), .Y(n_375) );
OAI22xp5_ASAP7_75t_SL g376 ( .A1(n_330), .A2(n_317), .B1(n_323), .B2(n_262), .Y(n_376) );
OAI21x1_ASAP7_75t_L g377 ( .A1(n_327), .A2(n_280), .B(n_289), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_353), .A2(n_348), .B1(n_342), .B2(n_340), .C(n_333), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_375), .A2(n_121), .B(n_122), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_369), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_377), .Y(n_382) );
OAI21xp5_ASAP7_75t_SL g383 ( .A1(n_355), .A2(n_336), .B(n_314), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_368), .A2(n_295), .B1(n_253), .B2(n_245), .C(n_238), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_360), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_358), .B(n_361), .Y(n_386) );
OA222x2_ASAP7_75t_L g387 ( .A1(n_356), .A2(n_314), .B1(n_316), .B2(n_341), .C1(n_238), .C2(n_264), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_364), .B(n_263), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_358), .B(n_289), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_359), .A2(n_317), .B1(n_323), .B2(n_309), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_362), .A2(n_317), .B1(n_323), .B2(n_309), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_361), .Y(n_392) );
OAI33xp33_ASAP7_75t_L g393 ( .A1(n_372), .A2(n_188), .A3(n_162), .B1(n_138), .B2(n_122), .B3(n_123), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_367), .A2(n_323), .B1(n_314), .B2(n_309), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_374), .B(n_133), .C(n_132), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_365), .A2(n_336), .B1(n_269), .B2(n_311), .Y(n_396) );
AOI322xp5_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_8), .A3(n_9), .B1(n_11), .B2(n_12), .C1(n_14), .C2(n_15), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_362), .B(n_339), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_373), .A2(n_336), .B1(n_269), .B2(n_311), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_366), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_357), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_367), .A2(n_341), .B1(n_339), .B2(n_316), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_371), .B(n_263), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_363), .A2(n_232), .B(n_229), .Y(n_404) );
OAI33xp33_ASAP7_75t_L g405 ( .A1(n_378), .A2(n_188), .A3(n_162), .B1(n_138), .B2(n_123), .B3(n_122), .Y(n_405) );
OAI31xp33_ASAP7_75t_L g406 ( .A1(n_370), .A2(n_229), .A3(n_236), .B(n_237), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_374), .B(n_339), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_354), .B(n_263), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_376), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_353), .A2(n_264), .B1(n_238), .B2(n_245), .C(n_237), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g411 ( .A(n_368), .B(n_172), .C(n_179), .D(n_171), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_355), .A2(n_264), .B1(n_275), .B2(n_251), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_407), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_381), .Y(n_414) );
AOI211xp5_ASAP7_75t_L g415 ( .A1(n_409), .A2(n_133), .B(n_132), .C(n_236), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_382), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_407), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_386), .B(n_339), .Y(n_418) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_380), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_401), .A2(n_251), .B(n_133), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_382), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_392), .B(n_8), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_380), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_398), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_392), .B(n_9), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_386), .B(n_16), .Y(n_427) );
OAI31xp33_ASAP7_75t_L g428 ( .A1(n_383), .A2(n_409), .A3(n_411), .B(n_384), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_385), .B(n_16), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_385), .B(n_17), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_380), .Y(n_431) );
AOI33xp33_ASAP7_75t_L g432 ( .A1(n_401), .A2(n_165), .A3(n_171), .B1(n_172), .B2(n_179), .B3(n_217), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_398), .B(n_133), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_389), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_379), .A2(n_258), .B1(n_246), .B2(n_247), .C(n_263), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_389), .B(n_18), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_400), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_400), .B(n_258), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_404), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_388), .B(n_247), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_387), .B(n_133), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_410), .A2(n_246), .B1(n_275), .B2(n_251), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_395), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_395), .B(n_18), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_387), .B(n_24), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_412), .B(n_251), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_397), .B(n_28), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_403), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_397), .B(n_30), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_405), .A2(n_250), .B(n_251), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_402), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_390), .B(n_263), .Y(n_453) );
NOR2xp67_ASAP7_75t_L g454 ( .A(n_391), .B(n_31), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_394), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_396), .Y(n_456) );
AND2x2_ASAP7_75t_SL g457 ( .A(n_399), .B(n_250), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_393), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_408), .Y(n_459) );
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_406), .A2(n_165), .B1(n_242), .B2(n_217), .C(n_196), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_437), .B(n_196), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_435), .B(n_34), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_437), .B(n_36), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_425), .B(n_42), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_421), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_427), .B(n_43), .Y(n_467) );
AND3x1_ASAP7_75t_L g468 ( .A(n_448), .B(n_45), .C(n_46), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_425), .B(n_47), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_438), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_425), .B(n_48), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_459), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_414), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g474 ( .A(n_428), .B(n_448), .C(n_450), .D(n_427), .Y(n_474) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_419), .A2(n_213), .B(n_175), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_435), .B(n_50), .Y(n_476) );
INVx2_ASAP7_75t_SL g477 ( .A(n_414), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_438), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_413), .B(n_51), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_413), .B(n_61), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_418), .B(n_62), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_414), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_417), .B(n_63), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_418), .B(n_65), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_417), .B(n_66), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_416), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_418), .B(n_67), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_434), .B(n_70), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_429), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_430), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
OAI211xp5_ASAP7_75t_L g492 ( .A1(n_428), .A2(n_163), .B(n_175), .C(n_213), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_416), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_434), .B(n_71), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_430), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_423), .B(n_426), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_440), .B(n_73), .Y(n_497) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_445), .B(n_163), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_415), .A2(n_221), .B(n_175), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_459), .B(n_163), .C(n_175), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_450), .A2(n_163), .B1(n_175), .B2(n_213), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_423), .B(n_163), .Y(n_502) );
NAND5xp2_ASAP7_75t_SL g503 ( .A(n_446), .B(n_213), .C(n_221), .D(n_442), .E(n_457), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_449), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_449), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_434), .B(n_213), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_434), .B(n_221), .Y(n_507) );
AOI22x1_ASAP7_75t_L g508 ( .A1(n_446), .A2(n_221), .B1(n_452), .B2(n_442), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_422), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_449), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_442), .B(n_440), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_439), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_419), .B(n_433), .Y(n_513) );
NOR2xp67_ASAP7_75t_L g514 ( .A(n_492), .B(n_452), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_474), .B(n_452), .C(n_441), .D(n_415), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_511), .B(n_424), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_472), .B(n_452), .C(n_456), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_505), .B(n_422), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_513), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_461), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_511), .B(n_424), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_466), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_513), .B(n_424), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_508), .B(n_454), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_488), .B(n_454), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_482), .B(n_431), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_470), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_510), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_470), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_478), .Y(n_530) );
OAI21xp33_ASAP7_75t_L g531 ( .A1(n_501), .A2(n_457), .B(n_441), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_482), .B(n_431), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_478), .Y(n_533) );
INVxp67_ASAP7_75t_L g534 ( .A(n_504), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_489), .B(n_458), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_477), .B(n_422), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_490), .B(n_458), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_494), .Y(n_538) );
AOI211xp5_ASAP7_75t_SL g539 ( .A1(n_483), .A2(n_436), .B(n_455), .C(n_420), .Y(n_539) );
OAI211xp5_ASAP7_75t_SL g540 ( .A1(n_467), .A2(n_464), .B(n_495), .C(n_498), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_496), .B(n_444), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_512), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_473), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_477), .B(n_479), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_479), .B(n_444), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_463), .B(n_431), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_468), .A2(n_436), .B(n_457), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_486), .B(n_433), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_463), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_476), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_480), .B(n_455), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_486), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_491), .B(n_433), .Y(n_553) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_462), .B(n_460), .C(n_453), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_491), .B(n_420), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_493), .B(n_439), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_476), .B(n_453), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_480), .B(n_432), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_483), .B(n_443), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_493), .B(n_447), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_520), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_522), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_527), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_528), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_529), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_530), .Y(n_566) );
OAI21xp5_ASAP7_75t_SL g567 ( .A1(n_515), .A2(n_494), .B(n_488), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_559), .A2(n_487), .B1(n_484), .B2(n_481), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_541), .B(n_509), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_547), .A2(n_503), .B(n_485), .C(n_497), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_533), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_534), .B(n_484), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_517), .A2(n_508), .B1(n_485), .B2(n_500), .C(n_497), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_538), .A2(n_487), .B1(n_488), .B2(n_465), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_518), .Y(n_575) );
NAND2xp33_ASAP7_75t_L g576 ( .A(n_525), .B(n_471), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_543), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_523), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_542), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g580 ( .A1(n_514), .A2(n_465), .B1(n_469), .B2(n_499), .C(n_502), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_518), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_544), .B(n_469), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_537), .B(n_506), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_539), .A2(n_443), .B(n_451), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_535), .B(n_475), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_554), .A2(n_503), .B1(n_506), .B2(n_460), .C(n_451), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_558), .B(n_507), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_516), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g589 ( .A1(n_531), .A2(n_447), .B1(n_475), .B2(n_507), .C(n_525), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_523), .B(n_549), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_521), .B(n_536), .Y(n_591) );
BUFx3_ASAP7_75t_L g592 ( .A(n_536), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_521), .Y(n_593) );
INVx2_ASAP7_75t_SL g594 ( .A(n_526), .Y(n_594) );
O2A1O1Ixp5_ASAP7_75t_L g595 ( .A1(n_524), .A2(n_545), .B(n_559), .C(n_550), .Y(n_595) );
BUFx2_ASAP7_75t_L g596 ( .A(n_548), .Y(n_596) );
NAND2x1_ASAP7_75t_L g597 ( .A(n_526), .B(n_532), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_532), .B(n_556), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_540), .A2(n_524), .B(n_551), .Y(n_599) );
AO22x1_ASAP7_75t_L g600 ( .A1(n_553), .A2(n_552), .B1(n_555), .B2(n_557), .Y(n_600) );
AO22x2_ASAP7_75t_SL g601 ( .A1(n_553), .A2(n_555), .B1(n_546), .B2(n_560), .Y(n_601) );
XNOR2x1_ASAP7_75t_L g602 ( .A(n_560), .B(n_468), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_519), .B(n_541), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_520), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_528), .Y(n_605) );
XNOR2x2_ASAP7_75t_L g606 ( .A(n_517), .B(n_474), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_520), .Y(n_607) );
AOI211xp5_ASAP7_75t_L g608 ( .A1(n_567), .A2(n_599), .B(n_589), .C(n_600), .Y(n_608) );
OAI31xp33_ASAP7_75t_L g609 ( .A1(n_605), .A2(n_602), .A3(n_606), .B(n_574), .Y(n_609) );
XNOR2x1_ASAP7_75t_L g610 ( .A(n_606), .B(n_602), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_603), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_564), .B(n_579), .Y(n_612) );
A2O1A1Ixp33_ASAP7_75t_L g613 ( .A1(n_570), .A2(n_595), .B(n_597), .C(n_576), .Y(n_613) );
INVxp33_ASAP7_75t_SL g614 ( .A(n_574), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_603), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_587), .A2(n_583), .B1(n_572), .B2(n_582), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_592), .B(n_596), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_561), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_607), .Y(n_619) );
AO21x1_ASAP7_75t_L g620 ( .A1(n_562), .A2(n_604), .B(n_584), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_617), .Y(n_621) );
AO22x2_ASAP7_75t_L g622 ( .A1(n_610), .A2(n_577), .B1(n_592), .B2(n_591), .Y(n_622) );
NAND4xp75_ASAP7_75t_L g623 ( .A(n_609), .B(n_584), .C(n_586), .D(n_568), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_618), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_614), .A2(n_594), .B1(n_563), .B2(n_565), .C(n_566), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_613), .A2(n_594), .B1(n_571), .B2(n_590), .C(n_578), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_619), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_626), .A2(n_620), .B1(n_615), .B2(n_611), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_623), .A2(n_613), .B1(n_608), .B2(n_616), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_625), .A2(n_612), .B(n_580), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_622), .A2(n_612), .B1(n_573), .B2(n_569), .C(n_575), .Y(n_631) );
NOR3x1_ASAP7_75t_L g632 ( .A(n_629), .B(n_622), .C(n_624), .Y(n_632) );
OR4x2_ASAP7_75t_L g633 ( .A(n_630), .B(n_601), .C(n_621), .D(n_627), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_632), .A2(n_628), .B(n_631), .Y(n_634) );
AOI22x1_ASAP7_75t_L g635 ( .A1(n_633), .A2(n_591), .B1(n_581), .B2(n_588), .Y(n_635) );
INVx2_ASAP7_75t_SL g636 ( .A(n_635), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_636), .A2(n_634), .B1(n_593), .B2(n_598), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_637), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_638), .A2(n_601), .B(n_585), .Y(n_639) );
endmodule