module fake_jpeg_26798_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_42),
.Y(n_60)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_58),
.Y(n_70)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_59),
.Y(n_72)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_16),
.B1(n_42),
.B2(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_41),
.B1(n_24),
.B2(n_25),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_16),
.B1(n_19),
.B2(n_30),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_86),
.B1(n_61),
.B2(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_79),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_41),
.B1(n_39),
.B2(n_42),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_51),
.B1(n_50),
.B2(n_45),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_40),
.C(n_37),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_40),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_37),
.B(n_25),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_26),
.B(n_27),
.C(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_30),
.B(n_43),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_21),
.B(n_33),
.Y(n_95)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_43),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_95),
.B1(n_62),
.B2(n_59),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_93),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_69),
.B(n_68),
.Y(n_91)
);

BUFx12f_ASAP7_75t_SL g118 ( 
.A(n_91),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_46),
.C(n_56),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_33),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_108),
.Y(n_129)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_20),
.C(n_23),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_21),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_64),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_112),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_64),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_36),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_115),
.B(n_84),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_16),
.B1(n_41),
.B2(n_61),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_65),
.B1(n_62),
.B2(n_46),
.Y(n_132)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_122),
.Y(n_147)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_120),
.A2(n_80),
.B1(n_81),
.B2(n_22),
.Y(n_177)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_127),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_126),
.B(n_55),
.Y(n_166)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_130),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_30),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_132),
.B1(n_86),
.B2(n_111),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_33),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_139),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_62),
.B1(n_16),
.B2(n_65),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_135),
.A2(n_89),
.B1(n_108),
.B2(n_102),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_136),
.A2(n_17),
.B1(n_88),
.B2(n_80),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_32),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_32),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_32),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

CKINVDCx12_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_144),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_137),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_161),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_94),
.B1(n_104),
.B2(n_102),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_94),
.B1(n_110),
.B2(n_92),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_153),
.B(n_162),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_21),
.A3(n_112),
.B1(n_114),
.B2(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_92),
.B1(n_111),
.B2(n_103),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_169),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_136),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_29),
.A3(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_106),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_122),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_174),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_27),
.B(n_29),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_172),
.B(n_22),
.C(n_31),
.Y(n_208)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_26),
.B(n_55),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_125),
.B1(n_134),
.B2(n_124),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_177),
.B1(n_127),
.B2(n_164),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_130),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_181),
.B(n_10),
.Y(n_232)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_193),
.Y(n_219)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_190),
.B1(n_31),
.B2(n_23),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_136),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_189),
.C(n_191),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_141),
.C(n_140),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_119),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_133),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_119),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_202),
.B(n_208),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_20),
.C(n_120),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_204),
.C(n_207),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_155),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_205),
.Y(n_225)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_152),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_147),
.A2(n_120),
.B(n_28),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_147),
.B(n_20),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_138),
.C(n_121),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_209),
.B(n_215),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_170),
.B1(n_148),
.B2(n_154),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_210),
.A2(n_230),
.B1(n_23),
.B2(n_18),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_172),
.B(n_157),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_157),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_182),
.A2(n_146),
.B1(n_156),
.B2(n_172),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_220),
.B1(n_229),
.B2(n_198),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_180),
.A2(n_158),
.B1(n_167),
.B2(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_226),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_171),
.B(n_162),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_28),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_227),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_138),
.Y(n_224)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_152),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_180),
.A2(n_31),
.B1(n_18),
.B2(n_17),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_178),
.A2(n_31),
.B1(n_17),
.B2(n_18),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_186),
.B1(n_197),
.B2(n_189),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_232),
.B(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_234),
.Y(n_248)
);

NOR2x1_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_20),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_179),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_250),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_237),
.B(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_193),
.B1(n_196),
.B2(n_204),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_188),
.B1(n_183),
.B2(n_18),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_18),
.B1(n_20),
.B2(n_2),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_249),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_210),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_216),
.C(n_211),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_253),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_236),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_10),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_218),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_228),
.B(n_230),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_259),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_216),
.C(n_211),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_261),
.C(n_264),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_217),
.B(n_213),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_212),
.C(n_233),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_228),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_263),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_212),
.C(n_221),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_254),
.B1(n_240),
.B2(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_213),
.C(n_223),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_270),
.C(n_272),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_224),
.C(n_209),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_229),
.C(n_234),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_280),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_246),
.B(n_245),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_279),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_240),
.B(n_248),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_278),
.A2(n_267),
.B(n_12),
.Y(n_292)
);

FAx1_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_252),
.CI(n_244),
.CON(n_279),
.SN(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_270),
.B(n_256),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_249),
.B1(n_3),
.B2(n_4),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_284),
.A2(n_268),
.B1(n_258),
.B2(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_7),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_287),
.Y(n_289)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_274),
.B1(n_279),
.B2(n_286),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_267),
.B(n_11),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_297),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_278),
.B(n_279),
.Y(n_305)
);

OAI321xp33_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_9),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C(n_7),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_298),
.B(n_13),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_28),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_23),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_287),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_7),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_9),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_284),
.Y(n_302)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_304),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_293),
.B(n_286),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_295),
.B(n_292),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_295),
.C(n_288),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_308),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_317),
.C(n_314),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_288),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_311),
.C(n_318),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_310),
.B(n_312),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_9),
.A3(n_23),
.B1(n_5),
.B2(n_6),
.C1(n_1),
.C2(n_4),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_5),
.B(n_6),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_5),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_6),
.B(n_23),
.Y(n_325)
);


endmodule