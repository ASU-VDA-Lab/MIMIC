module real_aes_2272_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_787, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_787;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g174 ( .A(n_0), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_1), .B(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_2), .B(n_180), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_3), .B(n_177), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_4), .A2(n_44), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_4), .Y(n_450) );
INVx1_ASAP7_75t_L g140 ( .A(n_5), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_6), .B(n_180), .Y(n_202) );
NAND2xp33_ASAP7_75t_SL g160 ( .A(n_7), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g131 ( .A(n_8), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_9), .Y(n_117) );
AND2x2_ASAP7_75t_L g200 ( .A(n_10), .B(n_183), .Y(n_200) );
AND2x2_ASAP7_75t_L g501 ( .A(n_11), .B(n_156), .Y(n_501) );
AND2x2_ASAP7_75t_L g552 ( .A(n_12), .B(n_211), .Y(n_552) );
INVx2_ASAP7_75t_L g134 ( .A(n_13), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_14), .B(n_177), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_15), .Y(n_110) );
AOI221x1_ASAP7_75t_L g152 ( .A1(n_16), .A2(n_153), .B1(n_155), .B2(n_156), .C(n_159), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_17), .B(n_180), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_18), .B(n_180), .Y(n_557) );
INVx1_ASAP7_75t_L g113 ( .A(n_19), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_20), .A2(n_92), .B1(n_135), .B2(n_180), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_21), .A2(n_155), .B(n_204), .Y(n_203) );
AOI221xp5_ASAP7_75t_SL g247 ( .A1(n_22), .A2(n_36), .B1(n_155), .B2(n_180), .C(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_23), .B(n_175), .Y(n_205) );
OR2x2_ASAP7_75t_L g133 ( .A(n_24), .B(n_91), .Y(n_133) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_24), .A2(n_91), .B(n_134), .Y(n_158) );
INVxp67_ASAP7_75t_L g151 ( .A(n_25), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_26), .B(n_177), .Y(n_242) );
AND2x2_ASAP7_75t_L g194 ( .A(n_27), .B(n_182), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_28), .A2(n_155), .B(n_173), .Y(n_172) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_29), .A2(n_156), .B(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_30), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_31), .B(n_177), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_32), .A2(n_155), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_33), .B(n_177), .Y(n_533) );
AND2x2_ASAP7_75t_L g142 ( .A(n_34), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g146 ( .A(n_34), .Y(n_146) );
AND2x2_ASAP7_75t_L g161 ( .A(n_34), .B(n_140), .Y(n_161) );
OR2x6_ASAP7_75t_L g111 ( .A(n_35), .B(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_37), .B(n_180), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_38), .A2(n_84), .B1(n_144), .B2(n_155), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_39), .B(n_177), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_40), .A2(n_49), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_40), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_41), .B(n_180), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_42), .B(n_175), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_43), .A2(n_155), .B(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_44), .Y(n_451) );
AND2x2_ASAP7_75t_L g181 ( .A(n_45), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_46), .B(n_175), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_47), .B(n_182), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_48), .B(n_180), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_49), .Y(n_777) );
INVx1_ASAP7_75t_L g138 ( .A(n_50), .Y(n_138) );
INVx1_ASAP7_75t_L g165 ( .A(n_50), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_51), .B(n_177), .Y(n_499) );
AND2x2_ASAP7_75t_L g511 ( .A(n_52), .B(n_182), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_53), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_54), .B(n_180), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_55), .B(n_175), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_56), .B(n_175), .Y(n_532) );
AND2x2_ASAP7_75t_L g223 ( .A(n_57), .B(n_182), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_58), .B(n_180), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_59), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_60), .B(n_180), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_61), .A2(n_155), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_62), .B(n_175), .Y(n_221) );
AND2x2_ASAP7_75t_SL g243 ( .A(n_63), .B(n_183), .Y(n_243) );
XNOR2xp5_ASAP7_75t_L g775 ( .A(n_64), .B(n_776), .Y(n_775) );
XNOR2x1_ASAP7_75t_SL g120 ( .A(n_65), .B(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g563 ( .A(n_65), .B(n_183), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_66), .A2(n_155), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_67), .B(n_177), .Y(n_206) );
AND2x2_ASAP7_75t_SL g215 ( .A(n_68), .B(n_211), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_69), .B(n_175), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_70), .B(n_175), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_71), .A2(n_94), .B1(n_144), .B2(n_155), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_72), .B(n_466), .Y(n_465) );
XNOR2xp5_ASAP7_75t_L g774 ( .A(n_73), .B(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_74), .B(n_177), .Y(n_560) );
INVx1_ASAP7_75t_L g143 ( .A(n_75), .Y(n_143) );
INVx1_ASAP7_75t_L g167 ( .A(n_75), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_76), .B(n_175), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_77), .A2(n_155), .B(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_78), .A2(n_155), .B(n_489), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_79), .A2(n_155), .B(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g535 ( .A(n_80), .B(n_183), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_81), .B(n_182), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_82), .A2(n_86), .B1(n_135), .B2(n_180), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_83), .B(n_180), .Y(n_222) );
INVx1_ASAP7_75t_L g114 ( .A(n_85), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_87), .B(n_175), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_88), .B(n_175), .Y(n_250) );
AND2x2_ASAP7_75t_L g492 ( .A(n_89), .B(n_211), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_90), .A2(n_155), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_93), .B(n_177), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_95), .A2(n_155), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_96), .B(n_177), .Y(n_490) );
OAI22x1_ASAP7_75t_R g447 ( .A1(n_97), .A2(n_448), .B1(n_449), .B2(n_452), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_97), .Y(n_452) );
INVxp67_ASAP7_75t_L g154 ( .A(n_98), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_99), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_100), .B(n_177), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_101), .A2(n_155), .B(n_240), .Y(n_239) );
BUFx2_ASAP7_75t_L g562 ( .A(n_102), .Y(n_562) );
BUFx2_ASAP7_75t_L g454 ( .A(n_103), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_118), .B(n_782), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx3_ASAP7_75t_L g785 ( .A(n_106), .Y(n_785) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_115), .Y(n_107) );
INVx2_ASAP7_75t_SL g467 ( .A(n_108), .Y(n_467) );
INVx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_110), .B(n_460), .Y(n_459) );
AND2x6_ASAP7_75t_SL g475 ( .A(n_110), .B(n_111), .Y(n_475) );
OR2x6_ASAP7_75t_SL g479 ( .A(n_110), .B(n_460), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_111), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_462), .Y(n_118) );
AOI22x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_453), .B1(n_456), .B2(n_461), .Y(n_119) );
OAI22x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_446), .B2(n_447), .Y(n_121) );
OAI22x1_ASAP7_75t_L g780 ( .A1(n_122), .A2(n_474), .B1(n_477), .B2(n_781), .Y(n_780) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OA22x2_ASAP7_75t_L g473 ( .A1(n_123), .A2(n_474), .B1(n_476), .B2(n_480), .Y(n_473) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_323), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_266), .C(n_305), .D(n_312), .Y(n_124) );
OAI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_184), .B1(n_224), .B2(n_233), .C(n_252), .Y(n_125) );
OR2x2_ASAP7_75t_L g396 ( .A(n_126), .B(n_258), .Y(n_396) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g311 ( .A(n_127), .B(n_236), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_127), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_127), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_168), .Y(n_127) );
AND2x4_ASAP7_75t_SL g235 ( .A(n_128), .B(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g257 ( .A(n_128), .Y(n_257) );
AND2x2_ASAP7_75t_L g292 ( .A(n_128), .B(n_265), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_128), .B(n_169), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_128), .B(n_259), .Y(n_344) );
OR2x2_ASAP7_75t_L g422 ( .A(n_128), .B(n_236), .Y(n_422) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_152), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_135), .B1(n_144), .B2(n_150), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_132), .B(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_132), .B(n_154), .Y(n_153) );
NOR3xp33_ASAP7_75t_L g159 ( .A(n_132), .B(n_160), .C(n_162), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_132), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_132), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_132), .A2(n_522), .B(n_523), .Y(n_521) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_133), .B(n_134), .Y(n_183) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_141), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g149 ( .A(n_138), .B(n_140), .Y(n_149) );
AND2x4_ASAP7_75t_L g177 ( .A(n_138), .B(n_166), .Y(n_177) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g155 ( .A(n_142), .B(n_149), .Y(n_155) );
INVx2_ASAP7_75t_L g148 ( .A(n_143), .Y(n_148) );
AND2x6_ASAP7_75t_L g175 ( .A(n_143), .B(n_164), .Y(n_175) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
NOR2x1p5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g528 ( .A(n_156), .Y(n_528) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21x1_ASAP7_75t_L g170 ( .A1(n_157), .A2(n_171), .B(n_181), .Y(n_170) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_157), .A2(n_495), .B(n_501), .Y(n_494) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx4f_ASAP7_75t_L g211 ( .A(n_158), .Y(n_211) );
INVx5_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
AND2x4_ASAP7_75t_L g180 ( .A(n_161), .B(n_163), .Y(n_180) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_166), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g244 ( .A(n_169), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_169), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g270 ( .A(n_169), .Y(n_270) );
OR2x2_ASAP7_75t_L g275 ( .A(n_169), .B(n_259), .Y(n_275) );
AND2x2_ASAP7_75t_L g288 ( .A(n_169), .B(n_246), .Y(n_288) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_169), .Y(n_291) );
INVx1_ASAP7_75t_L g303 ( .A(n_169), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_169), .B(n_257), .Y(n_368) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_179), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .B(n_178), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_175), .B(n_562), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_178), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_178), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_178), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_178), .A2(n_241), .B(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_178), .A2(n_249), .B(n_250), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_178), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_178), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_178), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_178), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_178), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_178), .A2(n_549), .B(n_550), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_178), .A2(n_560), .B(n_561), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_182), .Y(n_193) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_182), .A2(n_247), .B(n_251), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_182), .A2(n_487), .B(n_488), .Y(n_486) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_182), .A2(n_505), .B(n_506), .Y(n_504) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_185), .B(n_195), .Y(n_184) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OR2x2_ASAP7_75t_L g232 ( .A(n_186), .B(n_216), .Y(n_232) );
AND2x4_ASAP7_75t_L g262 ( .A(n_186), .B(n_199), .Y(n_262) );
INVx2_ASAP7_75t_L g296 ( .A(n_186), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_186), .B(n_216), .Y(n_354) );
AND2x2_ASAP7_75t_L g401 ( .A(n_186), .B(n_230), .Y(n_401) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_193), .B(n_194), .Y(n_186) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_187), .A2(n_193), .B(n_194), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_192), .Y(n_187) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_193), .A2(n_217), .B(n_223), .Y(n_216) );
AOI21x1_ASAP7_75t_L g545 ( .A1(n_193), .A2(n_546), .B(n_552), .Y(n_545) );
AOI222xp33_ASAP7_75t_L g389 ( .A1(n_195), .A2(n_261), .B1(n_304), .B2(n_364), .C1(n_390), .C2(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_207), .Y(n_196) );
AND2x2_ASAP7_75t_L g308 ( .A(n_197), .B(n_228), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_197), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g437 ( .A(n_197), .B(n_277), .Y(n_437) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_198), .A2(n_268), .B(n_272), .Y(n_267) );
AND2x2_ASAP7_75t_L g348 ( .A(n_198), .B(n_231), .Y(n_348) );
OR2x2_ASAP7_75t_L g373 ( .A(n_198), .B(n_232), .Y(n_373) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx5_ASAP7_75t_L g227 ( .A(n_199), .Y(n_227) );
AND2x2_ASAP7_75t_L g314 ( .A(n_199), .B(n_296), .Y(n_314) );
AND2x2_ASAP7_75t_L g340 ( .A(n_199), .B(n_216), .Y(n_340) );
OR2x2_ASAP7_75t_L g343 ( .A(n_199), .B(n_230), .Y(n_343) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_199), .Y(n_361) );
AND2x4_ASAP7_75t_SL g418 ( .A(n_199), .B(n_295), .Y(n_418) );
OR2x2_ASAP7_75t_L g427 ( .A(n_199), .B(n_254), .Y(n_427) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g260 ( .A(n_207), .Y(n_260) );
AOI221xp5_ASAP7_75t_SL g378 ( .A1(n_207), .A2(n_262), .B1(n_379), .B2(n_381), .C(n_382), .Y(n_378) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_216), .Y(n_207) );
OR2x2_ASAP7_75t_L g317 ( .A(n_208), .B(n_287), .Y(n_317) );
OR2x2_ASAP7_75t_L g327 ( .A(n_208), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g353 ( .A(n_208), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g359 ( .A(n_208), .B(n_278), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_208), .B(n_342), .Y(n_371) );
INVx2_ASAP7_75t_L g384 ( .A(n_208), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_208), .B(n_262), .Y(n_405) );
AND2x2_ASAP7_75t_L g409 ( .A(n_208), .B(n_231), .Y(n_409) );
AND2x2_ASAP7_75t_L g417 ( .A(n_208), .B(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g230 ( .A(n_209), .Y(n_230) );
AOI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_212), .B(n_215), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_211), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_211), .A2(n_557), .B(n_558), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_216), .B(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g261 ( .A(n_216), .B(n_230), .Y(n_261) );
INVx2_ASAP7_75t_L g278 ( .A(n_216), .Y(n_278) );
AND2x4_ASAP7_75t_L g295 ( .A(n_216), .B(n_296), .Y(n_295) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_216), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_222), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_228), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g407 ( .A(n_226), .B(n_229), .Y(n_407) );
AND2x4_ASAP7_75t_L g253 ( .A(n_227), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g294 ( .A(n_227), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g321 ( .A(n_227), .B(n_261), .Y(n_321) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
AND2x2_ASAP7_75t_L g425 ( .A(n_229), .B(n_426), .Y(n_425) );
BUFx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g277 ( .A(n_230), .B(n_278), .Y(n_277) );
OAI21xp5_ASAP7_75t_SL g297 ( .A1(n_231), .A2(n_298), .B(n_304), .Y(n_297) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_244), .Y(n_234) );
INVx1_ASAP7_75t_SL g351 ( .A(n_235), .Y(n_351) );
AND2x2_ASAP7_75t_L g381 ( .A(n_235), .B(n_291), .Y(n_381) );
AND2x4_ASAP7_75t_L g392 ( .A(n_235), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g258 ( .A(n_236), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g265 ( .A(n_236), .Y(n_265) );
AND2x4_ASAP7_75t_L g271 ( .A(n_236), .B(n_257), .Y(n_271) );
INVx2_ASAP7_75t_L g282 ( .A(n_236), .Y(n_282) );
INVx1_ASAP7_75t_L g331 ( .A(n_236), .Y(n_331) );
OR2x2_ASAP7_75t_L g352 ( .A(n_236), .B(n_336), .Y(n_352) );
OR2x2_ASAP7_75t_L g366 ( .A(n_236), .B(n_246), .Y(n_366) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_236), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_236), .B(n_288), .Y(n_438) );
OR2x6_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
INVx1_ASAP7_75t_L g283 ( .A(n_244), .Y(n_283) );
AND2x2_ASAP7_75t_L g416 ( .A(n_244), .B(n_282), .Y(n_416) );
AND2x2_ASAP7_75t_L g441 ( .A(n_244), .B(n_271), .Y(n_441) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g259 ( .A(n_246), .Y(n_259) );
BUFx3_ASAP7_75t_L g301 ( .A(n_246), .Y(n_301) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_246), .Y(n_328) );
INVx1_ASAP7_75t_L g337 ( .A(n_246), .Y(n_337) );
AOI33xp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_255), .A3(n_260), .B1(n_261), .B2(n_262), .B3(n_263), .Y(n_252) );
AOI21x1_ASAP7_75t_SL g355 ( .A1(n_253), .A2(n_277), .B(n_339), .Y(n_355) );
INVx2_ASAP7_75t_L g385 ( .A(n_253), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_253), .B(n_384), .Y(n_391) );
AND2x2_ASAP7_75t_L g339 ( .A(n_254), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g302 ( .A(n_257), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g403 ( .A(n_258), .Y(n_403) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_259), .Y(n_393) );
OAI32xp33_ASAP7_75t_L g442 ( .A1(n_260), .A2(n_262), .A3(n_438), .B1(n_443), .B2(n_445), .Y(n_442) );
AND2x2_ASAP7_75t_L g360 ( .A(n_261), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_SL g350 ( .A(n_262), .Y(n_350) );
AND2x2_ASAP7_75t_L g415 ( .A(n_262), .B(n_359), .Y(n_415) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OAI221xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_276), .B1(n_279), .B2(n_293), .C(n_297), .Y(n_266) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_270), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_271), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_271), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_271), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g320 ( .A(n_275), .Y(n_320) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR3xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_284), .C(n_289), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_281), .A2(n_343), .B1(n_383), .B2(n_386), .Y(n_382) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g286 ( .A(n_282), .Y(n_286) );
NOR2x1p5_ASAP7_75t_L g300 ( .A(n_282), .B(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI322xp33_ASAP7_75t_L g349 ( .A1(n_285), .A2(n_327), .A3(n_350), .B1(n_351), .B2(n_352), .C1(n_353), .C2(n_355), .Y(n_349) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_287), .A2(n_306), .B(n_307), .C(n_309), .Y(n_305) );
OR2x2_ASAP7_75t_L g397 ( .A(n_287), .B(n_351), .Y(n_397) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g304 ( .A(n_288), .B(n_292), .Y(n_304) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g310 ( .A(n_294), .B(n_311), .Y(n_310) );
INVx3_ASAP7_75t_SL g342 ( .A(n_295), .Y(n_342) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_299), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_SL g346 ( .A(n_302), .Y(n_346) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_303), .Y(n_388) );
OR2x6_ASAP7_75t_SL g443 ( .A(n_306), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI211xp5_ASAP7_75t_L g433 ( .A1(n_311), .A2(n_434), .B(n_435), .C(n_442), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_315), .B(n_318), .C(n_322), .Y(n_312) );
OAI211xp5_ASAP7_75t_SL g324 ( .A1(n_313), .A2(n_325), .B(n_332), .C(n_356), .Y(n_324) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NOR3xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_369), .C(n_413), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_328), .Y(n_420) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g375 ( .A(n_331), .Y(n_375) );
NOR3xp33_ASAP7_75t_SL g332 ( .A(n_333), .B(n_345), .C(n_349), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_338), .B1(n_341), .B2(n_344), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g377 ( .A(n_337), .Y(n_377) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_337), .Y(n_444) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_SL g430 ( .A(n_343), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OR2x2_ASAP7_75t_L g380 ( .A(n_346), .B(n_366), .Y(n_380) );
OR2x2_ASAP7_75t_L g431 ( .A(n_346), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g429 ( .A(n_354), .Y(n_429) );
OR2x2_ASAP7_75t_L g445 ( .A(n_354), .B(n_384), .Y(n_445) );
OAI21xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_362), .Y(n_356) );
OAI31xp33_ASAP7_75t_L g370 ( .A1(n_357), .A2(n_371), .A3(n_372), .B(n_374), .Y(n_370) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g402 ( .A(n_367), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND4xp25_ASAP7_75t_SL g369 ( .A(n_370), .B(n_378), .C(n_389), .D(n_394), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_377), .Y(n_412) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_398), .B1(n_402), .B2(n_404), .C(n_406), .Y(n_394) );
NAND2xp33_ASAP7_75t_SL g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g439 ( .A(n_398), .Y(n_439) );
AND2x2_ASAP7_75t_SL g398 ( .A(n_399), .B(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI21xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g434 ( .A(n_408), .Y(n_434) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_414), .B(n_433), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_417), .B2(n_419), .C(n_423), .Y(n_414) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_428), .B(n_431), .Y(n_423) );
INVxp33_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B1(n_439), .B2(n_440), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVxp33_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
NOR2x1_ASAP7_75t_R g461 ( .A(n_454), .B(n_459), .Y(n_461) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_454), .Y(n_471) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_456), .B(n_465), .C(n_468), .Y(n_464) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_779), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_472), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_774), .Y(n_472) );
CKINVDCx11_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
BUFx4f_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
CKINVDCx11_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
INVx3_ASAP7_75t_SL g781 ( .A(n_480), .Y(n_781) );
AND2x4_ASAP7_75t_SL g480 ( .A(n_481), .B(n_670), .Y(n_480) );
NOR3xp33_ASAP7_75t_SL g481 ( .A(n_482), .B(n_579), .C(n_611), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_507), .B1(n_536), .B2(n_553), .C(n_564), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g542 ( .A(n_485), .B(n_494), .Y(n_542) );
INVx4_ASAP7_75t_L g570 ( .A(n_485), .Y(n_570) );
AND2x4_ASAP7_75t_SL g610 ( .A(n_485), .B(n_544), .Y(n_610) );
BUFx2_ASAP7_75t_L g620 ( .A(n_485), .Y(n_620) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_485), .B(n_625), .Y(n_686) );
AND2x2_ASAP7_75t_L g695 ( .A(n_485), .B(n_623), .Y(n_695) );
OR2x2_ASAP7_75t_L g703 ( .A(n_485), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g729 ( .A(n_485), .B(n_568), .Y(n_729) );
AND2x4_ASAP7_75t_L g748 ( .A(n_485), .B(n_749), .Y(n_748) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
INVx2_ASAP7_75t_SL g661 ( .A(n_493), .Y(n_661) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_502), .Y(n_493) );
AND2x2_ASAP7_75t_L g568 ( .A(n_494), .B(n_545), .Y(n_568) );
INVx2_ASAP7_75t_L g595 ( .A(n_494), .Y(n_595) );
INVx2_ASAP7_75t_L g625 ( .A(n_494), .Y(n_625) );
AND2x2_ASAP7_75t_L g639 ( .A(n_494), .B(n_544), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_500), .Y(n_495) );
AND2x2_ASAP7_75t_L g569 ( .A(n_502), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g592 ( .A(n_502), .Y(n_592) );
BUFx3_ASAP7_75t_L g606 ( .A(n_502), .Y(n_606) );
AND2x2_ASAP7_75t_L g635 ( .A(n_502), .B(n_636), .Y(n_635) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
AND2x4_ASAP7_75t_L g540 ( .A(n_503), .B(n_504), .Y(n_540) );
INVx1_ASAP7_75t_L g641 ( .A(n_507), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .Y(n_507) );
OR2x2_ASAP7_75t_L g752 ( .A(n_508), .B(n_553), .Y(n_752) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g608 ( .A(n_509), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_509), .B(n_518), .Y(n_669) );
OR2x2_ASAP7_75t_L g767 ( .A(n_509), .B(n_689), .Y(n_767) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g578 ( .A(n_510), .B(n_554), .Y(n_578) );
OR2x2_ASAP7_75t_SL g588 ( .A(n_510), .B(n_589), .Y(n_588) );
INVx4_ASAP7_75t_L g599 ( .A(n_510), .Y(n_599) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_510), .Y(n_650) );
NAND2x1_ASAP7_75t_L g656 ( .A(n_510), .B(n_555), .Y(n_656) );
AND2x2_ASAP7_75t_L g681 ( .A(n_510), .B(n_520), .Y(n_681) );
OR2x2_ASAP7_75t_L g702 ( .A(n_510), .B(n_585), .Y(n_702) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g597 ( .A(n_518), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_518), .A2(n_691), .B(n_694), .C(n_696), .Y(n_690) );
AND2x2_ASAP7_75t_L g763 ( .A(n_518), .B(n_539), .Y(n_763) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_527), .Y(n_518) );
INVx1_ASAP7_75t_L g630 ( .A(n_519), .Y(n_630) );
AND2x2_ASAP7_75t_L g700 ( .A(n_519), .B(n_555), .Y(n_700) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g574 ( .A(n_520), .Y(n_574) );
OR2x2_ASAP7_75t_L g589 ( .A(n_520), .B(n_555), .Y(n_589) );
INVx1_ASAP7_75t_L g605 ( .A(n_520), .Y(n_605) );
AND2x2_ASAP7_75t_L g617 ( .A(n_520), .B(n_527), .Y(n_617) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_520), .Y(n_723) );
NOR2x1_ASAP7_75t_SL g554 ( .A(n_527), .B(n_555), .Y(n_554) );
AO21x1_ASAP7_75t_SL g527 ( .A1(n_528), .A2(n_529), .B(n_535), .Y(n_527) );
AO21x2_ASAP7_75t_L g586 ( .A1(n_528), .A2(n_529), .B(n_535), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
INVxp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .Y(n_537) );
OR2x2_ASAP7_75t_L g687 ( .A(n_538), .B(n_622), .Y(n_687) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_539), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g769 ( .A(n_539), .B(n_666), .Y(n_769) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g614 ( .A(n_540), .B(n_595), .Y(n_614) );
AND2x2_ASAP7_75t_L g710 ( .A(n_540), .B(n_623), .Y(n_710) );
INVx1_ASAP7_75t_L g627 ( .A(n_541), .Y(n_627) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g677 ( .A(n_542), .Y(n_677) );
INVx2_ASAP7_75t_L g644 ( .A(n_543), .Y(n_644) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g594 ( .A(n_544), .B(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g624 ( .A(n_544), .Y(n_624) );
INVx1_ASAP7_75t_L g749 ( .A(n_544), .Y(n_749) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_545), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_551), .Y(n_546) );
OR2x2_ASAP7_75t_L g720 ( .A(n_553), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_SL g575 ( .A(n_555), .Y(n_575) );
OR2x2_ASAP7_75t_L g598 ( .A(n_555), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g609 ( .A(n_555), .B(n_585), .Y(n_609) );
AND2x2_ASAP7_75t_L g683 ( .A(n_555), .B(n_599), .Y(n_683) );
BUFx2_ASAP7_75t_L g766 ( .A(n_555), .Y(n_766) );
OR2x6_ASAP7_75t_L g555 ( .A(n_556), .B(n_563), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_571), .B(n_576), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
AND2x2_ASAP7_75t_L g718 ( .A(n_567), .B(n_640), .Y(n_718) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g577 ( .A(n_568), .B(n_570), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_569), .B(n_639), .Y(n_740) );
INVx1_ASAP7_75t_L g770 ( .A(n_569), .Y(n_770) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_570), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_570), .B(n_706), .Y(n_743) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
AND2x4_ASAP7_75t_SL g607 ( .A(n_573), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_573), .B(n_601), .Y(n_754) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_574), .B(n_656), .Y(n_712) );
AND2x2_ASAP7_75t_L g730 ( .A(n_574), .B(n_683), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_575), .B(n_617), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g662 ( .A1(n_575), .A2(n_621), .B(n_663), .C(n_668), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_575), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_577), .A2(n_650), .B1(n_758), .B2(n_764), .C(n_768), .Y(n_757) );
INVx1_ASAP7_75t_SL g745 ( .A(n_578), .Y(n_745) );
OAI221xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_590), .B1(n_596), .B2(n_600), .C(n_787), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_582), .B(n_587), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g655 ( .A(n_584), .Y(n_655) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g629 ( .A(n_585), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g660 ( .A(n_585), .B(n_605), .Y(n_660) );
INVx2_ASAP7_75t_L g693 ( .A(n_585), .Y(n_693) );
INVx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI32xp33_ASAP7_75t_L g744 ( .A1(n_588), .A2(n_635), .A3(n_666), .B1(n_745), .B2(n_746), .Y(n_744) );
OR2x2_ASAP7_75t_L g715 ( .A(n_589), .B(n_702), .Y(n_715) );
INVx1_ASAP7_75t_L g725 ( .A(n_590), .Y(n_725) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx2_ASAP7_75t_L g640 ( .A(n_591), .Y(n_640) );
AND2x2_ASAP7_75t_L g711 ( .A(n_591), .B(n_686), .Y(n_711) );
OR2x2_ASAP7_75t_L g742 ( .A(n_591), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_592), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g636 ( .A(n_595), .Y(n_636) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx2_ASAP7_75t_SL g601 ( .A(n_598), .Y(n_601) );
OR2x2_ASAP7_75t_L g688 ( .A(n_598), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_599), .B(n_617), .Y(n_616) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_599), .B(n_723), .Y(n_722) );
BUFx2_ASAP7_75t_L g735 ( .A(n_599), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_607), .C(n_610), .Y(n_600) );
AND2x2_ASAP7_75t_L g750 ( .A(n_602), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g676 ( .A(n_606), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_606), .B(n_610), .Y(n_697) );
AND2x2_ASAP7_75t_L g728 ( .A(n_606), .B(n_729), .Y(n_728) );
O2A1O1Ixp33_ASAP7_75t_L g738 ( .A1(n_608), .A2(n_739), .B(n_741), .C(n_744), .Y(n_738) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_609), .A2(n_613), .B1(n_615), .B2(n_618), .C1(n_626), .C2(n_628), .Y(n_612) );
AND2x2_ASAP7_75t_L g680 ( .A(n_609), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g613 ( .A(n_610), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_SL g634 ( .A(n_610), .Y(n_634) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_631), .C(n_652), .D(n_662), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_614), .B(n_620), .Y(n_674) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g682 ( .A(n_617), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_SL g689 ( .A(n_617), .Y(n_689) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_619), .A2(n_653), .B(n_657), .C(n_661), .Y(n_652) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_620), .B(n_635), .Y(n_756) );
OR2x2_ASAP7_75t_L g760 ( .A(n_620), .B(n_646), .Y(n_760) );
INVx1_ASAP7_75t_L g733 ( .A(n_621), .Y(n_733) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_SL g667 ( .A(n_624), .Y(n_667) );
INVx1_ASAP7_75t_L g647 ( .A(n_625), .Y(n_647) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_627), .B(n_664), .Y(n_663) );
BUFx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g651 ( .A(n_629), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .A3(n_635), .B1(n_637), .B2(n_641), .C1(n_642), .C2(n_648), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_SL g713 ( .A1(n_634), .A2(n_714), .B(n_715), .C(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g736 ( .A(n_635), .Y(n_736) );
NOR2xp67_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g694 ( .A(n_640), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_646), .Y(n_716) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx3_ASAP7_75t_L g659 ( .A(n_656), .Y(n_659) );
OR2x2_ASAP7_75t_L g727 ( .A(n_656), .B(n_689), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_656), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_SL g759 ( .A(n_660), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_661), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND3xp33_ASAP7_75t_SL g764 ( .A(n_669), .B(n_765), .C(n_767), .Y(n_764) );
NOR3xp33_ASAP7_75t_SL g670 ( .A(n_671), .B(n_708), .C(n_737), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_672), .B(n_690), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B(n_678), .C(n_684), .Y(n_672) );
OAI31xp33_ASAP7_75t_L g717 ( .A1(n_673), .A2(n_695), .A3(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
INVx2_ASAP7_75t_L g732 ( .A(n_680), .Y(n_732) );
INVx1_ASAP7_75t_L g707 ( .A(n_682), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g734 ( .A(n_692), .B(n_735), .Y(n_734) );
INVxp67_ASAP7_75t_L g773 ( .A(n_693), .Y(n_773) );
OAI22xp33_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_698), .B1(n_703), .B2(n_707), .Y(n_696) );
INVx3_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x4_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_702), .Y(n_714) );
OR2x2_ASAP7_75t_L g765 ( .A(n_702), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_709), .B(n_717), .C(n_724), .Y(n_708) );
O2A1O1Ixp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B(n_712), .C(n_713), .Y(n_709) );
INVx2_ASAP7_75t_L g746 ( .A(n_710), .Y(n_746) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B1(n_728), .B2(n_730), .C(n_731), .Y(n_724) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_734), .B2(n_736), .Y(n_731) );
NAND3xp33_ASAP7_75t_SL g737 ( .A(n_738), .B(n_747), .C(n_757), .Y(n_737) );
INVxp33_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_750), .B1(n_753), .B2(n_755), .Y(n_747) );
INVx2_ASAP7_75t_L g761 ( .A(n_748), .Y(n_761) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_758) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OAI22xp33_ASAP7_75t_SL g768 ( .A1(n_767), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND2xp33_ASAP7_75t_SL g779 ( .A(n_774), .B(n_780), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
endmodule