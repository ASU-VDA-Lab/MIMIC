module fake_jpeg_27191_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_32),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_45),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_51),
.B1(n_57),
.B2(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_0),
.B(n_2),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_40),
.C(n_23),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_25),
.B1(n_30),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_24),
.B1(n_17),
.B2(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_33),
.B1(n_21),
.B2(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_40),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_66),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_39),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_89),
.C(n_40),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_69),
.B1(n_46),
.B2(n_48),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_43),
.B1(n_41),
.B2(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_76),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_42),
.B1(n_35),
.B2(n_32),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_77),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_82),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_38),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_85),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_52),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_53),
.Y(n_93)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_38),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_48),
.B1(n_73),
.B2(n_75),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_93),
.A2(n_101),
.B(n_105),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_100),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_86),
.C(n_70),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_89),
.B(n_67),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_51),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_93),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_48),
.B1(n_43),
.B2(n_42),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_84),
.B1(n_71),
.B2(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_40),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_28),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_2),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_49),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_116),
.B1(n_111),
.B2(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_123),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_97),
.B1(n_102),
.B2(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_138),
.B1(n_106),
.B2(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_119),
.B(n_120),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_R g120 ( 
.A(n_108),
.B(n_59),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_62),
.Y(n_123)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_112),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_137),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_65),
.B1(n_73),
.B2(n_83),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_127),
.B1(n_135),
.B2(n_113),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_105),
.B1(n_100),
.B2(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_23),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_136),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_90),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_50),
.B1(n_42),
.B2(n_20),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_20),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_50),
.B1(n_18),
.B2(n_17),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_15),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_14),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_98),
.C(n_95),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_142),
.C(n_154),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_98),
.C(n_95),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_146),
.Y(n_177)
);

BUFx24_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_145),
.B(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_150),
.B(n_18),
.Y(n_180)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_143),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_103),
.C(n_104),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_136),
.B1(n_132),
.B2(n_124),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_111),
.C(n_106),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_18),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_161),
.B1(n_115),
.B2(n_137),
.Y(n_167)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_160),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_2),
.B(n_4),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_117),
.B(n_5),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_171),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_141),
.B(n_118),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_184),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_160),
.B1(n_157),
.B2(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_185),
.C(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_4),
.Y(n_183)
);

OAI322xp33_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_5),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_179),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_156),
.C(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_189),
.B(n_194),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_146),
.B1(n_162),
.B2(n_164),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_158),
.B1(n_153),
.B2(n_148),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_144),
.B1(n_9),
.B2(n_10),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_178),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_144),
.B1(n_9),
.B2(n_10),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_183),
.B1(n_174),
.B2(n_13),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_8),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

NAND2x1p5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_168),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_205),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_169),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_212),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_182),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_191),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_214),
.Y(n_219)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

OA21x2_ASAP7_75t_SL g215 ( 
.A1(n_188),
.A2(n_185),
.B(n_177),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_193),
.B(n_177),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_190),
.C(n_187),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_225),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_205),
.B(n_200),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_209),
.B(n_197),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_190),
.B1(n_202),
.B2(n_192),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_211),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_233),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_223),
.B(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_231),
.B(n_232),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_221),
.B(n_225),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_199),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_236),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_208),
.B(n_206),
.Y(n_236)
);

OAI221xp5_ASAP7_75t_L g239 ( 
.A1(n_237),
.A2(n_234),
.B1(n_232),
.B2(n_238),
.C(n_229),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_229),
.B(n_217),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_217),
.C(n_227),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_11),
.B(n_12),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_SL g247 ( 
.A1(n_246),
.A2(n_245),
.B(n_11),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_13),
.Y(n_248)
);


endmodule