module fake_jpeg_18260_n_65 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_65);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_65;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx5_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx13_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_15),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_19),
.Y(n_23)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_0),
.B(n_1),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_20),
.B(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_15),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_30),
.B1(n_16),
.B2(n_13),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_31),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_18),
.B1(n_20),
.B2(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_12),
.B1(n_14),
.B2(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_28),
.B(n_31),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_35),
.B1(n_38),
.B2(n_14),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_28),
.C(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_47),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_12),
.B(n_32),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_51),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_35),
.C(n_37),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_10),
.C(n_5),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_50),
.B1(n_43),
.B2(n_11),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_46),
.B(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_56),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_5),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_1),
.B(n_2),
.Y(n_61)
);

AOI322xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_53),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_60),
.A2(n_61),
.B(n_58),
.Y(n_62)
);

BUFx24_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_3),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_3),
.Y(n_65)
);


endmodule