module fake_jpeg_1330_n_130 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_26),
.B(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

AO22x1_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_42),
.B1(n_10),
.B2(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_15),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_45),
.Y(n_55)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_3),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_38),
.Y(n_73)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx12_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_15),
.B(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_18),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_51),
.Y(n_76)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_4),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_5),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_19),
.C(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_19),
.B1(n_25),
.B2(n_8),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_6),
.B1(n_56),
.B2(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_27),
.B(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_30),
.Y(n_87)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_30),
.B(n_29),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_28),
.B1(n_48),
.B2(n_42),
.Y(n_82)
);

OAI22x1_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_75),
.B1(n_71),
.B2(n_57),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_29),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_35),
.B1(n_48),
.B2(n_34),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_91),
.B1(n_62),
.B2(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_35),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_87),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_6),
.B(n_7),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_54),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_55),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_101),
.B1(n_75),
.B2(n_71),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_78),
.C(n_87),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.C(n_109),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_83),
.C(n_80),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_90),
.B1(n_82),
.B2(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_110),
.B1(n_98),
.B2(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_102),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_90),
.B(n_89),
.C(n_91),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_68),
.B(n_61),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_76),
.C(n_63),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_113),
.B(n_114),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_99),
.B(n_94),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_116),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_61),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_112),
.A2(n_108),
.B1(n_104),
.B2(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_118),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_79),
.C(n_58),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_88),
.B(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_123),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_70),
.B(n_67),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_R g124 ( 
.A(n_122),
.B(n_118),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_119),
.C(n_77),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_119),
.C(n_86),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_86),
.C(n_57),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_6),
.Y(n_130)
);


endmodule