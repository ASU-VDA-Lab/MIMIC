module fake_ariane_2435_n_2258 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_34, n_404, n_172, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_636, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_2258);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2258;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_1107;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2233;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_2059;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_876;
wire n_791;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_1757;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_2158;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_683;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g655 ( 
.A(n_483),
.Y(n_655)
);

BUFx5_ASAP7_75t_L g656 ( 
.A(n_111),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_575),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_271),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_536),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_605),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_587),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_589),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_415),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_543),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_95),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_420),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_443),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_593),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_8),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_371),
.Y(n_670)
);

BUFx8_ASAP7_75t_SL g671 ( 
.A(n_642),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_230),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_89),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_181),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_481),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_230),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_246),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_541),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_577),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_53),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_650),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_406),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_254),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_67),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_111),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_142),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_576),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_485),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_652),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_91),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_128),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_621),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_632),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_38),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_508),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_351),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_288),
.Y(n_697)
);

CKINVDCx14_ASAP7_75t_R g698 ( 
.A(n_641),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_606),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_445),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_124),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_297),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_79),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_396),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_221),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_640),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_377),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_232),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_61),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_40),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_56),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_190),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_393),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_490),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_349),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_624),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_607),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_633),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_594),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_181),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_34),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_229),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_121),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_93),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_506),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_225),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_540),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_644),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_482),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_645),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_251),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_488),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_224),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_151),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_638),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_625),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_330),
.Y(n_737)
);

CKINVDCx16_ASAP7_75t_R g738 ( 
.A(n_116),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_628),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_514),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_72),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_512),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_597),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_611),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_409),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_627),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_583),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_367),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_1),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_245),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_61),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_385),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_521),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_280),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_434),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_538),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_619),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_466),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_291),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_651),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_643),
.Y(n_761)
);

CKINVDCx16_ASAP7_75t_R g762 ( 
.A(n_17),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_17),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_630),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_518),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_361),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_42),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_513),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_82),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_296),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_93),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_307),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_459),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_170),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_372),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_525),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_473),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_388),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_586),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_596),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_649),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_13),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_578),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_581),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_209),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_617),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_524),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_491),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_364),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_614),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_562),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_591),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_82),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_609),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_239),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_612),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_590),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_223),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_398),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_159),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_358),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_162),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_21),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_120),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_615),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_574),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_634),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_618),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_595),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_598),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_174),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_600),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_132),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_108),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_211),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_610),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_616),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_384),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_646),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_222),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_236),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_201),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_134),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_613),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_460),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_580),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_141),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_603),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_608),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_148),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_177),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_373),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_282),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_307),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_623),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_465),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_515),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_531),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_41),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_584),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_602),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_635),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_78),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_517),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_249),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_302),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_202),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_338),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_435),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_108),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_112),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_497),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_529),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_383),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_192),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_186),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_509),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_268),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_167),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_629),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_478),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_542),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_81),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_527),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_572),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_571),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_262),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_240),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_563),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_26),
.Y(n_870)
);

CKINVDCx16_ASAP7_75t_R g871 ( 
.A(n_592),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_502),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_319),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_141),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_280),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_97),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_566),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_620),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_599),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_622),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_119),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_336),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_118),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_403),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_579),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_184),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_423),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_80),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_192),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_626),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_332),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_149),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_437),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_484),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_648),
.Y(n_895)
);

BUFx8_ASAP7_75t_SL g896 ( 
.A(n_639),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_58),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_159),
.Y(n_898)
);

BUFx10_ASAP7_75t_L g899 ( 
.A(n_334),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_588),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_363),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_242),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_281),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_516),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_601),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_221),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_489),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_285),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_604),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_582),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_138),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_407),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_246),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_339),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_631),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_395),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_115),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_510),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_585),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_647),
.Y(n_920)
);

BUFx10_ASAP7_75t_L g921 ( 
.A(n_13),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_637),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_172),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_636),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_134),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_320),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_295),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_671),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_675),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_656),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_896),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_656),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_656),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_917),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_656),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_760),
.B(n_1),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_656),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_888),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_658),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_665),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_669),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_738),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_674),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_661),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_717),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_762),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_719),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_691),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_697),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_701),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_748),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_814),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_733),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_690),
.Y(n_954)
);

CKINVDCx16_ASAP7_75t_R g955 ( 
.A(n_718),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_870),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_752),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_944),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_930),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_942),
.Y(n_960)
);

OA21x2_ASAP7_75t_L g961 ( 
.A1(n_932),
.A2(n_659),
.B(n_655),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_933),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_944),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_935),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_944),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_946),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_956),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_937),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_939),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_940),
.B(n_807),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_952),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_941),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_947),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_955),
.B(n_871),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_943),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_948),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_949),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_936),
.B(n_909),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_950),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_954),
.B(n_698),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_SL g981 ( 
.A(n_928),
.B(n_814),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_953),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_931),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_938),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_951),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_934),
.B(n_957),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_929),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_945),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_975),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_975),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_978),
.B(n_895),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_961),
.A2(n_763),
.B1(n_708),
.B2(n_710),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_977),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_967),
.B(n_986),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_961),
.A2(n_845),
.B1(n_840),
.B2(n_788),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_982),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_973),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_969),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_985),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_971),
.Y(n_1000)
);

AND2x6_ASAP7_75t_L g1001 ( 
.A(n_980),
.B(n_683),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_959),
.B(n_695),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_972),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_984),
.B(n_792),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_963),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_962),
.B(n_727),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_976),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_983),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_963),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_979),
.Y(n_1010)
);

AO22x2_ASAP7_75t_L g1011 ( 
.A1(n_987),
.A2(n_898),
.B1(n_851),
.B2(n_926),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_958),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_965),
.Y(n_1013)
);

OR2x6_ASAP7_75t_L g1014 ( 
.A(n_988),
.B(n_741),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_960),
.Y(n_1015)
);

AND2x6_ASAP7_75t_L g1016 ( 
.A(n_970),
.B(n_814),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_964),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_966),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_965),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_968),
.B(n_825),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_974),
.Y(n_1021)
);

AND2x6_ASAP7_75t_L g1022 ( 
.A(n_981),
.B(n_751),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_965),
.B(n_660),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_967),
.B(n_724),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_977),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_985),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_983),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_978),
.A2(n_891),
.B1(n_805),
.B2(n_780),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_973),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_987),
.B(n_767),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_978),
.B(n_672),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_978),
.B(n_673),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_998),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_1029),
.B(n_999),
.Y(n_1034)
);

AO22x2_ASAP7_75t_L g1035 ( 
.A1(n_1004),
.A2(n_802),
.B1(n_811),
.B2(n_782),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_993),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_996),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1003),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1007),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1010),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1025),
.B(n_829),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1017),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1002),
.B(n_862),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_994),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1000),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_990),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_1026),
.Y(n_1047)
);

AND2x2_ASAP7_75t_SL g1048 ( 
.A(n_1028),
.B(n_813),
.Y(n_1048)
);

AO22x2_ASAP7_75t_L g1049 ( 
.A1(n_997),
.A2(n_874),
.B1(n_846),
.B2(n_772),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_989),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_1015),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_989),
.Y(n_1052)
);

BUFx8_ASAP7_75t_L g1053 ( 
.A(n_1018),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_1014),
.B(n_798),
.Y(n_1054)
);

AO22x2_ASAP7_75t_L g1055 ( 
.A1(n_991),
.A2(n_1011),
.B1(n_1024),
.B2(n_1031),
.Y(n_1055)
);

AO22x2_ASAP7_75t_L g1056 ( 
.A1(n_1032),
.A2(n_774),
.B1(n_795),
.B2(n_785),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_1008),
.Y(n_1057)
);

AO22x2_ASAP7_75t_L g1058 ( 
.A1(n_995),
.A2(n_800),
.B1(n_823),
.B2(n_821),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1012),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1006),
.B(n_880),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1005),
.Y(n_1061)
);

NAND2xp33_ASAP7_75t_L g1062 ( 
.A(n_1022),
.B(n_676),
.Y(n_1062)
);

BUFx8_ASAP7_75t_L g1063 ( 
.A(n_1001),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1020),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1013),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1013),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1019),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1019),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_992),
.A2(n_657),
.B1(n_790),
.B2(n_666),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1023),
.Y(n_1070)
);

AO22x2_ASAP7_75t_L g1071 ( 
.A1(n_1030),
.A2(n_831),
.B1(n_839),
.B2(n_834),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1009),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1009),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1016),
.Y(n_1074)
);

AO22x2_ASAP7_75t_L g1075 ( 
.A1(n_1027),
.A2(n_856),
.B1(n_892),
.B2(n_873),
.Y(n_1075)
);

AO22x2_ASAP7_75t_L g1076 ( 
.A1(n_1021),
.A2(n_906),
.B1(n_908),
.B2(n_897),
.Y(n_1076)
);

BUFx8_ASAP7_75t_L g1077 ( 
.A(n_1022),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_993),
.Y(n_1078)
);

AO22x2_ASAP7_75t_L g1079 ( 
.A1(n_1029),
.A2(n_925),
.B1(n_911),
.B2(n_890),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_998),
.Y(n_1080)
);

AO22x2_ASAP7_75t_L g1081 ( 
.A1(n_1029),
.A2(n_921),
.B1(n_724),
.B2(n_799),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_1026),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_998),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_993),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_998),
.B(n_677),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_998),
.Y(n_1086)
);

BUFx8_ASAP7_75t_L g1087 ( 
.A(n_999),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_997),
.B(n_923),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_993),
.Y(n_1089)
);

AO22x2_ASAP7_75t_L g1090 ( 
.A1(n_1029),
.A2(n_921),
.B1(n_692),
.B2(n_857),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_998),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_998),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_991),
.A2(n_684),
.B1(n_685),
.B2(n_680),
.Y(n_1093)
);

AO22x2_ASAP7_75t_L g1094 ( 
.A1(n_1029),
.A2(n_861),
.B1(n_894),
.B2(n_819),
.Y(n_1094)
);

AO22x2_ASAP7_75t_L g1095 ( 
.A1(n_1029),
.A2(n_761),
.B1(n_794),
.B2(n_678),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_998),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_998),
.Y(n_1097)
);

OAI221xp5_ASAP7_75t_L g1098 ( 
.A1(n_991),
.A2(n_702),
.B1(n_703),
.B2(n_694),
.C(n_686),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_L g1099 ( 
.A(n_1026),
.B(n_705),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_998),
.B(n_709),
.Y(n_1100)
);

OAI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_991),
.A2(n_720),
.B1(n_721),
.B2(n_712),
.C(n_711),
.Y(n_1101)
);

AO22x2_ASAP7_75t_L g1102 ( 
.A1(n_1029),
.A2(n_768),
.B1(n_789),
.B2(n_745),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_998),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_998),
.B(n_722),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_998),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_994),
.B(n_657),
.Y(n_1106)
);

AO22x2_ASAP7_75t_L g1107 ( 
.A1(n_1029),
.A2(n_826),
.B1(n_837),
.B2(n_681),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_998),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1029),
.B(n_723),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_1026),
.Y(n_1110)
);

AO22x2_ASAP7_75t_L g1111 ( 
.A1(n_1029),
.A2(n_776),
.B1(n_786),
.B2(n_700),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_1029),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_1029),
.Y(n_1113)
);

AO22x2_ASAP7_75t_L g1114 ( 
.A1(n_1029),
.A2(n_716),
.B1(n_668),
.B2(n_670),
.Y(n_1114)
);

INVx8_ASAP7_75t_L g1115 ( 
.A(n_1026),
.Y(n_1115)
);

OAI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_991),
.A2(n_734),
.B1(n_749),
.B2(n_731),
.C(n_726),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_998),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_998),
.B(n_750),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1029),
.B(n_754),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_1029),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_993),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_1029),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_998),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_998),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_998),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1029),
.B(n_759),
.Y(n_1126)
);

AO22x2_ASAP7_75t_L g1127 ( 
.A1(n_1029),
.A2(n_920),
.B1(n_922),
.B2(n_810),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1008),
.B(n_927),
.Y(n_1128)
);

BUFx8_ASAP7_75t_L g1129 ( 
.A(n_999),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1051),
.B(n_769),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1106),
.B(n_770),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1113),
.B(n_663),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1106),
.B(n_771),
.Y(n_1133)
);

NAND2xp33_ASAP7_75t_SL g1134 ( 
.A(n_1057),
.B(n_1047),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1064),
.B(n_793),
.Y(n_1135)
);

NAND2xp33_ASAP7_75t_SL g1136 ( 
.A(n_1082),
.B(n_803),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1044),
.B(n_1034),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1043),
.B(n_1060),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1120),
.B(n_804),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1070),
.B(n_815),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1112),
.B(n_820),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1122),
.B(n_822),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1088),
.B(n_827),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1119),
.B(n_830),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_SL g1145 ( 
.A(n_1110),
.B(n_1128),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1033),
.B(n_833),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1109),
.B(n_843),
.Y(n_1147)
);

NAND2xp33_ASAP7_75t_SL g1148 ( 
.A(n_1038),
.B(n_847),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1053),
.B(n_850),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1048),
.B(n_855),
.Y(n_1150)
);

NAND2xp33_ASAP7_75t_SL g1151 ( 
.A(n_1039),
.B(n_858),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1040),
.B(n_859),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1080),
.B(n_863),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1083),
.B(n_867),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1086),
.B(n_868),
.Y(n_1155)
);

NAND2xp33_ASAP7_75t_SL g1156 ( 
.A(n_1091),
.B(n_875),
.Y(n_1156)
);

NAND2xp33_ASAP7_75t_R g1157 ( 
.A(n_1126),
.B(n_1054),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1092),
.B(n_1096),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1097),
.B(n_876),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1103),
.B(n_881),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1105),
.B(n_883),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1108),
.B(n_886),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_SL g1163 ( 
.A(n_1117),
.B(n_889),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1123),
.B(n_902),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1124),
.B(n_903),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_SL g1166 ( 
.A(n_1125),
.B(n_913),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_SL g1167 ( 
.A(n_1085),
.B(n_919),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1042),
.B(n_707),
.Y(n_1168)
);

NAND2xp33_ASAP7_75t_SL g1169 ( 
.A(n_1100),
.B(n_662),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1115),
.B(n_666),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1058),
.B(n_900),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1115),
.B(n_790),
.Y(n_1172)
);

NAND2xp33_ASAP7_75t_SL g1173 ( 
.A(n_1104),
.B(n_664),
.Y(n_1173)
);

NAND2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1118),
.B(n_916),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1065),
.B(n_918),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1036),
.B(n_901),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1050),
.B(n_899),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1052),
.B(n_899),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1037),
.B(n_905),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1077),
.B(n_679),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1098),
.B(n_1101),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1078),
.B(n_915),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_SL g1183 ( 
.A(n_1066),
.B(n_910),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1041),
.B(n_687),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1067),
.B(n_924),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1068),
.B(n_693),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1087),
.B(n_696),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1084),
.B(n_884),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1129),
.B(n_699),
.Y(n_1189)
);

NAND2xp33_ASAP7_75t_SL g1190 ( 
.A(n_1046),
.B(n_872),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1059),
.B(n_704),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1089),
.B(n_725),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1045),
.B(n_706),
.Y(n_1193)
);

NAND2xp33_ASAP7_75t_SL g1194 ( 
.A(n_1072),
.B(n_887),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1121),
.B(n_713),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1074),
.B(n_777),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1069),
.B(n_714),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1056),
.B(n_779),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1073),
.B(n_914),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1093),
.B(n_728),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1062),
.B(n_860),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1061),
.B(n_729),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1063),
.B(n_730),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1099),
.B(n_732),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1116),
.B(n_735),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1075),
.B(n_736),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1054),
.B(n_737),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1055),
.B(n_739),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1095),
.B(n_740),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1102),
.B(n_742),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1107),
.B(n_743),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_L g1212 ( 
.A(n_1111),
.B(n_744),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1035),
.B(n_0),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1114),
.B(n_746),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1127),
.B(n_747),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1076),
.B(n_864),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1071),
.B(n_753),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1079),
.B(n_0),
.Y(n_1218)
);

NAND2xp33_ASAP7_75t_SL g1219 ( 
.A(n_1094),
.B(n_865),
.Y(n_1219)
);

AND2x2_ASAP7_75t_SL g1220 ( 
.A(n_1049),
.B(n_682),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1090),
.B(n_755),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1081),
.B(n_758),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1051),
.B(n_764),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1051),
.B(n_765),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_SL g1225 ( 
.A(n_1057),
.B(n_766),
.Y(n_1225)
);

NAND2xp33_ASAP7_75t_SL g1226 ( 
.A(n_1057),
.B(n_885),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1051),
.B(n_773),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1051),
.B(n_775),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1051),
.B(n_778),
.Y(n_1229)
);

NAND2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1057),
.B(n_912),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1051),
.B(n_781),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1051),
.B(n_783),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1051),
.B(n_784),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1051),
.B(n_791),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_SL g1235 ( 
.A(n_1057),
.B(n_797),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1051),
.B(n_806),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1051),
.B(n_808),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1064),
.B(n_787),
.Y(n_1238)
);

NAND2xp33_ASAP7_75t_SL g1239 ( 
.A(n_1057),
.B(n_877),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1120),
.B(n_2),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1051),
.B(n_809),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1051),
.B(n_812),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1051),
.B(n_816),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1051),
.B(n_817),
.Y(n_1244)
);

NAND2xp33_ASAP7_75t_SL g1245 ( 
.A(n_1057),
.B(n_818),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1064),
.B(n_828),
.Y(n_1246)
);

NAND2xp33_ASAP7_75t_SL g1247 ( 
.A(n_1057),
.B(n_824),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1064),
.B(n_852),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1051),
.B(n_832),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1051),
.B(n_835),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1051),
.B(n_838),
.Y(n_1251)
);

NAND2xp33_ASAP7_75t_SL g1252 ( 
.A(n_1057),
.B(n_893),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1051),
.B(n_842),
.Y(n_1253)
);

NAND2xp33_ASAP7_75t_SL g1254 ( 
.A(n_1057),
.B(n_854),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1120),
.B(n_2),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1064),
.B(n_836),
.Y(n_1256)
);

NAND2xp33_ASAP7_75t_SL g1257 ( 
.A(n_1057),
.B(n_879),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1120),
.B(n_3),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1120),
.B(n_3),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1051),
.B(n_866),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1051),
.B(n_869),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1051),
.B(n_878),
.Y(n_1262)
);

NAND2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1057),
.B(n_907),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1051),
.B(n_844),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_SL g1265 ( 
.A(n_1057),
.B(n_853),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1051),
.B(n_801),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1064),
.B(n_4),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1051),
.B(n_841),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1051),
.B(n_849),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1051),
.B(n_667),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1064),
.B(n_4),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1051),
.B(n_689),
.Y(n_1272)
);

NAND2xp33_ASAP7_75t_SL g1273 ( 
.A(n_1057),
.B(n_715),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1051),
.B(n_661),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1051),
.B(n_661),
.Y(n_1275)
);

NOR2xp67_ASAP7_75t_L g1276 ( 
.A(n_1138),
.B(n_321),
.Y(n_1276)
);

AO22x2_ASAP7_75t_L g1277 ( 
.A1(n_1209),
.A2(n_757),
.B1(n_848),
.B2(n_756),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1181),
.B(n_5),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1150),
.B(n_5),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1176),
.A2(n_323),
.B(n_322),
.Y(n_1280)
);

BUFx4f_ASAP7_75t_L g1281 ( 
.A(n_1132),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1196),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1158),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1240),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1238),
.B(n_6),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_L g1286 ( 
.A(n_1170),
.B(n_324),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1196),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1246),
.B(n_7),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1134),
.B(n_882),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1148),
.B(n_904),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1248),
.B(n_7),
.Y(n_1291)
);

OA22x2_ASAP7_75t_L g1292 ( 
.A1(n_1217),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1267),
.A2(n_796),
.B(n_688),
.C(n_11),
.Y(n_1293)
);

NOR2x1_ASAP7_75t_SL g1294 ( 
.A(n_1271),
.B(n_688),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1179),
.A2(n_326),
.B(n_325),
.Y(n_1295)
);

NAND2xp33_ASAP7_75t_L g1296 ( 
.A(n_1167),
.B(n_688),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1182),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1137),
.B(n_9),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1184),
.A2(n_1143),
.B(n_1133),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1188),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1131),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_1301)
);

AOI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1192),
.A2(n_796),
.B(n_328),
.Y(n_1302)
);

INVx6_ASAP7_75t_L g1303 ( 
.A(n_1132),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1168),
.A2(n_329),
.B(n_327),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1198),
.A2(n_796),
.A3(n_333),
.B(n_335),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1201),
.A2(n_1193),
.B(n_1256),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_SL g1307 ( 
.A1(n_1146),
.A2(n_1154),
.B(n_1171),
.Y(n_1307)
);

AOI221x1_ASAP7_75t_L g1308 ( 
.A1(n_1219),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.C(n_16),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1135),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1212),
.B(n_18),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1169),
.A2(n_337),
.B(n_331),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1152),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1255),
.B(n_18),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_SL g1314 ( 
.A1(n_1216),
.A2(n_19),
.B(n_20),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_1136),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1151),
.B(n_19),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1274),
.A2(n_341),
.B(n_340),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1208),
.A2(n_343),
.A3(n_344),
.B(n_342),
.Y(n_1318)
);

AOI21x1_ASAP7_75t_SL g1319 ( 
.A1(n_1173),
.A2(n_20),
.B(n_21),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1157),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1275),
.A2(n_346),
.B(n_345),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1258),
.B(n_22),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1210),
.A2(n_348),
.A3(n_350),
.B(n_347),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1259),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1145),
.Y(n_1325)
);

AOI221x1_ASAP7_75t_L g1326 ( 
.A1(n_1218),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.C(n_26),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1140),
.A2(n_23),
.B(n_24),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1174),
.A2(n_353),
.B(n_352),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1204),
.A2(n_355),
.B(n_354),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1213),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1153),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1220),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1205),
.A2(n_25),
.B(n_27),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1155),
.Y(n_1334)
);

INVxp67_ASAP7_75t_L g1335 ( 
.A(n_1264),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1159),
.Y(n_1336)
);

INVx5_ASAP7_75t_L g1337 ( 
.A(n_1187),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1144),
.B(n_28),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1211),
.B(n_28),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1214),
.B(n_29),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1160),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1195),
.A2(n_1200),
.B(n_1202),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1161),
.A2(n_357),
.B(n_356),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1180),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1215),
.B(n_30),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1206),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1162),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1207),
.A2(n_1222),
.B(n_1221),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1191),
.A2(n_360),
.B(n_359),
.Y(n_1349)
);

CKINVDCx6p67_ASAP7_75t_R g1350 ( 
.A(n_1189),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1147),
.B(n_32),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1164),
.A2(n_365),
.B(n_362),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1197),
.B(n_33),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1165),
.A2(n_368),
.B(n_366),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1156),
.B(n_34),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1177),
.A2(n_370),
.B(n_369),
.Y(n_1356)
);

OR2x6_ASAP7_75t_L g1357 ( 
.A(n_1149),
.B(n_35),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1163),
.B(n_35),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1166),
.A2(n_375),
.A3(n_376),
.B(n_374),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1172),
.B(n_36),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1266),
.A2(n_379),
.B(n_378),
.Y(n_1361)
);

AOI21x1_ASAP7_75t_SL g1362 ( 
.A1(n_1190),
.A2(n_37),
.B(n_38),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1268),
.A2(n_381),
.B(n_380),
.Y(n_1363)
);

AO31x2_ASAP7_75t_L g1364 ( 
.A1(n_1175),
.A2(n_386),
.A3(n_387),
.B(n_382),
.Y(n_1364)
);

AOI21xp33_ASAP7_75t_L g1365 ( 
.A1(n_1269),
.A2(n_37),
.B(n_39),
.Y(n_1365)
);

AO31x2_ASAP7_75t_L g1366 ( 
.A1(n_1183),
.A2(n_390),
.A3(n_391),
.B(n_389),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1141),
.B(n_39),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1142),
.B(n_40),
.Y(n_1368)
);

AOI221x1_ASAP7_75t_L g1369 ( 
.A1(n_1185),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.C(n_44),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1273),
.A2(n_394),
.B(n_392),
.Y(n_1370)
);

O2A1O1Ixp5_ASAP7_75t_L g1371 ( 
.A1(n_1223),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1139),
.B(n_45),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1186),
.A2(n_1265),
.B(n_1194),
.C(n_1199),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1224),
.A2(n_399),
.B(n_397),
.Y(n_1374)
);

AO32x2_ASAP7_75t_L g1375 ( 
.A1(n_1178),
.A2(n_48),
.A3(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1225),
.B(n_46),
.Y(n_1376)
);

NAND3x1_ASAP7_75t_L g1377 ( 
.A(n_1203),
.B(n_49),
.C(n_48),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1130),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1227),
.A2(n_401),
.B(n_400),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1270),
.B(n_47),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1228),
.A2(n_1231),
.B(n_1229),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1226),
.B(n_50),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1272),
.B(n_50),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1232),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1230),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1233),
.B(n_51),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1263),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1235),
.B(n_52),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1282),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1283),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1332),
.A2(n_1236),
.B1(n_1237),
.B2(n_1234),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1281),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1297),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1337),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1280),
.A2(n_1242),
.B(n_1241),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1295),
.A2(n_1244),
.B(n_1243),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1284),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1325),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1279),
.B(n_1250),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1387),
.B(n_1239),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1324),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1278),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1331),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1300),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1287),
.B(n_1249),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1335),
.B(n_1320),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1378),
.B(n_1315),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1304),
.A2(n_1253),
.B(n_1251),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1307),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1344),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1312),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1330),
.A2(n_1261),
.B1(n_1262),
.B2(n_1260),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1302),
.A2(n_404),
.B(n_402),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1350),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1296),
.A2(n_1247),
.B(n_1245),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1285),
.A2(n_1254),
.B1(n_1257),
.B2(n_1252),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1288),
.B(n_54),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1384),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1336),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1334),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1298),
.B(n_405),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1313),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1277),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1361),
.A2(n_410),
.B(n_408),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1294),
.A2(n_412),
.B(n_411),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1291),
.B(n_55),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1347),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1276),
.A2(n_414),
.B(n_413),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1380),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1360),
.B(n_416),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1292),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1322),
.A2(n_63),
.B1(n_60),
.B2(n_62),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1286),
.B(n_417),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1383),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1381),
.Y(n_1435)
);

AND2x2_ASAP7_75t_SL g1436 ( 
.A(n_1388),
.B(n_62),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1311),
.A2(n_419),
.B(n_418),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1305),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1305),
.Y(n_1439)
);

OAI222xp33_ASAP7_75t_L g1440 ( 
.A1(n_1310),
.A2(n_65),
.B1(n_67),
.B2(n_63),
.C1(n_64),
.C2(n_66),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1338),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1373),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1353),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1349),
.A2(n_1354),
.B(n_1352),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1317),
.A2(n_422),
.B(n_421),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1357),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1306),
.A2(n_68),
.B(n_69),
.Y(n_1447)
);

AO31x2_ASAP7_75t_L g1448 ( 
.A1(n_1293),
.A2(n_425),
.A3(n_426),
.B(n_424),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1333),
.A2(n_70),
.B(n_71),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1299),
.A2(n_71),
.B(n_72),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1351),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1321),
.A2(n_428),
.B(n_427),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1372),
.B(n_73),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1342),
.A2(n_430),
.B(n_429),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1367),
.A2(n_75),
.B(n_76),
.C(n_74),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1314),
.A2(n_432),
.B(n_431),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1355),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1339),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1386),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1340),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1348),
.B(n_76),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1356),
.A2(n_1328),
.B(n_1362),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1345),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1358),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_SL g1465 ( 
.A1(n_1327),
.A2(n_1379),
.B(n_1374),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1289),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1371),
.A2(n_1290),
.B(n_1369),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1368),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.C(n_80),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1376),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1382),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1370),
.A2(n_436),
.B(n_433),
.Y(n_1471)
);

INVx8_ASAP7_75t_L g1472 ( 
.A(n_1377),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1309),
.A2(n_77),
.B(n_81),
.Y(n_1473)
);

A2O1A1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1301),
.A2(n_1316),
.B(n_1346),
.C(n_1385),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1365),
.A2(n_1343),
.B(n_1329),
.C(n_1341),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1308),
.A2(n_85),
.B(n_86),
.C(n_84),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1375),
.B(n_83),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1326),
.A2(n_86),
.B1(n_83),
.B2(n_85),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1375),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1363),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1319),
.A2(n_439),
.B(n_438),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1318),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1318),
.Y(n_1483)
);

BUFx4f_ASAP7_75t_SL g1484 ( 
.A(n_1323),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1323),
.A2(n_87),
.B(n_88),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1359),
.A2(n_1366),
.B(n_1364),
.Y(n_1486)
);

AND2x6_ASAP7_75t_L g1487 ( 
.A(n_1359),
.B(n_1364),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_SL g1488 ( 
.A(n_1366),
.B(n_87),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1283),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1281),
.B(n_90),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1278),
.A2(n_441),
.B(n_440),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1324),
.B(n_91),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1280),
.A2(n_444),
.B(n_442),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1303),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1283),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_SL g1496 ( 
.A(n_1281),
.B(n_446),
.Y(n_1496)
);

OAI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1278),
.A2(n_95),
.B1(n_92),
.B2(n_94),
.C(n_96),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1281),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1280),
.A2(n_448),
.B(n_447),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1280),
.A2(n_450),
.B(n_449),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1278),
.A2(n_92),
.B(n_97),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1303),
.Y(n_1502)
);

INVx5_ASAP7_75t_SL g1503 ( 
.A(n_1350),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1325),
.B(n_98),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1435),
.B(n_98),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1393),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1404),
.Y(n_1507)
);

BUFx2_ASAP7_75t_SL g1508 ( 
.A(n_1392),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1390),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1409),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1489),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1411),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1495),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1494),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1443),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1438),
.A2(n_452),
.B(n_451),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1502),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1420),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1410),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1401),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1458),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1455),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1498),
.B(n_99),
.Y(n_1523)
);

INVxp67_ASAP7_75t_SL g1524 ( 
.A(n_1403),
.Y(n_1524)
);

INVxp33_ASAP7_75t_L g1525 ( 
.A(n_1407),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1463),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1429),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1397),
.B(n_100),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1434),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1419),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1394),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1389),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1451),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1430),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1444),
.A2(n_454),
.B(n_453),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1418),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1398),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1414),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1422),
.B(n_101),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1406),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1402),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1479),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1472),
.B(n_455),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1490),
.B(n_1436),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1454),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1446),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1459),
.B(n_102),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1465),
.A2(n_102),
.B(n_103),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1437),
.A2(n_103),
.B(n_104),
.Y(n_1549)
);

INVx5_ASAP7_75t_L g1550 ( 
.A(n_1503),
.Y(n_1550)
);

BUFx4f_ASAP7_75t_SL g1551 ( 
.A(n_1469),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1417),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1477),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1464),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1492),
.B(n_104),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1421),
.B(n_105),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1461),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1462),
.A2(n_457),
.B(n_456),
.Y(n_1558)
);

OA21x2_ASAP7_75t_L g1559 ( 
.A1(n_1439),
.A2(n_461),
.B(n_458),
.Y(n_1559)
);

AOI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1483),
.A2(n_463),
.B(n_462),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1426),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1470),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1460),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1405),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1447),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1453),
.B(n_105),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1453),
.B(n_106),
.Y(n_1567)
);

BUFx5_ASAP7_75t_L g1568 ( 
.A(n_1487),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1456),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1501),
.B(n_107),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1466),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1503),
.B(n_107),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1450),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1441),
.B(n_109),
.Y(n_1574)
);

CKINVDCx11_ASAP7_75t_R g1575 ( 
.A(n_1433),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1536),
.B(n_1546),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1537),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1554),
.B(n_1400),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1543),
.B(n_1415),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1517),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1509),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1518),
.B(n_1504),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_R g1583 ( 
.A(n_1543),
.B(n_1399),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1550),
.B(n_1408),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1540),
.B(n_1416),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1519),
.Y(n_1586)
);

NAND2xp33_ASAP7_75t_R g1587 ( 
.A(n_1556),
.B(n_1481),
.Y(n_1587)
);

NAND2xp33_ASAP7_75t_SL g1588 ( 
.A(n_1570),
.B(n_1478),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1550),
.Y(n_1589)
);

XNOR2xp5_ASAP7_75t_L g1590 ( 
.A(n_1525),
.B(n_1412),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1553),
.B(n_1476),
.Y(n_1591)
);

BUFx10_ASAP7_75t_L g1592 ( 
.A(n_1523),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_R g1593 ( 
.A(n_1544),
.B(n_1486),
.Y(n_1593)
);

NAND2xp33_ASAP7_75t_R g1594 ( 
.A(n_1566),
.B(n_1473),
.Y(n_1594)
);

NAND2xp33_ASAP7_75t_R g1595 ( 
.A(n_1567),
.B(n_1449),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1550),
.B(n_1395),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1520),
.B(n_1431),
.Y(n_1597)
);

XNOR2xp5_ASAP7_75t_L g1598 ( 
.A(n_1514),
.B(n_1423),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1551),
.B(n_1440),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1534),
.B(n_1396),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1524),
.B(n_1485),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_R g1602 ( 
.A(n_1505),
.B(n_1496),
.Y(n_1602)
);

XNOR2xp5_ASAP7_75t_L g1603 ( 
.A(n_1539),
.B(n_1391),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1515),
.B(n_1457),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1564),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1532),
.B(n_1530),
.Y(n_1606)
);

CKINVDCx11_ASAP7_75t_R g1607 ( 
.A(n_1575),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_R g1608 ( 
.A(n_1538),
.B(n_1484),
.Y(n_1608)
);

OR2x6_ASAP7_75t_L g1609 ( 
.A(n_1508),
.B(n_1442),
.Y(n_1609)
);

CKINVDCx16_ASAP7_75t_R g1610 ( 
.A(n_1528),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1531),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1541),
.B(n_1468),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1512),
.Y(n_1613)
);

NAND2xp33_ASAP7_75t_R g1614 ( 
.A(n_1572),
.B(n_1467),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1571),
.Y(n_1615)
);

NAND2xp33_ASAP7_75t_R g1616 ( 
.A(n_1557),
.B(n_1482),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1562),
.B(n_1448),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_R g1618 ( 
.A(n_1555),
.B(n_1432),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1533),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1586),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1606),
.B(n_1510),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1619),
.B(n_1510),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1576),
.B(n_1507),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1581),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1605),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1613),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1577),
.B(n_1511),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1601),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1578),
.B(n_1610),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1604),
.Y(n_1630)
);

AND2x4_ASAP7_75t_SL g1631 ( 
.A(n_1592),
.B(n_1521),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1585),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1591),
.B(n_1513),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1582),
.B(n_1561),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_1616),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1617),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1597),
.B(n_1542),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1612),
.B(n_1552),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1584),
.B(n_1526),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1614),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1588),
.A2(n_1573),
.B1(n_1574),
.B2(n_1565),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1618),
.A2(n_1488),
.B1(n_1487),
.B2(n_1568),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1587),
.Y(n_1643)
);

BUFx2_ASAP7_75t_SL g1644 ( 
.A(n_1615),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1600),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1596),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1579),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1611),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1599),
.A2(n_1563),
.B1(n_1497),
.B2(n_1487),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1579),
.Y(n_1650)
);

NAND2x1p5_ASAP7_75t_L g1651 ( 
.A(n_1589),
.B(n_1529),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1608),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1593),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1589),
.B(n_1527),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1590),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1598),
.B(n_1547),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1609),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1609),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1580),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1603),
.Y(n_1660)
);

NOR2xp67_ASAP7_75t_L g1661 ( 
.A(n_1583),
.B(n_1548),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1607),
.B(n_1568),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1594),
.B(n_1568),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1595),
.B(n_1506),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1628),
.B(n_1630),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1625),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1640),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1629),
.B(n_1569),
.Y(n_1668)
);

AOI33xp33_ASAP7_75t_L g1669 ( 
.A1(n_1641),
.A2(n_1522),
.A3(n_112),
.B1(n_114),
.B2(n_109),
.B3(n_110),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1649),
.A2(n_1602),
.B1(n_1474),
.B2(n_1475),
.C(n_1427),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_1643),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1622),
.B(n_1623),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1646),
.B(n_1545),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1627),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1624),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1631),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1633),
.B(n_1632),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1659),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1648),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1637),
.Y(n_1680)
);

INVx4_ASAP7_75t_L g1681 ( 
.A(n_1662),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1661),
.A2(n_1549),
.B1(n_1425),
.B2(n_1491),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1657),
.A2(n_1471),
.B1(n_1559),
.B2(n_1516),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1626),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1658),
.Y(n_1685)
);

INVxp67_ASAP7_75t_SL g1686 ( 
.A(n_1650),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1639),
.B(n_1560),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1620),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1652),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1634),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1645),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1636),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1664),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1642),
.A2(n_1428),
.B1(n_1559),
.B2(n_1480),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1638),
.Y(n_1695)
);

AND2x4_ASAP7_75t_SL g1696 ( 
.A(n_1663),
.B(n_1535),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1653),
.B(n_113),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1647),
.B(n_1558),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1635),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1644),
.B(n_1493),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1654),
.B(n_1499),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_L g1702 ( 
.A(n_1655),
.B(n_1656),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1651),
.B(n_1660),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1621),
.B(n_1500),
.Y(n_1704)
);

OR2x6_ASAP7_75t_L g1705 ( 
.A(n_1662),
.B(n_1413),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1624),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1621),
.B(n_117),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1624),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1621),
.B(n_118),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1650),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1626),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1620),
.Y(n_1712)
);

AOI211xp5_ASAP7_75t_L g1713 ( 
.A1(n_1640),
.A2(n_1445),
.B(n_1452),
.C(n_1424),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1640),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1621),
.B(n_119),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1624),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1621),
.B(n_120),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1628),
.B(n_122),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1628),
.B(n_122),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1684),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1672),
.B(n_1710),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1699),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1665),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1667),
.B(n_123),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1710),
.B(n_123),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1681),
.B(n_1666),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1675),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1674),
.B(n_124),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1686),
.B(n_125),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1714),
.B(n_125),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1668),
.B(n_126),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1706),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1708),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1716),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1690),
.B(n_126),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1677),
.B(n_127),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1671),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1691),
.B(n_127),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1669),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1693),
.B(n_129),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1680),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1711),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1689),
.B(n_130),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1695),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1692),
.Y(n_1745)
);

NAND4xp25_ASAP7_75t_L g1746 ( 
.A(n_1670),
.B(n_135),
.C(n_132),
.D(n_133),
.Y(n_1746)
);

INVxp67_ASAP7_75t_SL g1747 ( 
.A(n_1697),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1685),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1698),
.Y(n_1749)
);

INVxp67_ASAP7_75t_L g1750 ( 
.A(n_1702),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1678),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1704),
.B(n_135),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1718),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1719),
.B(n_136),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1707),
.B(n_136),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1673),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1676),
.B(n_137),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1688),
.B(n_137),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1688),
.B(n_138),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1712),
.B(n_139),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1712),
.B(n_139),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1679),
.B(n_140),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1703),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1709),
.B(n_142),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1701),
.Y(n_1765)
);

NOR2x1_ASAP7_75t_L g1766 ( 
.A(n_1715),
.B(n_143),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1717),
.B(n_144),
.Y(n_1767)
);

INVxp67_ASAP7_75t_SL g1768 ( 
.A(n_1700),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1696),
.B(n_144),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1705),
.B(n_145),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1687),
.Y(n_1771)
);

CKINVDCx11_ASAP7_75t_R g1772 ( 
.A(n_1683),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1694),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1682),
.B(n_146),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1713),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1667),
.B(n_147),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1684),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1672),
.B(n_148),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_SL g1779 ( 
.A(n_1679),
.B(n_149),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1674),
.B(n_150),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1672),
.B(n_150),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1667),
.B(n_151),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1666),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1684),
.Y(n_1784)
);

AND2x6_ASAP7_75t_SL g1785 ( 
.A(n_1707),
.B(n_152),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1672),
.B(n_152),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1699),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1684),
.Y(n_1788)
);

NAND2xp67_ASAP7_75t_SL g1789 ( 
.A(n_1700),
.B(n_153),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1684),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1684),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1775),
.B(n_154),
.Y(n_1792)
);

NAND2xp33_ASAP7_75t_SL g1793 ( 
.A(n_1721),
.B(n_154),
.Y(n_1793)
);

OAI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1746),
.A2(n_1774),
.B1(n_1750),
.B2(n_1773),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1737),
.B(n_155),
.Y(n_1795)
);

NAND2x1_ASAP7_75t_L g1796 ( 
.A(n_1751),
.B(n_156),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1751),
.Y(n_1797)
);

CKINVDCx20_ASAP7_75t_R g1798 ( 
.A(n_1767),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1752),
.B(n_1726),
.Y(n_1799)
);

NAND2xp33_ASAP7_75t_SL g1800 ( 
.A(n_1725),
.B(n_156),
.Y(n_1800)
);

AO221x2_ASAP7_75t_L g1801 ( 
.A1(n_1724),
.A2(n_160),
.B1(n_157),
.B2(n_158),
.C(n_161),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1752),
.B(n_157),
.Y(n_1802)
);

AO221x2_ASAP7_75t_L g1803 ( 
.A1(n_1730),
.A2(n_161),
.B1(n_158),
.B2(n_160),
.C(n_162),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1785),
.B(n_163),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1744),
.B(n_164),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_R g1806 ( 
.A(n_1779),
.B(n_165),
.Y(n_1806)
);

AO221x2_ASAP7_75t_L g1807 ( 
.A1(n_1782),
.A2(n_169),
.B1(n_166),
.B2(n_168),
.C(n_170),
.Y(n_1807)
);

NAND2xp33_ASAP7_75t_SL g1808 ( 
.A(n_1738),
.B(n_166),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1720),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1723),
.B(n_171),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1787),
.B(n_171),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1736),
.B(n_173),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1728),
.B(n_1741),
.Y(n_1813)
);

AO221x2_ASAP7_75t_L g1814 ( 
.A1(n_1755),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.C(n_178),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1740),
.B(n_175),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1727),
.B(n_176),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1748),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_1778),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1732),
.B(n_179),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1749),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1777),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_L g1822 ( 
.A(n_1789),
.B(n_1776),
.Y(n_1822)
);

BUFx4f_ASAP7_75t_L g1823 ( 
.A(n_1758),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1766),
.B(n_180),
.Y(n_1824)
);

NOR4xp25_ASAP7_75t_SL g1825 ( 
.A(n_1771),
.B(n_183),
.C(n_180),
.D(n_182),
.Y(n_1825)
);

NOR2x1_ASAP7_75t_L g1826 ( 
.A(n_1776),
.B(n_182),
.Y(n_1826)
);

AO221x2_ASAP7_75t_L g1827 ( 
.A1(n_1765),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.C(n_186),
.Y(n_1827)
);

OAI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1780),
.A2(n_188),
.B1(n_189),
.B2(n_187),
.Y(n_1828)
);

NOR4xp25_ASAP7_75t_SL g1829 ( 
.A(n_1768),
.B(n_188),
.C(n_185),
.D(n_187),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1763),
.Y(n_1830)
);

AO221x2_ASAP7_75t_L g1831 ( 
.A1(n_1772),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.C(n_193),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1733),
.B(n_191),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1762),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1770),
.B(n_193),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1784),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1734),
.B(n_194),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1781),
.Y(n_1837)
);

OR2x6_ASAP7_75t_L g1838 ( 
.A(n_1786),
.B(n_195),
.Y(n_1838)
);

AO221x2_ASAP7_75t_L g1839 ( 
.A1(n_1735),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_1839)
);

AO221x2_ASAP7_75t_L g1840 ( 
.A1(n_1753),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1759),
.Y(n_1841)
);

AO221x2_ASAP7_75t_L g1842 ( 
.A1(n_1739),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1788),
.B(n_203),
.Y(n_1843)
);

AO221x2_ASAP7_75t_L g1844 ( 
.A1(n_1790),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.C(n_207),
.Y(n_1844)
);

A2O1A1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1761),
.A2(n_213),
.B(n_222),
.C(n_205),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1791),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1731),
.B(n_206),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1743),
.B(n_1769),
.Y(n_1848)
);

AO221x2_ASAP7_75t_L g1849 ( 
.A1(n_1729),
.A2(n_211),
.B1(n_208),
.B2(n_210),
.C(n_212),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1764),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_1850)
);

OAI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1754),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1760),
.B(n_217),
.Y(n_1852)
);

INVxp33_ASAP7_75t_SL g1853 ( 
.A(n_1757),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1745),
.B(n_218),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1742),
.B(n_219),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1756),
.A2(n_225),
.B1(n_220),
.B2(n_224),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1721),
.B(n_226),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1775),
.B(n_226),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1785),
.Y(n_1859)
);

AO221x2_ASAP7_75t_L g1860 ( 
.A1(n_1775),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.C(n_231),
.Y(n_1860)
);

OAI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1775),
.A2(n_231),
.B1(n_227),
.B2(n_228),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_R g1862 ( 
.A(n_1785),
.B(n_232),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1775),
.B(n_233),
.Y(n_1863)
);

OAI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1775),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_1864)
);

O2A1O1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1739),
.A2(n_237),
.B(n_234),
.C(n_235),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_R g1866 ( 
.A(n_1785),
.B(n_237),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1775),
.B(n_238),
.Y(n_1867)
);

INVxp33_ASAP7_75t_SL g1868 ( 
.A(n_1779),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1783),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1746),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_1870)
);

BUFx2_ASAP7_75t_L g1871 ( 
.A(n_1737),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1775),
.B(n_241),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1747),
.B(n_243),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1775),
.B(n_244),
.Y(n_1874)
);

NAND2xp33_ASAP7_75t_R g1875 ( 
.A(n_1776),
.B(n_244),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1747),
.B(n_245),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1722),
.Y(n_1877)
);

INVx3_ASAP7_75t_SL g1878 ( 
.A(n_1859),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1809),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1869),
.B(n_247),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1798),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1853),
.B(n_247),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1868),
.B(n_248),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1833),
.B(n_1792),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1797),
.B(n_248),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1821),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1818),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1837),
.B(n_249),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1835),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1871),
.B(n_250),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1858),
.B(n_252),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1848),
.B(n_253),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1817),
.B(n_254),
.Y(n_1893)
);

NOR2x1_ASAP7_75t_L g1894 ( 
.A(n_1826),
.B(n_255),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1862),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1846),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1854),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1822),
.Y(n_1898)
);

HB1xp67_ASAP7_75t_L g1899 ( 
.A(n_1813),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1866),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1855),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1795),
.B(n_255),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1831),
.A2(n_256),
.B(n_257),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1830),
.B(n_256),
.Y(n_1904)
);

CKINVDCx16_ASAP7_75t_R g1905 ( 
.A(n_1875),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1877),
.Y(n_1906)
);

OR2x6_ASAP7_75t_L g1907 ( 
.A(n_1796),
.B(n_257),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1857),
.B(n_1799),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1831),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1811),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1873),
.B(n_258),
.Y(n_1911)
);

AO21x2_ASAP7_75t_L g1912 ( 
.A1(n_1863),
.A2(n_259),
.B(n_260),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1876),
.B(n_261),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1810),
.B(n_261),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1843),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1836),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1842),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1805),
.B(n_263),
.Y(n_1918)
);

AO21x2_ASAP7_75t_L g1919 ( 
.A1(n_1867),
.A2(n_264),
.B(n_265),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1816),
.B(n_265),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1819),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1832),
.B(n_266),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_SL g1923 ( 
.A1(n_1804),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1838),
.B(n_267),
.Y(n_1924)
);

INVx2_ASAP7_75t_SL g1925 ( 
.A(n_1841),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1872),
.B(n_269),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1820),
.B(n_269),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1794),
.B(n_270),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1874),
.Y(n_1929)
);

INVx1_ASAP7_75t_SL g1930 ( 
.A(n_1806),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1815),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1852),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1847),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1840),
.B(n_272),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1842),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1849),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1824),
.Y(n_1937)
);

OAI21xp33_ASAP7_75t_L g1938 ( 
.A1(n_1870),
.A2(n_273),
.B(n_274),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1849),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1812),
.B(n_275),
.Y(n_1940)
);

OAI21x1_ASAP7_75t_L g1941 ( 
.A1(n_1802),
.A2(n_1834),
.B(n_1856),
.Y(n_1941)
);

INVx4_ASAP7_75t_L g1942 ( 
.A(n_1801),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1840),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1827),
.B(n_275),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1839),
.B(n_276),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1839),
.B(n_276),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1844),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1803),
.B(n_277),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1807),
.B(n_277),
.Y(n_1949)
);

INVx1_ASAP7_75t_SL g1950 ( 
.A(n_1808),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1860),
.A2(n_281),
.B1(n_278),
.B2(n_279),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1814),
.B(n_278),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1850),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1851),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1845),
.B(n_279),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1793),
.Y(n_1956)
);

INVx1_ASAP7_75t_SL g1957 ( 
.A(n_1800),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1829),
.B(n_1825),
.Y(n_1958)
);

NOR2x1_ASAP7_75t_L g1959 ( 
.A(n_1828),
.B(n_283),
.Y(n_1959)
);

BUFx12f_ASAP7_75t_L g1960 ( 
.A(n_1861),
.Y(n_1960)
);

INVx1_ASAP7_75t_SL g1961 ( 
.A(n_1864),
.Y(n_1961)
);

OA21x2_ASAP7_75t_L g1962 ( 
.A1(n_1865),
.A2(n_283),
.B(n_284),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1809),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1797),
.B(n_284),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1833),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1798),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1869),
.B(n_285),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1833),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1798),
.Y(n_1969)
);

INVx3_ASAP7_75t_SL g1970 ( 
.A(n_1859),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1869),
.B(n_286),
.Y(n_1971)
);

INVx4_ASAP7_75t_L g1972 ( 
.A(n_1838),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1797),
.B(n_286),
.Y(n_1973)
);

NOR2x1_ASAP7_75t_L g1974 ( 
.A(n_1826),
.B(n_287),
.Y(n_1974)
);

NAND3x1_ASAP7_75t_SL g1975 ( 
.A(n_1826),
.B(n_287),
.C(n_288),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1797),
.B(n_289),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1833),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1869),
.B(n_289),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1798),
.Y(n_1979)
);

BUFx3_ASAP7_75t_L g1980 ( 
.A(n_1823),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1869),
.B(n_290),
.Y(n_1981)
);

INVx1_ASAP7_75t_SL g1982 ( 
.A(n_1798),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1809),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1809),
.Y(n_1984)
);

INVx2_ASAP7_75t_SL g1985 ( 
.A(n_1823),
.Y(n_1985)
);

INVx1_ASAP7_75t_SL g1986 ( 
.A(n_1798),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1871),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1869),
.B(n_290),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1869),
.B(n_291),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1869),
.B(n_292),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1869),
.B(n_293),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1871),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1833),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1797),
.B(n_293),
.Y(n_1994)
);

CKINVDCx16_ASAP7_75t_R g1995 ( 
.A(n_1862),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1869),
.B(n_294),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1809),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1809),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_1823),
.Y(n_1999)
);

CKINVDCx16_ASAP7_75t_R g2000 ( 
.A(n_1862),
.Y(n_2000)
);

INVx1_ASAP7_75t_SL g2001 ( 
.A(n_1798),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1809),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1809),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1809),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1869),
.B(n_294),
.Y(n_2005)
);

INVxp67_ASAP7_75t_L g2006 ( 
.A(n_1875),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_1823),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1869),
.B(n_295),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1797),
.B(n_296),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1809),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1875),
.Y(n_2011)
);

INVx1_ASAP7_75t_SL g2012 ( 
.A(n_1798),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1809),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1797),
.B(n_297),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1797),
.B(n_298),
.Y(n_2015)
);

HB1xp67_ASAP7_75t_L g2016 ( 
.A(n_1871),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1833),
.Y(n_2017)
);

AOI211xp5_ASAP7_75t_L g2018 ( 
.A1(n_1936),
.A2(n_300),
.B(n_298),
.C(n_299),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1879),
.Y(n_2019)
);

AOI311xp33_ASAP7_75t_L g2020 ( 
.A1(n_1943),
.A2(n_1889),
.A3(n_1963),
.B(n_1896),
.C(n_1886),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1983),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1939),
.A2(n_1928),
.B(n_1942),
.Y(n_2022)
);

AOI222xp33_ASAP7_75t_L g2023 ( 
.A1(n_2006),
.A2(n_2011),
.B1(n_1946),
.B2(n_1960),
.C1(n_1952),
.C2(n_1949),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1984),
.Y(n_2024)
);

AOI21xp33_ASAP7_75t_SL g2025 ( 
.A1(n_1995),
.A2(n_299),
.B(n_300),
.Y(n_2025)
);

OAI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1909),
.A2(n_1974),
.B(n_1894),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1962),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1881),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1968),
.Y(n_2029)
);

INVx1_ASAP7_75t_SL g2030 ( 
.A(n_1878),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1970),
.B(n_2000),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1972),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1898),
.A2(n_1905),
.B1(n_1951),
.B2(n_1956),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_2017),
.B(n_301),
.Y(n_2034)
);

AOI21xp33_ASAP7_75t_L g2035 ( 
.A1(n_1962),
.A2(n_303),
.B(n_304),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1916),
.B(n_304),
.Y(n_2036)
);

OAI322xp33_ASAP7_75t_L g2037 ( 
.A1(n_1923),
.A2(n_311),
.A3(n_310),
.B1(n_308),
.B2(n_305),
.C1(n_306),
.C2(n_309),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1948),
.A2(n_305),
.B(n_306),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1980),
.B(n_308),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1899),
.B(n_309),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1987),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1938),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_2042)
);

NAND3xp33_ASAP7_75t_L g2043 ( 
.A(n_1917),
.B(n_1935),
.C(n_1959),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1908),
.B(n_312),
.Y(n_2044)
);

NAND3xp33_ASAP7_75t_L g2045 ( 
.A(n_1992),
.B(n_313),
.C(n_314),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1965),
.B(n_313),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1997),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1998),
.Y(n_2048)
);

INVxp67_ASAP7_75t_L g2049 ( 
.A(n_1932),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1977),
.B(n_314),
.Y(n_2050)
);

OAI21xp33_ASAP7_75t_L g2051 ( 
.A1(n_1945),
.A2(n_1934),
.B(n_1947),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1993),
.A2(n_317),
.B1(n_315),
.B2(n_316),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1929),
.B(n_315),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2002),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_2016),
.Y(n_2055)
);

NOR2x1_ASAP7_75t_L g2056 ( 
.A(n_1907),
.B(n_316),
.Y(n_2056)
);

INVxp67_ASAP7_75t_SL g2057 ( 
.A(n_1884),
.Y(n_2057)
);

OAI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1957),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_1931),
.B(n_318),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2003),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1950),
.A2(n_320),
.B(n_464),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1915),
.B(n_467),
.Y(n_2062)
);

AOI222xp33_ASAP7_75t_L g2063 ( 
.A1(n_1944),
.A2(n_470),
.B1(n_472),
.B2(n_468),
.C1(n_469),
.C2(n_471),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2004),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2010),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2013),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1910),
.Y(n_2067)
);

OAI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_1941),
.A2(n_474),
.B(n_475),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_SL g2069 ( 
.A1(n_1903),
.A2(n_1882),
.B(n_1955),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1937),
.A2(n_479),
.B1(n_476),
.B2(n_477),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1895),
.B(n_480),
.Y(n_2071)
);

INVxp33_ASAP7_75t_L g2072 ( 
.A(n_1937),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1897),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1901),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_1921),
.Y(n_2075)
);

OAI21xp33_ASAP7_75t_SL g2076 ( 
.A1(n_1890),
.A2(n_486),
.B(n_487),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_1887),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1927),
.Y(n_2078)
);

AOI322xp5_ASAP7_75t_L g2079 ( 
.A1(n_1953),
.A2(n_492),
.A3(n_493),
.B1(n_494),
.B2(n_495),
.C1(n_496),
.C2(n_498),
.Y(n_2079)
);

AOI22xp33_ASAP7_75t_L g2080 ( 
.A1(n_1961),
.A2(n_501),
.B1(n_499),
.B2(n_500),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1966),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1880),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_1900),
.B(n_503),
.Y(n_2083)
);

AND4x1_ASAP7_75t_L g2084 ( 
.A(n_1883),
.B(n_507),
.C(n_504),
.D(n_505),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1969),
.B(n_511),
.Y(n_2085)
);

INVxp67_ASAP7_75t_L g2086 ( 
.A(n_1958),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1967),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1978),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1979),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1989),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1991),
.Y(n_2091)
);

AOI211xp5_ASAP7_75t_SL g2092 ( 
.A1(n_1891),
.A2(n_522),
.B(n_519),
.C(n_520),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_1982),
.A2(n_2001),
.B1(n_2012),
.B2(n_1986),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1933),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2005),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1971),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1912),
.B(n_523),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_1919),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1985),
.B(n_526),
.Y(n_2099)
);

OAI21xp5_ASAP7_75t_SL g2100 ( 
.A1(n_1911),
.A2(n_528),
.B(n_530),
.Y(n_2100)
);

O2A1O1Ixp33_ASAP7_75t_L g2101 ( 
.A1(n_1926),
.A2(n_534),
.B(n_532),
.C(n_533),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_1930),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1907),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1981),
.Y(n_2104)
);

HB1xp67_ASAP7_75t_L g2105 ( 
.A(n_1954),
.Y(n_2105)
);

INVx1_ASAP7_75t_SL g2106 ( 
.A(n_1924),
.Y(n_2106)
);

XOR2x2_ASAP7_75t_L g2107 ( 
.A(n_1975),
.B(n_535),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1988),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1906),
.Y(n_2109)
);

NOR2xp67_ASAP7_75t_L g2110 ( 
.A(n_1999),
.B(n_537),
.Y(n_2110)
);

AOI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_1902),
.A2(n_1893),
.B1(n_1940),
.B2(n_1913),
.C(n_1920),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1990),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2007),
.B(n_539),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_1996),
.B(n_544),
.Y(n_2114)
);

INVxp67_ASAP7_75t_SL g2115 ( 
.A(n_2031),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2075),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2094),
.B(n_1918),
.Y(n_2117)
);

AOI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_2022),
.A2(n_2008),
.B(n_1925),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_2028),
.B(n_1892),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2081),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2077),
.B(n_1922),
.Y(n_2121)
);

INVxp67_ASAP7_75t_L g2122 ( 
.A(n_2093),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2098),
.B(n_1888),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_L g2124 ( 
.A(n_2030),
.B(n_1914),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_2072),
.B(n_1885),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2089),
.B(n_1964),
.Y(n_2126)
);

INVx2_ASAP7_75t_SL g2127 ( 
.A(n_2032),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2057),
.B(n_1973),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2036),
.Y(n_2129)
);

NAND2x1_ASAP7_75t_L g2130 ( 
.A(n_2029),
.B(n_1904),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2041),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2102),
.B(n_1976),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_2044),
.Y(n_2133)
);

NAND2x1_ASAP7_75t_L g2134 ( 
.A(n_2082),
.B(n_1994),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_2087),
.B(n_2009),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_2049),
.B(n_2014),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2106),
.B(n_2015),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2088),
.B(n_654),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2090),
.B(n_545),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2096),
.B(n_546),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_2091),
.B(n_2095),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2055),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2104),
.B(n_547),
.Y(n_2143)
);

AND2x4_ASAP7_75t_SL g2144 ( 
.A(n_2046),
.B(n_2050),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_2086),
.Y(n_2145)
);

NAND2xp33_ASAP7_75t_L g2146 ( 
.A(n_2020),
.B(n_548),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_2069),
.B(n_549),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_2034),
.B(n_550),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2034),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2059),
.B(n_551),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2108),
.B(n_2112),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_2040),
.B(n_552),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2043),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2051),
.B(n_556),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2038),
.B(n_557),
.Y(n_2155)
);

NOR3xp33_ASAP7_75t_L g2156 ( 
.A(n_2025),
.B(n_2037),
.C(n_2035),
.Y(n_2156)
);

NOR2x1_ASAP7_75t_L g2157 ( 
.A(n_2056),
.B(n_558),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2111),
.B(n_559),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2105),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2023),
.B(n_560),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2103),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2076),
.A2(n_565),
.B1(n_561),
.B2(n_564),
.Y(n_2162)
);

NOR2x1_ASAP7_75t_L g2163 ( 
.A(n_2045),
.B(n_567),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_2053),
.B(n_2039),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_2058),
.B(n_568),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2026),
.B(n_2071),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_2073),
.B(n_569),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2074),
.B(n_570),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2019),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2067),
.B(n_2021),
.Y(n_2170)
);

AND2x2_ASAP7_75t_SL g2171 ( 
.A(n_2078),
.B(n_573),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2027),
.B(n_653),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2141),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2151),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2170),
.Y(n_2175)
);

INVx1_ASAP7_75t_SL g2176 ( 
.A(n_2132),
.Y(n_2176)
);

CKINVDCx20_ASAP7_75t_R g2177 ( 
.A(n_2144),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2131),
.Y(n_2178)
);

CKINVDCx6p67_ASAP7_75t_R g2179 ( 
.A(n_2121),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2142),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2159),
.Y(n_2181)
);

INVxp67_ASAP7_75t_L g2182 ( 
.A(n_2145),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2169),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2116),
.Y(n_2184)
);

BUFx2_ASAP7_75t_L g2185 ( 
.A(n_2115),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2120),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2135),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2129),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2161),
.Y(n_2189)
);

INVxp33_ASAP7_75t_SL g2190 ( 
.A(n_2124),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2117),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2137),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2128),
.Y(n_2193)
);

INVx1_ASAP7_75t_SL g2194 ( 
.A(n_2146),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2119),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2123),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2119),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_2122),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2126),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2133),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2156),
.B(n_2164),
.Y(n_2201)
);

INVx1_ASAP7_75t_SL g2202 ( 
.A(n_2167),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2149),
.Y(n_2203)
);

CKINVDCx20_ASAP7_75t_R g2204 ( 
.A(n_2127),
.Y(n_2204)
);

NAND4xp75_ASAP7_75t_L g2205 ( 
.A(n_2201),
.B(n_2157),
.C(n_2163),
.D(n_2160),
.Y(n_2205)
);

AOI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_2194),
.A2(n_2033),
.B1(n_2166),
.B2(n_2147),
.C(n_2018),
.Y(n_2206)
);

AND2x2_ASAP7_75t_SL g2207 ( 
.A(n_2185),
.B(n_2136),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_2177),
.B(n_2125),
.Y(n_2208)
);

NAND3xp33_ASAP7_75t_L g2209 ( 
.A(n_2198),
.B(n_2042),
.C(n_2153),
.Y(n_2209)
);

AOI221xp5_ASAP7_75t_L g2210 ( 
.A1(n_2194),
.A2(n_2186),
.B1(n_2202),
.B2(n_2196),
.C(n_2173),
.Y(n_2210)
);

NAND3xp33_ASAP7_75t_L g2211 ( 
.A(n_2182),
.B(n_2063),
.C(n_2158),
.Y(n_2211)
);

OAI21xp33_ASAP7_75t_L g2212 ( 
.A1(n_2190),
.A2(n_2118),
.B(n_2134),
.Y(n_2212)
);

AOI311xp33_ASAP7_75t_L g2213 ( 
.A1(n_2191),
.A2(n_2048),
.A3(n_2054),
.B(n_2047),
.C(n_2024),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_2204),
.B(n_2061),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2195),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2176),
.B(n_2130),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2193),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2187),
.Y(n_2218)
);

AOI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_2174),
.A2(n_2155),
.B(n_2172),
.Y(n_2219)
);

NOR2xp67_ASAP7_75t_SL g2220 ( 
.A(n_2197),
.B(n_2100),
.Y(n_2220)
);

NAND4xp25_ASAP7_75t_SL g2221 ( 
.A(n_2199),
.B(n_2162),
.C(n_2060),
.D(n_2065),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2179),
.B(n_2064),
.Y(n_2222)
);

AOI22xp33_ASAP7_75t_SL g2223 ( 
.A1(n_2211),
.A2(n_2175),
.B1(n_2203),
.B2(n_2171),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2207),
.B(n_2200),
.Y(n_2224)
);

NAND4xp25_ASAP7_75t_L g2225 ( 
.A(n_2210),
.B(n_2192),
.C(n_2180),
.D(n_2178),
.Y(n_2225)
);

OAI21xp33_ASAP7_75t_L g2226 ( 
.A1(n_2212),
.A2(n_2184),
.B(n_2181),
.Y(n_2226)
);

NOR4xp25_ASAP7_75t_L g2227 ( 
.A(n_2213),
.B(n_2188),
.C(n_2183),
.D(n_2189),
.Y(n_2227)
);

AOI21xp33_ASAP7_75t_SL g2228 ( 
.A1(n_2214),
.A2(n_2052),
.B(n_2066),
.Y(n_2228)
);

NAND4xp75_ASAP7_75t_L g2229 ( 
.A(n_2216),
.B(n_2154),
.C(n_2110),
.D(n_2165),
.Y(n_2229)
);

OA22x2_ASAP7_75t_L g2230 ( 
.A1(n_2208),
.A2(n_2068),
.B1(n_2109),
.B2(n_2138),
.Y(n_2230)
);

OAI211xp5_ASAP7_75t_SL g2231 ( 
.A1(n_2206),
.A2(n_2092),
.B(n_2101),
.C(n_2079),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2228),
.B(n_2208),
.Y(n_2232)
);

NOR3xp33_ASAP7_75t_L g2233 ( 
.A(n_2224),
.B(n_2205),
.C(n_2221),
.Y(n_2233)
);

NOR2x1_ASAP7_75t_L g2234 ( 
.A(n_2225),
.B(n_2222),
.Y(n_2234)
);

OAI22x1_ASAP7_75t_L g2235 ( 
.A1(n_2227),
.A2(n_2215),
.B1(n_2218),
.B2(n_2217),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2223),
.B(n_2219),
.Y(n_2236)
);

NOR2x1_ASAP7_75t_L g2237 ( 
.A(n_2226),
.B(n_2209),
.Y(n_2237)
);

XNOR2x1_ASAP7_75t_L g2238 ( 
.A(n_2229),
.B(n_2107),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2230),
.B(n_2220),
.Y(n_2239)
);

NAND2xp33_ASAP7_75t_SL g2240 ( 
.A(n_2235),
.B(n_2085),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_R g2241 ( 
.A(n_2232),
.B(n_2083),
.Y(n_2241)
);

XNOR2xp5_ASAP7_75t_L g2242 ( 
.A(n_2238),
.B(n_2084),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_2233),
.B(n_2231),
.Y(n_2243)
);

NAND3xp33_ASAP7_75t_L g2244 ( 
.A(n_2234),
.B(n_2152),
.C(n_2150),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2243),
.Y(n_2245)
);

NAND2x1_ASAP7_75t_SL g2246 ( 
.A(n_2240),
.B(n_2237),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2245),
.Y(n_2247)
);

INVxp67_ASAP7_75t_SL g2248 ( 
.A(n_2247),
.Y(n_2248)
);

AOI22xp33_ASAP7_75t_L g2249 ( 
.A1(n_2248),
.A2(n_2239),
.B1(n_2244),
.B2(n_2236),
.Y(n_2249)
);

AOI22xp33_ASAP7_75t_L g2250 ( 
.A1(n_2248),
.A2(n_2241),
.B1(n_2242),
.B2(n_2097),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2249),
.B(n_2250),
.Y(n_2251)
);

OAI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_2249),
.A2(n_2246),
.B1(n_2139),
.B2(n_2114),
.Y(n_2252)
);

OAI21xp5_ASAP7_75t_SL g2253 ( 
.A1(n_2251),
.A2(n_2252),
.B(n_2113),
.Y(n_2253)
);

OAI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2252),
.A2(n_2143),
.B(n_2140),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2253),
.Y(n_2255)
);

HB1xp67_ASAP7_75t_L g2256 ( 
.A(n_2254),
.Y(n_2256)
);

OAI221xp5_ASAP7_75t_R g2257 ( 
.A1(n_2256),
.A2(n_2080),
.B1(n_2070),
.B2(n_2168),
.C(n_2099),
.Y(n_2257)
);

AOI211xp5_ASAP7_75t_L g2258 ( 
.A1(n_2257),
.A2(n_2255),
.B(n_2148),
.C(n_2062),
.Y(n_2258)
);


endmodule