module real_jpeg_33261_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_0),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g300 ( 
.A(n_0),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_L g53 ( 
.A(n_1),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_1),
.B(n_244),
.Y(n_243)
);

NAND2x1_ASAP7_75t_L g258 ( 
.A(n_1),
.B(n_259),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_R g264 ( 
.A(n_1),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_1),
.B(n_309),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g328 ( 
.A(n_1),
.B(n_146),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_1),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_1),
.B(n_256),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_2),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_2),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_2),
.B(n_115),
.Y(n_114)
);

NAND2x1p5_ASAP7_75t_L g179 ( 
.A(n_2),
.B(n_98),
.Y(n_179)
);

NAND2x1_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_3),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_3),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_3),
.B(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_3),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_3),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_3),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_4),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_4),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_4),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_4),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_4),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_4),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_4),
.B(n_356),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_5),
.Y(n_168)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_7),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_7),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_7),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_37),
.Y(n_44)
);

NAND2x1_ASAP7_75t_L g60 ( 
.A(n_8),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_8),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_8),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_8),
.B(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_10),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_29),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_11),
.B(n_51),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_11),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_11),
.B(n_26),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_11),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_12),
.B(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_12),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_12),
.B(n_256),
.Y(n_263)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_13),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_14),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_15),
.B(n_67),
.Y(n_66)
);

NAND2x1_ASAP7_75t_L g97 ( 
.A(n_15),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_15),
.B(n_112),
.Y(n_111)
);

AND2x4_ASAP7_75t_SL g166 ( 
.A(n_15),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_15),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_15),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_15),
.B(n_283),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_15),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_220),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_217),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_182),
.Y(n_19)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_20),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_106),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_69),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_46),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.C(n_31),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_25),
.A2(n_28),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_25),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_25),
.A2(n_102),
.B1(n_194),
.B2(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_28),
.A2(n_103),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_28),
.B(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_28),
.B(n_282),
.Y(n_306)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_30),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_31),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_33),
.Y(n_200)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_33),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_40),
.Y(n_246)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_43),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_59),
.C(n_64),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2x1_ASAP7_75t_L g137 ( 
.A(n_48),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.C(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_53),
.B(n_56),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_56),
.B(n_175),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g286 ( 
.A1(n_56),
.A2(n_174),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_56),
.B(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_60),
.A2(n_66),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_62),
.Y(n_311)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_68),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_85),
.C(n_100),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_70),
.A2(n_71),
.B1(n_85),
.B2(n_86),
.Y(n_213)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

OAI22x1_ASAP7_75t_L g170 ( 
.A1(n_72),
.A2(n_82),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2x1_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_78),
.B(n_82),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_80),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.C(n_97),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2x2_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_89),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_90),
.Y(n_358)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_100),
.Y(n_212)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_102),
.B(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_161),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_136),
.C(n_141),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_109),
.B(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_123),
.C(n_133),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_110),
.B(n_133),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.C(n_118),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_111),
.B(n_163),
.Y(n_267)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_117),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_118),
.B(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_123),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.C(n_129),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_124),
.B(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_129),
.Y(n_192)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_131),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_132),
.Y(n_241)
);

BUFx2_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_137),
.B(n_142),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.C(n_155),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_143),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_155),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_159),
.Y(n_265)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2x2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_169),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_175),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_210),
.C(n_214),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_183),
.B(n_400),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.C(n_207),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_184),
.B(n_208),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

XOR2x2_ASAP7_75t_SL g395 ( 
.A(n_190),
.B(n_396),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_196),
.Y(n_190)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_193),
.B(n_197),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.C(n_204),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_204),
.B1(n_205),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_211),
.B(n_215),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_382),
.B(n_401),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_289),
.B(n_380),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_268),
.Y(n_223)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_224),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_250),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_247),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_226),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.C(n_233),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_227),
.B(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.C(n_242),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_234),
.A2(n_235),
.B1(n_242),
.B2(n_243),
.Y(n_372)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_239),
.B(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_247),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_250),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_266),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_262),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_252),
.B(n_262),
.C(n_266),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.C(n_258),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_254),
.B(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_258),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_269),
.B(n_381),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.C(n_276),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_270),
.B(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_276),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.C(n_286),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_277),
.A2(n_278),
.B1(n_286),
.B2(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_280),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_286),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_374),
.B(n_379),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_363),
.B(n_373),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_333),
.B(n_362),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_325),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_307),
.B1(n_323),
.B2(n_324),
.Y(n_293)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

AOI221xp5_ASAP7_75t_L g362 ( 
.A1(n_294),
.A2(n_307),
.B1(n_323),
.B2(n_324),
.C(n_325),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_305),
.B2(n_306),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_295),
.B(n_306),
.C(n_324),
.Y(n_364)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_301),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_301),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_300),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_312),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_308),
.B(n_313),
.C(n_317),
.Y(n_370)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_317),
.B1(n_321),
.B2(n_322),
.Y(n_312)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.C(n_329),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_326),
.A2(n_327),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_328),
.A2(n_329),
.B1(n_330),
.B2(n_347),
.Y(n_346)
);

CKINVDCx12_ASAP7_75t_R g347 ( 
.A(n_328),
.Y(n_347)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_348),
.B(n_361),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_344),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_344),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_341),
.Y(n_350)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_354),
.B(n_360),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_351),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.Y(n_354)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_365),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_369),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_370),
.C(n_371),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_378),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_SL g379 ( 
.A(n_375),
.B(n_378),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR2x1_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_397),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_389),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_389),
.Y(n_403)
);

MAJx2_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.C(n_388),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_395),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_392),
.C(n_395),
.Y(n_398)
);

XNOR2x2_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_397),
.A2(n_403),
.B(n_404),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_399),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);


endmodule