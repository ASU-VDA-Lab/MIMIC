module fake_jpeg_18531_n_311 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_10),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_16),
.B1(n_19),
.B2(n_13),
.Y(n_38)
);

AO22x1_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_34),
.B1(n_25),
.B2(n_28),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_31),
.B1(n_16),
.B2(n_32),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_39),
.B1(n_35),
.B2(n_43),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_31),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_34),
.B1(n_25),
.B2(n_33),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_52),
.B1(n_39),
.B2(n_35),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_36),
.B1(n_28),
.B2(n_27),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_30),
.B1(n_16),
.B2(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_16),
.B1(n_24),
.B2(n_28),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_19),
.B1(n_22),
.B2(n_13),
.Y(n_78)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_59),
.Y(n_77)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_68),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_38),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_33),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_43),
.B1(n_19),
.B2(n_14),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_13),
.B(n_12),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_48),
.B(n_61),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_60),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_19),
.B1(n_15),
.B2(n_12),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_58),
.B1(n_55),
.B2(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_48),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_73),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_93),
.B1(n_73),
.B2(n_76),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_86),
.B1(n_88),
.B2(n_74),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_66),
.C(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_84),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_67),
.B1(n_70),
.B2(n_65),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_72),
.B(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_95),
.Y(n_113)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_48),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_46),
.C(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_98),
.Y(n_119)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_46),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_67),
.B1(n_69),
.B2(n_75),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_112),
.B1(n_97),
.B2(n_81),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_102),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_110),
.B(n_116),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_72),
.B(n_77),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_0),
.B(n_1),
.Y(n_153)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_78),
.B(n_64),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_114),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_47),
.B1(n_50),
.B2(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_123),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_73),
.B1(n_63),
.B2(n_76),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_85),
.B(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_22),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_118),
.B(n_22),
.Y(n_129)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_27),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_133),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_83),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_135),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_129),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_110),
.B(n_115),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_90),
.B(n_88),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_136),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_83),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_123),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_86),
.A3(n_93),
.B1(n_96),
.B2(n_99),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_26),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_139),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_100),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_116),
.B1(n_36),
.B2(n_27),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_148),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_81),
.B1(n_97),
.B2(n_92),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_121),
.B1(n_109),
.B2(n_112),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_80),
.B(n_62),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_153),
.B(n_116),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_63),
.Y(n_147)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_106),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_81),
.B1(n_92),
.B2(n_29),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_106),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_15),
.B1(n_21),
.B2(n_49),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_116),
.B(n_15),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_119),
.C(n_117),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_164),
.C(n_170),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_117),
.B1(n_113),
.B2(n_101),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_182),
.B1(n_160),
.B2(n_169),
.Y(n_205)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_134),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_171),
.B1(n_173),
.B2(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_181),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_119),
.C(n_115),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_111),
.C(n_116),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_172),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_140),
.B1(n_142),
.B2(n_131),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_23),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_29),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_178),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_183),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_132),
.A2(n_130),
.B(n_141),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_171),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_194),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_142),
.C(n_128),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_161),
.C(n_174),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_129),
.Y(n_195)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_133),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_181),
.B(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_124),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_167),
.B(n_163),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_165),
.B(n_148),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_203),
.B(n_7),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_18),
.B1(n_23),
.B2(n_11),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_138),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_157),
.B1(n_169),
.B2(n_173),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_214),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_172),
.B1(n_159),
.B2(n_178),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_162),
.C(n_125),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_201),
.C(n_185),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_136),
.B1(n_151),
.B2(n_178),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_151),
.B(n_153),
.C(n_180),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_154),
.B1(n_26),
.B2(n_18),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_229),
.B1(n_7),
.B2(n_10),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_190),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_7),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_192),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_193),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_245),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_201),
.B(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_238),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_202),
.C(n_191),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_184),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_241),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_188),
.C(n_186),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_244),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_186),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_20),
.C(n_18),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_21),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_222),
.B1(n_225),
.B2(n_224),
.Y(n_252)
);

OAI321xp33_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_220),
.A3(n_230),
.B1(n_219),
.B2(n_214),
.C(n_213),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_228),
.B(n_216),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_264),
.B1(n_245),
.B2(n_243),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_6),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_235),
.A2(n_221),
.B(n_218),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_255),
.A2(n_0),
.B(n_1),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_6),
.B1(n_10),
.B2(n_8),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_232),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_234),
.A2(n_220),
.B1(n_249),
.B2(n_236),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_240),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_220),
.B(n_21),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_265),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_268),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_257),
.B(n_276),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_11),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_11),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_271),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_270),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_11),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_273),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_18),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_20),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_275),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_20),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_6),
.C(n_1),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_0),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_3),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_262),
.B1(n_20),
.B2(n_3),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_2),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_290),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_20),
.C(n_3),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_280),
.C(n_281),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_2),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_292),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_277),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_296),
.B(n_297),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_3),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_4),
.Y(n_298)
);

NAND4xp25_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_299),
.C(n_284),
.D(n_289),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_4),
.B(n_5),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_291),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_304),
.A2(n_305),
.B(n_293),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_287),
.B(n_295),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_307),
.B(n_302),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_301),
.B(n_4),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_5),
.B(n_301),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_5),
.Y(n_311)
);


endmodule