module fake_jpeg_25622_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx16f_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

INVx8_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_2),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_15),
.B(n_16),
.Y(n_18)
);

AO22x2_ASAP7_75t_L g16 ( 
.A1(n_9),
.A2(n_6),
.B1(n_5),
.B2(n_12),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_18),
.B(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_17),
.Y(n_20)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_21),
.B(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_16),
.B1(n_20),
.B2(n_12),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

AO221x1_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_16),
.B1(n_6),
.B2(n_14),
.C(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_14),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_22),
.B(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_29),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_3),
.B(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_7),
.Y(n_33)
);


endmodule