module fake_jpeg_1821_n_195 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_12),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_66),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_70),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_73),
.Y(n_77)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_57),
.Y(n_74)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_72),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_62),
.B1(n_63),
.B2(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_81),
.B1(n_83),
.B2(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_84),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_SL g80 ( 
.A(n_66),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_68),
.B1(n_63),
.B2(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_50),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_70),
.B1(n_52),
.B2(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_100),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_102),
.Y(n_110)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_68),
.B1(n_83),
.B2(n_71),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_116),
.B1(n_17),
.B2(n_42),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_60),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_114),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_82),
.B(n_58),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_115),
.B(n_1),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_54),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_59),
.B(n_55),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_53),
.B1(n_67),
.B2(n_70),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_20),
.C(n_45),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_43),
.C(n_41),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_0),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_18),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_65),
.B(n_2),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_6),
.B(n_9),
.Y(n_141)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_131),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_140),
.B1(n_141),
.B2(n_105),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_129),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_1),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_3),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_5),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_140)
);

NAND2x1_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_120),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_158),
.B(n_33),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_105),
.B1(n_119),
.B2(n_11),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_117),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_128),
.C(n_35),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_28),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_154),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_27),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_105),
.B(n_10),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_9),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_159),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_10),
.B(n_12),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_131),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_163),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_164),
.B1(n_171),
.B2(n_144),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_13),
.B1(n_15),
.B2(n_22),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_23),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_167),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_143),
.B(n_158),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_40),
.B1(n_36),
.B2(n_37),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_174),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_168),
.B(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

AOI321xp33_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_150),
.A3(n_148),
.B1(n_152),
.B2(n_154),
.C(n_156),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_163),
.B1(n_175),
.B2(n_178),
.Y(n_182)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_172),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_184),
.A2(n_162),
.B1(n_165),
.B2(n_179),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_SL g189 ( 
.A(n_188),
.B(n_185),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_186),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_190),
.B(n_183),
.Y(n_191)
);

AOI21x1_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_187),
.B(n_181),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_184),
.B(n_38),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_34),
.Y(n_195)
);


endmodule