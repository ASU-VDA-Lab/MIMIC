module fake_jpeg_82_n_64 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_19),
.B(n_21),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_20),
.B1(n_14),
.B2(n_17),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_22),
.B(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AO22x1_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_19),
.B1(n_22),
.B2(n_18),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_38),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_12),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_50),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_38),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_44),
.C(n_40),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_44),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_12),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_31),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_41),
.B(n_39),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_47),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_52),
.Y(n_58)
);

MAJx2_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_11),
.C(n_35),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_56),
.B(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_61),
.B(n_4),
.Y(n_63)
);

AOI322xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_2),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_24),
.C2(n_54),
.Y(n_64)
);


endmodule