module fake_jpeg_22835_n_313 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_24),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_32),
.Y(n_56)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_57),
.Y(n_78)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_19),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_81),
.Y(n_90)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_37),
.B1(n_21),
.B2(n_26),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_37),
.B1(n_58),
.B2(n_72),
.Y(n_86)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_72),
.Y(n_92)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g93 ( 
.A(n_74),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_19),
.B1(n_33),
.B2(n_31),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_38),
.B1(n_49),
.B2(n_44),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_19),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_71),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_102),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_80),
.B1(n_63),
.B2(n_40),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_26),
.B1(n_25),
.B2(n_46),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_45),
.B1(n_41),
.B2(n_26),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_103),
.B1(n_77),
.B2(n_38),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_19),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_62),
.B(n_76),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_43),
.A3(n_50),
.B1(n_25),
.B2(n_26),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_25),
.B1(n_45),
.B2(n_29),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_55),
.C(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_64),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_33),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_76),
.B(n_66),
.C(n_40),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_106),
.A2(n_117),
.B(n_120),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_80),
.B1(n_59),
.B2(n_78),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_78),
.B1(n_67),
.B2(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_122),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_84),
.A2(n_16),
.B(n_14),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_94),
.Y(n_136)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_33),
.B(n_31),
.C(n_22),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_16),
.B1(n_14),
.B2(n_62),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_92),
.B1(n_91),
.B2(n_78),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_127),
.Y(n_134)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_130),
.Y(n_149)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_145),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_90),
.B(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_138),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_154),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_99),
.C(n_83),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_143),
.C(n_155),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_139),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_85),
.C(n_96),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_150),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_115),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_153),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_89),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_122),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_85),
.C(n_92),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_172),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_119),
.B1(n_128),
.B2(n_125),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_133),
.B1(n_140),
.B2(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_161),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_125),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_143),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_108),
.C(n_97),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_120),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_113),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_179),
.Y(n_201)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_148),
.B(n_126),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_143),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_183),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_177),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_185),
.B(n_161),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_137),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_191),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_141),
.A3(n_136),
.B1(n_138),
.B2(n_135),
.C1(n_95),
.C2(n_140),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_190),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_131),
.Y(n_191)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_196),
.C(n_197),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_106),
.B(n_144),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_195),
.B1(n_171),
.B2(n_178),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_106),
.B1(n_144),
.B2(n_124),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_151),
.C(n_118),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_129),
.C(n_127),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_180),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_124),
.C(n_88),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_167),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_175),
.A2(n_101),
.B1(n_91),
.B2(n_130),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_203),
.A2(n_156),
.B1(n_173),
.B2(n_160),
.Y(n_208)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_208),
.A2(n_222),
.B1(n_195),
.B2(n_187),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_159),
.B(n_174),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_209),
.A2(n_21),
.B(n_23),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_213),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_216),
.B1(n_204),
.B2(n_200),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_188),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_201),
.Y(n_214)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_226),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_163),
.B1(n_162),
.B2(n_166),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_109),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_223),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_183),
.B(n_163),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_130),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_184),
.C(n_109),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_191),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_231),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_182),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_235),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_SL g234 ( 
.A(n_226),
.B(n_197),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_240),
.C(n_212),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_196),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_194),
.B1(n_200),
.B2(n_192),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_209),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_242),
.B1(n_245),
.B2(n_16),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_202),
.B1(n_203),
.B2(n_193),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_158),
.C(n_101),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_244),
.C(n_208),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_109),
.C(n_75),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_91),
.B1(n_61),
.B2(n_14),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_246),
.A2(n_221),
.B(n_23),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_257),
.B1(n_18),
.B2(n_27),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_104),
.Y(n_266)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_18),
.B(n_24),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_220),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_29),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_254),
.A2(n_238),
.B1(n_235),
.B2(n_230),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_221),
.C(n_74),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_256),
.C(n_259),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_104),
.C(n_21),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_229),
.C(n_233),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_246),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_262),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_236),
.B(n_17),
.Y(n_262)
);

OAI322xp33_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_29),
.A3(n_18),
.B1(n_23),
.B2(n_21),
.C1(n_17),
.C2(n_22),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_264),
.A2(n_28),
.B(n_27),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_276),
.C(n_277),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_274),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_270),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_251),
.B1(n_28),
.B2(n_13),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_249),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_250),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_15),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_15),
.C(n_27),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_22),
.C(n_28),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_280),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_260),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_277),
.C(n_1),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_285),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_260),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_273),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_13),
.B(n_11),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_289),
.A2(n_278),
.B(n_269),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_11),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_0),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_292),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_297),
.C(n_282),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_280),
.B(n_0),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_0),
.B(n_1),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_1),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_0),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_299),
.A2(n_304),
.B1(n_293),
.B2(n_4),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_286),
.A3(n_287),
.B1(n_281),
.B2(n_279),
.C1(n_4),
.C2(n_5),
.Y(n_300)
);

A2O1A1O1Ixp25_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_301),
.B(n_3),
.C(n_6),
.D(n_7),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_298),
.A2(n_1),
.B(n_2),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_302),
.A2(n_3),
.B(n_5),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_306),
.A3(n_307),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_308),
.A2(n_303),
.B(n_7),
.Y(n_309)
);

AOI32xp33_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_6),
.B(n_8),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_10),
.Y(n_313)
);


endmodule