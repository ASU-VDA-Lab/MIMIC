module fake_jpeg_28465_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_34),
.B(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_59),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_20),
.B1(n_33),
.B2(n_30),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_50),
.B1(n_37),
.B2(n_5),
.Y(n_67)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_39),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_3),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_59),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_42),
.B1(n_4),
.B2(n_6),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_72),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_44),
.C(n_46),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_88),
.C(n_38),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_47),
.B(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_81),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_82),
.B1(n_87),
.B2(n_22),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_47),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_43),
.B(n_7),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_9),
.B(n_10),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_83),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_47),
.B1(n_38),
.B2(n_9),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_23),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_93),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_96),
.B(n_100),
.Y(n_105)
);

OAI22x1_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_35),
.B1(n_12),
.B2(n_17),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_11),
.C(n_18),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_99),
.C(n_88),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_88),
.C(n_76),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_19),
.B(n_21),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_107),
.C(n_96),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_24),
.C(n_25),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_110),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_92),
.C(n_90),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_99),
.B1(n_97),
.B2(n_94),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_111),
.B(n_106),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_105),
.C(n_103),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_26),
.C(n_27),
.Y(n_115)
);

HAxp5_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_28),
.CON(n_116),
.SN(n_116)
);


endmodule