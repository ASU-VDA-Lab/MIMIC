module fake_jpeg_20269_n_254 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_149;
wire n_35;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_24),
.B(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_47),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_24),
.B1(n_26),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_27),
.B1(n_32),
.B2(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_30),
.B1(n_34),
.B2(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_23),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_23),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_34),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_54),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_74),
.B1(n_50),
.B2(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_41),
.B1(n_42),
.B2(n_34),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_41),
.B1(n_42),
.B2(n_34),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_55),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_36),
.B(n_42),
.C(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_78),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_89),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_75),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_45),
.B1(n_46),
.B2(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_85),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_25),
.B1(n_38),
.B2(n_21),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_71),
.B1(n_68),
.B2(n_11),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_22),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_73),
.B(n_21),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_38),
.C(n_25),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_60),
.C(n_38),
.Y(n_94)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_74),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_84),
.B(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_106),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_97),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_108),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_72),
.C(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_11),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_60),
.C(n_70),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_60),
.B1(n_14),
.B2(n_68),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_15),
.B(n_12),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_71),
.B1(n_25),
.B2(n_68),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_112),
.A2(n_92),
.B1(n_85),
.B2(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_120),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_77),
.B(n_84),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_114),
.A2(n_116),
.B(n_117),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_126),
.B1(n_99),
.B2(n_105),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_89),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_84),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_136),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_92),
.B1(n_91),
.B2(n_81),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_0),
.B(n_1),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_133),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_14),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_10),
.Y(n_153)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_137),
.Y(n_146)
);

XOR2x1_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_15),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_139),
.B(n_151),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_106),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_145),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_98),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_94),
.B1(n_109),
.B2(n_108),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_161),
.B1(n_152),
.B2(n_158),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_100),
.B1(n_62),
.B2(n_2),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_157),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_162),
.B(n_120),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_10),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_156),
.B(n_132),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_62),
.B1(n_1),
.B2(n_2),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_15),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_138),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_38),
.C(n_51),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_117),
.C(n_114),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_62),
.B1(n_1),
.B2(n_3),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_118),
.A2(n_35),
.A3(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_168),
.C(n_149),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_116),
.C(n_127),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_130),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_177),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_133),
.B1(n_116),
.B2(n_137),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_180),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_121),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_181),
.B(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_144),
.B1(n_139),
.B2(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_192),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_143),
.B(n_124),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_188),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_143),
.B(n_147),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_145),
.C(n_160),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_168),
.C(n_176),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_197),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_162),
.B(n_147),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_206),
.C(n_197),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_163),
.C(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_205),
.Y(n_215)
);

OAI322xp33_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_155),
.A3(n_178),
.B1(n_169),
.B2(n_174),
.C1(n_165),
.C2(n_136),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_192),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_113),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_165),
.C(n_51),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_184),
.C(n_191),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_10),
.Y(n_207)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_35),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_212),
.B(n_220),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_202),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_217),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_198),
.B1(n_208),
.B2(n_182),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_35),
.B1(n_15),
.B2(n_56),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_188),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_195),
.C(n_190),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_51),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_187),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_200),
.B(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_214),
.B(n_222),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_226),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_16),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_43),
.C(n_38),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_227),
.C(n_43),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_217),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_239),
.B1(n_232),
.B2(n_16),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_0),
.B(n_4),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_0),
.B(n_4),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_35),
.B(n_43),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_235),
.A2(n_19),
.B(n_20),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_35),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_237),
.A2(n_238),
.B1(n_12),
.B2(n_6),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_230),
.A3(n_20),
.B1(n_19),
.B2(n_17),
.C1(n_16),
.C2(n_12),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_244),
.B(n_239),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_5),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_19),
.A3(n_20),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_5),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_248),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_251),
.A2(n_249),
.B1(n_245),
.B2(n_8),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_8),
.C(n_6),
.Y(n_253)
);

OAI311xp33_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_6),
.A3(n_7),
.B1(n_178),
.C1(n_251),
.Y(n_254)
);


endmodule