module fake_jpeg_30229_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx6f_ASAP7_75t_SL g72 ( 
.A(n_7),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_95),
.Y(n_102)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_57),
.B1(n_63),
.B2(n_71),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_93),
.B1(n_55),
.B2(n_58),
.Y(n_101)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_68),
.B1(n_71),
.B2(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_52),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_51),
.B1(n_58),
.B2(n_55),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_57),
.B1(n_63),
.B2(n_51),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_98),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_103),
.B1(n_91),
.B2(n_112),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_103),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_79),
.B1(n_65),
.B2(n_66),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_67),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_70),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_65),
.B(n_53),
.C(n_70),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_0),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_4),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_122),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_126),
.B1(n_127),
.B2(n_13),
.Y(n_147)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_69),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_114),
.A2(n_92),
.B1(n_61),
.B2(n_53),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_92),
.B1(n_53),
.B2(n_70),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_134),
.B(n_135),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_25),
.B(n_48),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_6),
.B(n_9),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_136),
.A2(n_135),
.B(n_134),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_49),
.B(n_26),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_139),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_141),
.B1(n_147),
.B2(n_23),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_11),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_145),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_29),
.B1(n_46),
.B2(n_45),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_12),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_144),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_115),
.C(n_117),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_131),
.B(n_16),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_16),
.Y(n_152)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_153),
.B(n_18),
.C(n_20),
.D(n_21),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_32),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_124),
.B(n_121),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_151),
.B(n_147),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_160),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_161),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_137),
.C(n_150),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_145),
.C(n_153),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_154),
.B(n_137),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_162),
.B1(n_167),
.B2(n_146),
.Y(n_169)
);

OAI221xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_165),
.B1(n_162),
.B2(n_141),
.C(n_164),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_47),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_24),
.C(n_27),
.Y(n_172)
);

AOI321xp33_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_34),
.A3(n_36),
.B1(n_37),
.B2(n_40),
.C(n_41),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_42),
.Y(n_174)
);


endmodule