module real_jpeg_14256_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_1),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_1),
.A2(n_60),
.B1(n_63),
.B2(n_71),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_46),
.B1(n_48),
.B2(n_71),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_1),
.A2(n_34),
.B1(n_41),
.B2(n_71),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_3),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_3),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_3),
.A2(n_65),
.B(n_201),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g226 ( 
.A1(n_3),
.A2(n_46),
.B1(n_48),
.B2(n_192),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_3),
.A2(n_48),
.B(n_51),
.C(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_3),
.B(n_84),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_3),
.B(n_38),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_3),
.B(n_56),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_3),
.A2(n_63),
.B(n_78),
.C(n_263),
.Y(n_262)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_5),
.A2(n_60),
.B1(n_63),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_5),
.A2(n_46),
.B1(n_48),
.B2(n_77),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_5),
.A2(n_34),
.B1(n_41),
.B2(n_77),
.Y(n_182)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_7),
.A2(n_60),
.B1(n_63),
.B2(n_69),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_7),
.A2(n_46),
.B1(n_48),
.B2(n_69),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_7),
.A2(n_34),
.B1(n_41),
.B2(n_69),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_8),
.A2(n_45),
.B1(n_60),
.B2(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_8),
.A2(n_45),
.B1(n_65),
.B2(n_66),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_8),
.A2(n_34),
.B1(n_41),
.B2(n_45),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_9),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_9),
.A2(n_40),
.B1(n_60),
.B2(n_63),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_9),
.A2(n_40),
.B1(n_65),
.B2(n_66),
.Y(n_329)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_11),
.A2(n_60),
.B1(n_63),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_11),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_174),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_11),
.A2(n_46),
.B1(n_48),
.B2(n_174),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_11),
.A2(n_34),
.B1(n_41),
.B2(n_174),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_12),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_12),
.A2(n_60),
.B1(n_63),
.B2(n_161),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_12),
.A2(n_46),
.B1(n_48),
.B2(n_161),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_12),
.A2(n_34),
.B1(n_41),
.B2(n_161),
.Y(n_241)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_14),
.Y(n_341)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_17),
.A2(n_65),
.B1(n_66),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_17),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_17),
.A2(n_46),
.B1(n_48),
.B2(n_125),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_17),
.A2(n_60),
.B1(n_63),
.B2(n_125),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_17),
.A2(n_34),
.B1(n_41),
.B2(n_125),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_18),
.A2(n_46),
.B1(n_48),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_18),
.A2(n_55),
.B1(n_60),
.B2(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_18),
.A2(n_34),
.B1(n_41),
.B2(n_55),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_18),
.A2(n_55),
.B1(n_65),
.B2(n_66),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_21),
.B(n_340),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_19),
.B(n_341),
.Y(n_340)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_335),
.B(n_338),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_327),
.B(n_331),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_314),
.B(n_326),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_139),
.B(n_311),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_126),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_101),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_27),
.B(n_101),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_72),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_28),
.B(n_87),
.C(n_99),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_57),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_29),
.A2(n_30),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_42),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_31),
.A2(n_32),
.B1(n_57),
.B2(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_31),
.A2(n_32),
.B1(n_42),
.B2(n_43),
.Y(n_145)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_38),
.B(n_39),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_33),
.A2(n_38),
.B1(n_39),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_33),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_33),
.A2(n_38),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_33),
.A2(n_38),
.B1(n_181),
.B2(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_33),
.A2(n_38),
.B1(n_152),
.B2(n_182),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_33),
.A2(n_38),
.B1(n_195),
.B2(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_33),
.A2(n_38),
.B1(n_192),
.B2(n_248),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_33),
.A2(n_38),
.B1(n_241),
.B2(n_248),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_34),
.B(n_250),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_37),
.A2(n_115),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_37),
.A2(n_150),
.B1(n_240),
.B2(n_242),
.Y(n_239)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_41),
.A2(n_52),
.B(n_192),
.Y(n_229)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_44),
.A2(n_49),
.B1(n_56),
.B2(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_48),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_46),
.A2(n_63),
.A3(n_80),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_48),
.B(n_81),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_54),
.B1(n_56),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_56),
.B(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_49),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_49),
.A2(n_56),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_49),
.A2(n_56),
.B1(n_155),
.B2(n_186),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_49),
.A2(n_56),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_49),
.A2(n_56),
.B1(n_227),
.B2(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_53),
.A2(n_119),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_53),
.A2(n_156),
.B1(n_185),
.B2(n_265),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_57),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_68),
.B2(n_70),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_59),
.B1(n_70),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_58),
.A2(n_59),
.B1(n_68),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_58),
.A2(n_59),
.B1(n_90),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_58),
.A2(n_59),
.B1(n_124),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_58),
.A2(n_59),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_58),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_59),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_63),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_60),
.B(n_192),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_60),
.A2(n_62),
.A3(n_65),
.B1(n_202),
.B2(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_61),
.B(n_63),
.Y(n_216)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_66),
.B(n_192),
.Y(n_202)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_87),
.B1(n_99),
.B2(n_100),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_74),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_85),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_82),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_83),
.B1(n_84),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_78),
.A2(n_84),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_78),
.A2(n_84),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_78),
.A2(n_84),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_82),
.A2(n_96),
.B1(n_121),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_82),
.A2(n_121),
.B1(n_122),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_82),
.A2(n_121),
.B1(n_176),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_82),
.A2(n_173),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_89),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_94),
.C(n_97),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_89),
.B(n_129),
.C(n_132),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_98),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_97),
.B(n_135),
.C(n_137),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_109),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_120),
.C(n_123),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_111),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_296)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_123),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_126),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_127),
.B(n_128),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_136),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_138),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_164),
.B(n_310),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_162),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_141),
.B(n_162),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_146),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_142),
.B(n_145),
.Y(n_308)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_146),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_157),
.C(n_159),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_147),
.A2(n_148),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_149),
.B(n_153),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_157),
.B(n_159),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_158),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_160),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_305),
.B(n_309),
.Y(n_164)
);

OAI221xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_292),
.B1(n_303),
.B2(n_304),
.C(n_343),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_276),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_219),
.B(n_275),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_196),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_169),
.B(n_196),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_183),
.C(n_187),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_170),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_178),
.C(n_180),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_179),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_179),
.A2(n_289),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_179),
.A2(n_289),
.B1(n_322),
.B2(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_179),
.A2(n_289),
.B(n_329),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_183),
.A2(n_187),
.B1(n_188),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_189),
.A2(n_190),
.B1(n_194),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_191),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_210),
.B2(n_218),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_197),
.B(n_211),
.C(n_217),
.Y(n_277)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_199),
.B(n_205),
.C(n_209),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_206),
.Y(n_285)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_217),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_212),
.B(n_215),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_269),
.B(n_274),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_257),
.B(n_268),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_237),
.B(n_256),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_223),
.B(n_230),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_233),
.C(n_235),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_245),
.B(n_255),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_239),
.B(n_243),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_251),
.B(n_254),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_252),
.B(n_253),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_264),
.C(n_266),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_278),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_281),
.C(n_282),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_291),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_287),
.C(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_302),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_300),
.B2(n_301),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_296),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_301),
.C(n_302),
.Y(n_306)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_316),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_320),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_323),
.C(n_325),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_328),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_336),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_337),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);


endmodule