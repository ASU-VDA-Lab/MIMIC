module fake_jpeg_10100_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g13 ( 
.A(n_12),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_18),
.B(n_24),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_46),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_45),
.B1(n_14),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_22),
.B1(n_13),
.B2(n_24),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_14),
.B1(n_15),
.B2(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_18),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_28),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_52),
.Y(n_76)
);

AOI22x1_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_33),
.B1(n_21),
.B2(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_60),
.B1(n_23),
.B2(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_33),
.B1(n_14),
.B2(n_17),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_56),
.B1(n_61),
.B2(n_67),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_50),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_32),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_40),
.C(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_14),
.B1(n_21),
.B2(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_17),
.B1(n_25),
.B2(n_15),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_77),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_45),
.CI(n_39),
.CON(n_70),
.SN(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_72),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_44),
.CI(n_14),
.CON(n_72),
.SN(n_72)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_85),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_44),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_80),
.B1(n_88),
.B2(n_49),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_64),
.C(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_15),
.B1(n_44),
.B2(n_19),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_48),
.C(n_50),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_89),
.B1(n_68),
.B2(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_2),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_19),
.C(n_5),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_19),
.B1(n_5),
.B2(n_6),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_108),
.C(n_19),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_85),
.B1(n_82),
.B2(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_49),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_56),
.B1(n_52),
.B2(n_55),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_102),
.B1(n_109),
.B2(n_90),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_65),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_19),
.B(n_58),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_59),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_124),
.B1(n_97),
.B2(n_7),
.Y(n_139)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_70),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_91),
.C(n_103),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_72),
.B(n_75),
.C(n_73),
.D(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_131),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_134),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_108),
.C(n_101),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_93),
.B1(n_97),
.B2(n_87),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_111),
.B1(n_124),
.B2(n_115),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_136),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_120),
.B(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_121),
.B1(n_117),
.B2(n_113),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

AOI31xp67_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_149),
.A3(n_110),
.B(n_7),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_127),
.C(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_153),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_145),
.C(n_131),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_140),
.Y(n_161)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_129),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_155),
.A2(n_157),
.B(n_149),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_135),
.B1(n_138),
.B2(n_110),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_3),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_8),
.B(n_9),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_147),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_155),
.A3(n_152),
.B1(n_154),
.B2(n_151),
.C1(n_11),
.C2(n_7),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_160),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_167),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_170),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_165),
.C(n_166),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_167),
.C(n_11),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_12),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_173),
.Y(n_176)
);


endmodule