module fake_jpeg_16802_n_114 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_25),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_17),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_34),
.B(n_35),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_13),
.B1(n_21),
.B2(n_17),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_13),
.B1(n_21),
.B2(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_52),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_27),
.B1(n_16),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_50),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_16),
.B(n_22),
.C(n_18),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_14),
.B(n_2),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_32),
.B1(n_30),
.B2(n_36),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_67),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_25),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_68),
.C(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_36),
.B1(n_18),
.B2(n_14),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_19),
.B(n_14),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_45),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_14),
.C(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_40),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_79),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_57),
.C(n_54),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_46),
.B1(n_53),
.B2(n_41),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_64),
.B1(n_60),
.B2(n_59),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_63),
.C(n_54),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_74),
.B1(n_58),
.B2(n_67),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_72),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_75),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_19),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_78),
.B(n_58),
.C(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_64),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_81),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_1),
.B(n_2),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_93),
.B1(n_99),
.B2(n_3),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_5),
.Y(n_108)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_1),
.B(n_2),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_6),
.B(n_7),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_107),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_4),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_108),
.A2(n_109),
.B(n_5),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_6),
.C(n_10),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_111),
.B(n_107),
.Y(n_114)
);


endmodule