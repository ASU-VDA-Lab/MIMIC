module real_jpeg_32492_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_75, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_74, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_75;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_74;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_57;
wire n_65;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_55;
wire n_69;
wire n_58;
wire n_31;
wire n_49;
wire n_52;
wire n_67;
wire n_63;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_44;
wire n_60;
wire n_28;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_61;
wire n_71;
wire n_42;
wire n_22;
wire n_53;
wire n_39;
wire n_40;
wire n_36;
wire n_70;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_32;
wire n_48;
wire n_30;
wire n_56;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

OAI211xp5_ASAP7_75t_L g29 ( 
.A1(n_2),
.A2(n_30),
.B(n_33),
.C(n_41),
.Y(n_29)
);

AOI211xp5_ASAP7_75t_SL g42 ( 
.A1(n_2),
.A2(n_30),
.B(n_33),
.C(n_41),
.Y(n_42)
);

AOI321xp33_ASAP7_75t_L g19 ( 
.A1(n_3),
.A2(n_20),
.A3(n_23),
.B1(n_24),
.B2(n_58),
.C(n_62),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_4),
.A2(n_9),
.B1(n_26),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_4),
.B(n_14),
.C(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_5),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_8),
.C(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_9),
.A2(n_26),
.B(n_43),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_11),
.C(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_15),
.B(n_74),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_18),
.A2(n_22),
.B1(n_26),
.B2(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_20),
.A2(n_47),
.B(n_59),
.Y(n_58)
);

NOR4xp25_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_45),
.C(n_47),
.D(n_55),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_25),
.A2(n_45),
.B(n_60),
.C(n_61),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B(n_42),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_39),
.C(n_40),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.C(n_38),
.Y(n_35)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_75),
.Y(n_37)
);


endmodule