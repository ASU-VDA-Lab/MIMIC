module real_aes_4484_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_370;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_1049;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_1070;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_973;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_1006;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_1031;
wire n_432;
wire n_880;
wire n_1037;
wire n_1008;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_288;
wire n_1073;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_997;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1003;
wire n_1000;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_649;
wire n_293;
wire n_385;
wire n_358;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_314;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_756;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_0), .A2(n_21), .B1(n_670), .B2(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_1), .A2(n_51), .B1(n_812), .B2(n_813), .Y(n_811) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_2), .Y(n_294) );
AND2x4_ASAP7_75t_L g775 ( .A(n_2), .B(n_276), .Y(n_775) );
AND2x4_ASAP7_75t_L g780 ( .A(n_2), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_SL g302 ( .A(n_3), .Y(n_302) );
INVx1_ASAP7_75t_L g706 ( .A(n_4), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_5), .A2(n_111), .B1(n_355), .B2(n_356), .Y(n_604) );
XOR2x2_ASAP7_75t_L g525 ( .A(n_6), .B(n_526), .Y(n_525) );
XNOR2xp5_ASAP7_75t_L g580 ( .A(n_6), .B(n_526), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_7), .A2(n_181), .B1(n_383), .B2(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_8), .B(n_554), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_9), .A2(n_94), .B1(n_554), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_10), .A2(n_119), .B1(n_499), .B2(n_500), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_11), .A2(n_218), .B1(n_397), .B2(n_626), .Y(n_625) );
AOI21xp33_ASAP7_75t_SL g712 ( .A1(n_12), .A2(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g374 ( .A(n_13), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_14), .A2(n_232), .B1(n_424), .B2(n_591), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_15), .A2(n_85), .B1(n_784), .B2(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g538 ( .A(n_16), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_17), .A2(n_28), .B1(n_513), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_18), .A2(n_133), .B1(n_414), .B2(n_651), .Y(n_694) );
INVx1_ASAP7_75t_L g802 ( .A(n_19), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_20), .A2(n_154), .B1(n_523), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_22), .A2(n_57), .B1(n_649), .B2(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_23), .A2(n_203), .B1(n_419), .B2(n_421), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_24), .A2(n_220), .B1(n_435), .B2(n_437), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_25), .A2(n_83), .B1(n_772), .B2(n_776), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_26), .A2(n_115), .B1(n_504), .B2(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g612 ( .A(n_27), .Y(n_612) );
INVx1_ASAP7_75t_SL g886 ( .A(n_29), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_30), .A2(n_139), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g549 ( .A(n_31), .Y(n_549) );
INVx1_ASAP7_75t_L g1008 ( .A(n_32), .Y(n_1008) );
AOI22xp5_ASAP7_75t_L g1046 ( .A1(n_33), .A2(n_262), .B1(n_510), .B2(n_512), .Y(n_1046) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_34), .B(n_221), .Y(n_292) );
INVx1_ASAP7_75t_L g327 ( .A(n_34), .Y(n_327) );
INVxp67_ASAP7_75t_L g391 ( .A(n_34), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_35), .A2(n_97), .B1(n_779), .B2(n_791), .Y(n_817) );
INVx1_ASAP7_75t_L g1014 ( .A(n_36), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_37), .A2(n_135), .B1(n_421), .B2(n_577), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_38), .A2(n_230), .B1(n_478), .B2(n_614), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_39), .A2(n_76), .B1(n_522), .B2(n_619), .Y(n_1047) );
AOI21xp33_ASAP7_75t_SL g561 ( .A1(n_40), .A2(n_540), .B(n_562), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_41), .A2(n_158), .B1(n_419), .B2(n_619), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_42), .A2(n_75), .B1(n_361), .B2(n_363), .C(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_43), .B(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_44), .A2(n_93), .B1(n_737), .B2(n_738), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_45), .B(n_312), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_46), .A2(n_174), .B1(n_504), .B2(n_722), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_47), .A2(n_273), .B1(n_406), .B2(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g1023 ( .A(n_48), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_49), .A2(n_233), .B1(n_379), .B2(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g1062 ( .A(n_50), .Y(n_1062) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_51), .A2(n_587), .B(n_605), .Y(n_586) );
NAND4xp25_ASAP7_75t_L g605 ( .A(n_51), .B(n_588), .C(n_594), .D(n_601), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_52), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_53), .A2(n_281), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_54), .A2(n_78), .B1(n_397), .B2(n_399), .C(n_402), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_55), .A2(n_259), .B1(n_412), .B2(n_414), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_56), .A2(n_199), .B1(n_590), .B2(n_591), .Y(n_589) );
INVxp67_ASAP7_75t_R g804 ( .A(n_58), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_59), .A2(n_227), .B1(n_626), .B2(n_649), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_60), .A2(n_130), .B1(n_523), .B2(n_722), .Y(n_1000) );
INVx1_ASAP7_75t_L g1064 ( .A(n_61), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_62), .A2(n_252), .B1(n_307), .B2(n_330), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_63), .A2(n_172), .B1(n_532), .B2(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_64), .A2(n_120), .B1(n_412), .B2(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g289 ( .A(n_65), .Y(n_289) );
XNOR2x1_ASAP7_75t_L g677 ( .A(n_66), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g479 ( .A(n_67), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_68), .A2(n_229), .B1(n_406), .B2(n_408), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_69), .A2(n_189), .B1(n_505), .B2(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g774 ( .A(n_70), .Y(n_774) );
AND2x4_ASAP7_75t_L g777 ( .A(n_70), .B(n_289), .Y(n_777) );
INVx1_ASAP7_75t_SL g810 ( .A(n_70), .Y(n_810) );
INVx1_ASAP7_75t_L g381 ( .A(n_71), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_72), .A2(n_213), .B1(n_339), .B2(n_352), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_73), .A2(n_74), .B1(n_424), .B2(n_426), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_77), .A2(n_609), .B(n_611), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_79), .A2(n_210), .B1(n_784), .B2(n_809), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_80), .A2(n_167), .B1(n_511), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_81), .A2(n_121), .B1(n_753), .B2(n_1002), .Y(n_1001) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_82), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_84), .A2(n_200), .B1(n_376), .B2(n_379), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_86), .B(n_744), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_87), .A2(n_192), .B1(n_383), .B2(n_385), .Y(n_599) );
INVx1_ASAP7_75t_L g1059 ( .A(n_88), .Y(n_1059) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_89), .A2(n_268), .B1(n_334), .B2(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_90), .A2(n_239), .B1(n_419), .B2(n_603), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_91), .A2(n_250), .B1(n_508), .B2(n_531), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_92), .B(n_385), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_95), .A2(n_146), .B1(n_431), .B2(n_529), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_96), .A2(n_109), .B1(n_752), .B2(n_753), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_98), .A2(n_138), .B1(n_696), .B2(n_697), .Y(n_695) );
CKINVDCx16_ASAP7_75t_R g800 ( .A(n_99), .Y(n_800) );
AO22x2_ASAP7_75t_L g1004 ( .A1(n_100), .A2(n_178), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_101), .A2(n_175), .B1(n_779), .B2(n_782), .Y(n_778) );
XOR2x2_ASAP7_75t_L g996 ( .A(n_101), .B(n_997), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_101), .A2(n_1033), .B1(n_1035), .B2(n_1070), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_102), .B(n_1055), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_103), .A2(n_236), .B1(n_603), .B2(n_663), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_104), .A2(n_182), .B1(n_349), .B2(n_356), .Y(n_460) );
INVx1_ASAP7_75t_L g313 ( .A(n_105), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_105), .B(n_219), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_106), .A2(n_254), .B1(n_553), .B2(n_554), .Y(n_1027) );
INVx1_ASAP7_75t_L g597 ( .A(n_107), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_108), .A2(n_113), .B1(n_435), .B2(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_110), .A2(n_134), .B1(n_740), .B2(n_741), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_112), .A2(n_169), .B1(n_511), .B2(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g485 ( .A(n_114), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_116), .A2(n_209), .B1(n_424), .B2(n_426), .Y(n_533) );
INVx1_ASAP7_75t_L g832 ( .A(n_117), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_118), .A2(n_176), .B1(n_772), .B2(n_789), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_122), .A2(n_196), .B1(n_349), .B2(n_352), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_123), .A2(n_193), .B1(n_424), .B2(n_426), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_124), .A2(n_243), .B1(n_531), .B2(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_125), .B(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_126), .A2(n_155), .B1(n_744), .B2(n_745), .C(n_746), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_126), .A2(n_155), .B1(n_744), .B2(n_745), .C(n_746), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_127), .A2(n_187), .B1(n_334), .B2(n_355), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_128), .A2(n_211), .B1(n_435), .B2(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g715 ( .A(n_129), .Y(n_715) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_131), .A2(n_444), .B(n_462), .Y(n_443) );
INVx1_ASAP7_75t_L g465 ( .A(n_131), .Y(n_465) );
INVx1_ASAP7_75t_L g654 ( .A(n_132), .Y(n_654) );
XNOR2x1_ASAP7_75t_L g637 ( .A(n_136), .B(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_137), .A2(n_194), .B1(n_424), .B2(n_591), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_140), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_140), .A2(n_179), .B1(n_776), .B2(n_788), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_141), .A2(n_151), .B1(n_571), .B2(n_572), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_142), .A2(n_204), .B1(n_426), .B2(n_571), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_143), .A2(n_201), .B1(n_515), .B2(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g1016 ( .A(n_144), .Y(n_1016) );
INVx1_ASAP7_75t_L g547 ( .A(n_145), .Y(n_547) );
INVx1_ASAP7_75t_L g1011 ( .A(n_147), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_148), .A2(n_241), .B1(n_419), .B2(n_421), .Y(n_640) );
INVx1_ASAP7_75t_L g1044 ( .A(n_149), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_150), .A2(n_244), .B1(n_429), .B2(n_431), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_152), .A2(n_249), .B1(n_435), .B2(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g377 ( .A(n_153), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_156), .A2(n_162), .B1(n_487), .B2(n_491), .Y(n_568) );
INVx1_ASAP7_75t_L g676 ( .A(n_157), .Y(n_676) );
INVx1_ASAP7_75t_L g1041 ( .A(n_159), .Y(n_1041) );
AOI21xp33_ASAP7_75t_SL g1057 ( .A1(n_160), .A2(n_540), .B(n_1058), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_161), .A2(n_171), .B1(n_505), .B2(n_663), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_163), .A2(n_260), .B1(n_812), .B2(n_813), .Y(n_821) );
INVx1_ASAP7_75t_L g835 ( .A(n_164), .Y(n_835) );
INVx1_ASAP7_75t_L g833 ( .A(n_165), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_166), .B(n_495), .Y(n_560) );
INVx1_ASAP7_75t_L g452 ( .A(n_168), .Y(n_452) );
INVx1_ASAP7_75t_L g493 ( .A(n_170), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_173), .A2(n_258), .B1(n_579), .B2(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g476 ( .A(n_177), .Y(n_476) );
INVx1_ASAP7_75t_L g366 ( .A(n_180), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_183), .A2(n_255), .B1(n_435), .B2(n_535), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_184), .A2(n_235), .B1(n_651), .B2(n_652), .C(n_653), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_185), .A2(n_251), .B1(n_553), .B2(n_554), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_186), .A2(n_265), .B1(n_355), .B2(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g690 ( .A(n_188), .Y(n_690) );
OA22x2_ASAP7_75t_L g318 ( .A1(n_190), .A2(n_221), .B1(n_312), .B2(n_316), .Y(n_318) );
INVx1_ASAP7_75t_L g344 ( .A(n_190), .Y(n_344) );
INVx1_ASAP7_75t_L g545 ( .A(n_191), .Y(n_545) );
AOI21xp5_ASAP7_75t_SL g362 ( .A1(n_195), .A2(n_363), .B(n_365), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_197), .A2(n_215), .B1(n_510), .B2(n_512), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_198), .A2(n_280), .B1(n_419), .B2(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_202), .A2(n_222), .B1(n_307), .B2(n_330), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_205), .A2(n_226), .B1(n_614), .B2(n_626), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_206), .A2(n_274), .B1(n_424), .B2(n_426), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_207), .A2(n_263), .B1(n_590), .B2(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g1050 ( .A(n_208), .Y(n_1050) );
INVx1_ASAP7_75t_L g563 ( .A(n_212), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_214), .B(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_216), .A2(n_245), .B1(n_532), .B2(n_579), .Y(n_578) );
CKINVDCx6p67_ASAP7_75t_R g798 ( .A(n_217), .Y(n_798) );
INVx1_ASAP7_75t_L g329 ( .A(n_219), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_219), .B(n_342), .Y(n_372) );
OAI21xp33_ASAP7_75t_L g345 ( .A1(n_221), .A2(n_240), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g359 ( .A(n_223), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_224), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_225), .A2(n_266), .B1(n_334), .B2(n_339), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_228), .A2(n_242), .B1(n_779), .B2(n_791), .Y(n_790) );
XOR2xp5_ASAP7_75t_L g1035 ( .A(n_231), .B(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g557 ( .A(n_234), .Y(n_557) );
INVxp67_ASAP7_75t_SL g748 ( .A(n_237), .Y(n_748) );
INVx1_ASAP7_75t_SL g1067 ( .A(n_238), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_240), .B(n_269), .Y(n_293) );
INVx1_ASAP7_75t_L g315 ( .A(n_240), .Y(n_315) );
INVx1_ASAP7_75t_L g489 ( .A(n_246), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_247), .A2(n_257), .B1(n_648), .B2(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g887 ( .A(n_248), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_253), .A2(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_SL g1049 ( .A(n_256), .Y(n_1049) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_261), .A2(n_376), .B(n_451), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_264), .A2(n_272), .B1(n_435), .B2(n_437), .Y(n_666) );
INVx1_ASAP7_75t_L g747 ( .A(n_267), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_269), .B(n_322), .Y(n_321) );
XNOR2x1_ASAP7_75t_L g472 ( .A(n_270), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g1019 ( .A(n_271), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_275), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g781 ( .A(n_276), .Y(n_781) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_276), .Y(n_1072) );
INVx1_ASAP7_75t_L g1021 ( .A(n_277), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_278), .Y(n_403) );
INVx1_ASAP7_75t_L g542 ( .A(n_279), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_295), .B(n_765), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND3xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .C(n_294), .Y(n_286) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_287), .B(n_1030), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_287), .B(n_1031), .Y(n_1034) );
AOI21xp5_ASAP7_75t_L g1073 ( .A1(n_287), .A2(n_294), .B(n_810), .Y(n_1073) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AO21x1_ASAP7_75t_L g1071 ( .A1(n_288), .A2(n_1072), .B(n_1073), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g773 ( .A(n_289), .B(n_774), .Y(n_773) );
AND3x4_ASAP7_75t_L g809 ( .A(n_289), .B(n_780), .C(n_810), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g1030 ( .A(n_290), .B(n_1031), .Y(n_1030) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AO21x2_ASAP7_75t_L g368 ( .A1(n_291), .A2(n_369), .B(n_371), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g1031 ( .A(n_294), .Y(n_1031) );
XNOR2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_466), .Y(n_295) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_442), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
OA22x2_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_392), .B1(n_440), .B2(n_441), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
XNOR2x1_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
XNOR2xp5_ASAP7_75t_L g441 ( .A(n_302), .B(n_303), .Y(n_441) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_357), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_347), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_333), .Y(n_305) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_319), .Y(n_307) );
AND2x4_ASAP7_75t_L g330 ( .A(n_308), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g349 ( .A(n_308), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g352 ( .A(n_308), .B(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g420 ( .A(n_308), .B(n_350), .Y(n_420) );
AND2x4_ASAP7_75t_L g422 ( .A(n_308), .B(n_336), .Y(n_422) );
AND2x4_ASAP7_75t_L g425 ( .A(n_308), .B(n_319), .Y(n_425) );
AND2x2_ASAP7_75t_L g427 ( .A(n_308), .B(n_331), .Y(n_427) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_317), .Y(n_308) );
AND2x2_ASAP7_75t_L g364 ( .A(n_309), .B(n_318), .Y(n_364) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g335 ( .A(n_310), .B(n_318), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
NAND2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx2_ASAP7_75t_L g316 ( .A(n_312), .Y(n_316) );
INVx3_ASAP7_75t_L g322 ( .A(n_312), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g328 ( .A(n_312), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g346 ( .A(n_312), .Y(n_346) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_312), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_313), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
OAI21xp5_ASAP7_75t_L g390 ( .A1(n_315), .A2(n_346), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g389 ( .A(n_318), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g376 ( .A(n_319), .B(n_364), .Y(n_376) );
AND2x4_ASAP7_75t_L g383 ( .A(n_319), .B(n_335), .Y(n_383) );
AND2x4_ASAP7_75t_L g398 ( .A(n_319), .B(n_364), .Y(n_398) );
AND2x2_ASAP7_75t_L g407 ( .A(n_319), .B(n_335), .Y(n_407) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .Y(n_319) );
INVx2_ASAP7_75t_L g332 ( .A(n_320), .Y(n_332) );
OR2x2_ASAP7_75t_L g337 ( .A(n_320), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g350 ( .A(n_320), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g386 ( .A(n_320), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_322), .B(n_327), .Y(n_326) );
INVxp67_ASAP7_75t_L g342 ( .A(n_322), .Y(n_342) );
NAND3xp33_ASAP7_75t_L g371 ( .A(n_323), .B(n_341), .C(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g331 ( .A(n_324), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g338 ( .A(n_325), .Y(n_338) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g361 ( .A(n_331), .B(n_335), .Y(n_361) );
AND2x2_ASAP7_75t_L g363 ( .A(n_331), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g379 ( .A(n_331), .B(n_340), .Y(n_379) );
AND2x2_ASAP7_75t_L g401 ( .A(n_331), .B(n_335), .Y(n_401) );
AND2x4_ASAP7_75t_L g413 ( .A(n_331), .B(n_364), .Y(n_413) );
AND2x4_ASAP7_75t_L g416 ( .A(n_331), .B(n_340), .Y(n_416) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
AND2x4_ASAP7_75t_L g355 ( .A(n_335), .B(n_350), .Y(n_355) );
AND2x4_ASAP7_75t_L g430 ( .A(n_335), .B(n_353), .Y(n_430) );
AND2x2_ASAP7_75t_L g436 ( .A(n_335), .B(n_350), .Y(n_436) );
AND2x2_ASAP7_75t_L g683 ( .A(n_335), .B(n_350), .Y(n_683) );
AND2x4_ASAP7_75t_L g339 ( .A(n_336), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g433 ( .A(n_336), .B(n_340), .Y(n_433) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g353 ( .A(n_337), .Y(n_353) );
INVx1_ASAP7_75t_L g351 ( .A(n_338), .Y(n_351) );
AND2x4_ASAP7_75t_L g356 ( .A(n_340), .B(n_350), .Y(n_356) );
AND2x4_ASAP7_75t_L g439 ( .A(n_340), .B(n_350), .Y(n_439) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_345), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_354), .Y(n_347) );
NOR3xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_373), .C(n_380), .Y(n_357) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B(n_362), .Y(n_358) );
INVx2_ASAP7_75t_L g652 ( .A(n_360), .Y(n_652) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_367), .Y(n_404) );
INVx2_ASAP7_75t_L g565 ( .A(n_367), .Y(n_565) );
INVx2_ASAP7_75t_SL g656 ( .A(n_367), .Y(n_656) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g454 ( .A(n_368), .Y(n_454) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_370), .B(n_388), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_377), .B2(n_378), .Y(n_373) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI21xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_382), .B(n_384), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx4_ASAP7_75t_L g691 ( .A(n_385), .Y(n_691) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
AND2x4_ASAP7_75t_L g410 ( .A(n_386), .B(n_389), .Y(n_410) );
AND2x2_ASAP7_75t_L g449 ( .A(n_386), .B(n_389), .Y(n_449) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_392), .Y(n_440) );
XNOR2x1_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_417), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_405), .C(n_411), .Y(n_395) );
INVx4_ASAP7_75t_L g1015 ( .A(n_397), .Y(n_1015) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx3_ASAP7_75t_L g478 ( .A(n_398), .Y(n_478) );
INVx1_ASAP7_75t_L g541 ( .A(n_398), .Y(n_541) );
BUFx3_ASAP7_75t_L g670 ( .A(n_398), .Y(n_670) );
INVx2_ASAP7_75t_L g610 ( .A(n_399), .Y(n_610) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g456 ( .A(n_400), .Y(n_456) );
INVx2_ASAP7_75t_L g551 ( .A(n_400), .Y(n_551) );
INVx2_ASAP7_75t_L g688 ( .A(n_400), .Y(n_688) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g497 ( .A(n_401), .Y(n_497) );
BUFx3_ASAP7_75t_L g675 ( .A(n_401), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx2_ASAP7_75t_L g693 ( .A(n_404), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_404), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g543 ( .A(n_406), .Y(n_543) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g483 ( .A(n_407), .Y(n_483) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_407), .Y(n_626) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx3_ASAP7_75t_L g499 ( .A(n_409), .Y(n_499) );
INVx4_ASAP7_75t_L g614 ( .A(n_409), .Y(n_614) );
INVx2_ASAP7_75t_L g744 ( .A(n_409), .Y(n_744) );
INVx5_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx4f_ASAP7_75t_L g553 ( .A(n_410), .Y(n_553) );
BUFx2_ASAP7_75t_L g711 ( .A(n_410), .Y(n_711) );
INVx2_ASAP7_75t_L g546 ( .A(n_412), .Y(n_546) );
BUFx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_413), .Y(n_447) );
INVx2_ASAP7_75t_L g488 ( .A(n_413), .Y(n_488) );
INVx2_ASAP7_75t_L g673 ( .A(n_413), .Y(n_673) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_413), .Y(n_713) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_415), .A2(n_545), .B1(n_546), .B2(n_547), .Y(n_544) );
INVx3_ASAP7_75t_L g628 ( .A(n_415), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_415), .A2(n_1019), .B1(n_1020), .B2(n_1021), .Y(n_1018) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_416), .Y(n_649) );
NAND4xp25_ASAP7_75t_SL g417 ( .A(n_418), .B(n_423), .C(n_428), .D(n_434), .Y(n_417) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx12f_ASAP7_75t_L g511 ( .A(n_420), .Y(n_511) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_420), .Y(n_577) );
BUFx3_ASAP7_75t_L g752 ( .A(n_421), .Y(n_752) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_422), .Y(n_513) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_422), .Y(n_529) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_422), .Y(n_603) );
BUFx12f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g516 ( .A(n_425), .Y(n_516) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_425), .Y(n_571) );
BUFx2_ASAP7_75t_SL g1006 ( .A(n_426), .Y(n_1006) );
INVx1_ASAP7_75t_L g1051 ( .A(n_426), .Y(n_1051) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g520 ( .A(n_427), .Y(n_520) );
BUFx5_ASAP7_75t_L g572 ( .A(n_427), .Y(n_572) );
BUFx3_ASAP7_75t_L g591 ( .A(n_427), .Y(n_591) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx12f_ASAP7_75t_L g505 ( .A(n_430), .Y(n_505) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_430), .Y(n_531) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_430), .Y(n_579) );
BUFx3_ASAP7_75t_L g623 ( .A(n_430), .Y(n_623) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g508 ( .A(n_432), .Y(n_508) );
INVx3_ASAP7_75t_L g593 ( .A(n_432), .Y(n_593) );
INVx5_ASAP7_75t_L g663 ( .A(n_432), .Y(n_663) );
INVx6_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx12f_ASAP7_75t_L g532 ( .A(n_433), .Y(n_532) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx8_ASAP7_75t_L g522 ( .A(n_436), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_437), .Y(n_523) );
INVx4_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx4_ASAP7_75t_L g535 ( .A(n_438), .Y(n_535) );
INVx2_ASAP7_75t_L g574 ( .A(n_438), .Y(n_574) );
INVx4_ASAP7_75t_L g619 ( .A(n_438), .Y(n_619) );
INVx1_ASAP7_75t_L g724 ( .A(n_438), .Y(n_724) );
INVx8_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_457), .Y(n_444) );
INVxp67_ASAP7_75t_L g463 ( .A(n_445), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .C(n_450), .D(n_455), .Y(n_445) );
INVx2_ASAP7_75t_L g1020 ( .A(n_447), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx4_ASAP7_75t_L g554 ( .A(n_453), .Y(n_554) );
INVx4_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g501 ( .A(n_454), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_457), .B(n_465), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .C(n_460), .D(n_461), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_631), .B2(n_632), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B1(n_581), .B2(n_630), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
XOR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_524), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_502), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .C(n_492), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_479), .B2(n_480), .Y(n_475) );
INVx2_ASAP7_75t_L g737 ( .A(n_477), .Y(n_737) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g1017 ( .A(n_482), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g648 ( .A(n_483), .Y(n_648) );
INVx1_ASAP7_75t_L g697 ( .A(n_483), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_489), .B2(n_490), .Y(n_484) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_SL g651 ( .A(n_488), .Y(n_651) );
INVx4_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI21xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B(n_498), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g717 ( .A(n_496), .Y(n_717) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g1056 ( .A(n_497), .Y(n_1056) );
INVx4_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_501), .B(n_597), .Y(n_596) );
AND4x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_509), .C(n_514), .D(n_521), .Y(n_502) );
BUFx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g1043 ( .A(n_507), .Y(n_1043) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx12f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_511), .Y(n_759) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g590 ( .A(n_516), .Y(n_590) );
INVx1_ASAP7_75t_L g1005 ( .A(n_516), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_516), .A2(n_1049), .B1(n_1050), .B2(n_1051), .Y(n_1048) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI22x1_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_555), .B1(n_556), .B2(n_580), .Y(n_524) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_536), .Y(n_526) );
AND4x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .C(n_533), .D(n_534), .Y(n_527) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_531), .Y(n_1002) );
BUFx3_ASAP7_75t_L g753 ( .A(n_532), .Y(n_753) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_544), .C(n_548), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B1(n_542), .B2(n_543), .Y(n_537) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g696 ( .A(n_541), .Y(n_696) );
OAI21xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B(n_552), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g1060 ( .A(n_554), .Y(n_1060) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
XNOR2x1_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NOR4xp75_ASAP7_75t_L g558 ( .A(n_559), .B(n_566), .C(n_569), .D(n_575), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_570), .B(n_573), .Y(n_569) );
BUFx3_ASAP7_75t_L g757 ( .A(n_572), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_576), .B(n_578), .Y(n_575) );
INVx1_ASAP7_75t_L g630 ( .A(n_581), .Y(n_630) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_606), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND3x1_ASAP7_75t_L g587 ( .A(n_588), .B(n_594), .C(n_601), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
XNOR2x1_ASAP7_75t_L g606 ( .A(n_607), .B(n_629), .Y(n_606) );
NAND4xp75_ASAP7_75t_L g607 ( .A(n_608), .B(n_616), .C(n_620), .D(n_624), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_615), .Y(n_611) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
BUFx3_ASAP7_75t_L g738 ( .A(n_626), .Y(n_738) );
INVx3_ASAP7_75t_L g1068 ( .A(n_626), .Y(n_1068) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI22x1_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_699), .B2(n_700), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OA22x2_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_657), .B1(n_658), .B2(n_698), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g698 ( .A(n_636), .Y(n_698) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND4xp75_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .C(n_645), .D(n_650), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
BUFx3_ASAP7_75t_L g741 ( .A(n_649), .Y(n_741) );
INVx3_ASAP7_75t_L g1065 ( .A(n_649), .Y(n_1065) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NOR2xp33_ASAP7_75t_R g746 ( .A(n_655), .B(n_747), .Y(n_746) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
XNOR2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_677), .Y(n_658) );
XOR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_676), .Y(n_659) );
NOR2x1_ASAP7_75t_L g660 ( .A(n_661), .B(n_667), .Y(n_660) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .C(n_665), .D(n_666), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .C(n_671), .D(n_674), .Y(n_667) );
INVx2_ASAP7_75t_L g1063 ( .A(n_672), .Y(n_1063) );
INVx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g1026 ( .A(n_675), .Y(n_1026) );
OR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_686), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .C(n_684), .D(n_685), .Y(n_679) );
BUFx4f_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_683), .Y(n_722) );
NAND3xp33_ASAP7_75t_SL g686 ( .A(n_687), .B(n_694), .C(n_695), .Y(n_686) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_688), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B(n_692), .Y(n_689) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_732), .B1(n_762), .B2(n_763), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g762 ( .A(n_703), .Y(n_762) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI21x1_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B(n_726), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_705), .B(n_718), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
NOR2xp67_ASAP7_75t_L g707 ( .A(n_708), .B(n_719), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_716), .C(n_718), .Y(n_708) );
INVx1_ASAP7_75t_L g730 ( .A(n_709), .Y(n_730) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
BUFx3_ASAP7_75t_L g740 ( .A(n_713), .Y(n_740) );
INVxp67_ASAP7_75t_L g728 ( .A(n_716), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_719), .Y(n_731) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .C(n_723), .D(n_725), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_731), .Y(n_726) );
NOR3xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .C(n_730), .Y(n_727) );
AO22x2_ASAP7_75t_SL g732 ( .A1(n_733), .A2(n_748), .B1(n_749), .B2(n_760), .Y(n_732) );
AO22x2_ASAP7_75t_L g764 ( .A1(n_733), .A2(n_748), .B1(n_749), .B2(n_760), .Y(n_764) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_742), .C(n_748), .Y(n_733) );
INVxp67_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND4xp75_ASAP7_75t_SL g760 ( .A(n_735), .B(n_750), .C(n_755), .D(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_755), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g1010 ( .A(n_752), .Y(n_1010) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .Y(n_755) );
INVx1_ASAP7_75t_L g1009 ( .A(n_759), .Y(n_1009) );
INVx2_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
OAI221xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_992), .B1(n_995), .B2(n_1028), .C(n_1032), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_858), .B(n_883), .C(n_889), .Y(n_766) );
OAI211xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_792), .B(n_822), .C(n_841), .Y(n_767) );
INVx1_ASAP7_75t_L g943 ( .A(n_768), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_785), .Y(n_768) );
AND2x2_ASAP7_75t_L g839 ( .A(n_769), .B(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g869 ( .A(n_769), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_769), .B(n_884), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_769), .B(n_884), .Y(n_969) );
NOR3xp33_ASAP7_75t_L g988 ( .A(n_769), .B(n_874), .C(n_989), .Y(n_988) );
INVx3_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OR2x2_ASAP7_75t_L g852 ( .A(n_770), .B(n_785), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_770), .B(n_845), .Y(n_913) );
AND2x2_ASAP7_75t_L g949 ( .A(n_770), .B(n_950), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_770), .B(n_785), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_770), .B(n_877), .Y(n_975) );
AND2x2_ASAP7_75t_L g986 ( .A(n_770), .B(n_786), .Y(n_986) );
AND2x4_ASAP7_75t_L g770 ( .A(n_771), .B(n_778), .Y(n_770) );
AND2x2_ASAP7_75t_L g772 ( .A(n_773), .B(n_775), .Y(n_772) );
AND2x4_ASAP7_75t_L g779 ( .A(n_773), .B(n_780), .Y(n_779) );
AND2x4_ASAP7_75t_L g788 ( .A(n_773), .B(n_775), .Y(n_788) );
AND2x2_ASAP7_75t_L g812 ( .A(n_773), .B(n_775), .Y(n_812) );
AND2x4_ASAP7_75t_L g776 ( .A(n_775), .B(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g789 ( .A(n_775), .B(n_777), .Y(n_789) );
AND2x2_ASAP7_75t_L g813 ( .A(n_775), .B(n_777), .Y(n_813) );
INVx2_ASAP7_75t_L g805 ( .A(n_776), .Y(n_805) );
AND2x4_ASAP7_75t_L g784 ( .A(n_777), .B(n_780), .Y(n_784) );
AND2x4_ASAP7_75t_L g791 ( .A(n_777), .B(n_780), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_777), .B(n_780), .Y(n_799) );
INVx3_ASAP7_75t_L g797 ( .A(n_779), .Y(n_797) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
INVx3_ASAP7_75t_L g866 ( .A(n_785), .Y(n_866) );
AND2x2_ASAP7_75t_L g870 ( .A(n_785), .B(n_795), .Y(n_870) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g877 ( .A(n_786), .B(n_795), .Y(n_877) );
AND2x2_ASAP7_75t_L g908 ( .A(n_786), .B(n_840), .Y(n_908) );
OR2x2_ASAP7_75t_L g918 ( .A(n_786), .B(n_795), .Y(n_918) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_790), .Y(n_786) );
INVx3_ASAP7_75t_L g803 ( .A(n_788), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_806), .Y(n_792) );
INVx2_ASAP7_75t_L g896 ( .A(n_793), .Y(n_896) );
O2A1O1Ixp33_ASAP7_75t_SL g953 ( .A1(n_793), .A2(n_824), .B(n_954), .C(n_956), .Y(n_953) );
BUFx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_794), .B(n_843), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_794), .B(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g903 ( .A(n_794), .Y(n_903) );
AND2x2_ASAP7_75t_L g936 ( .A(n_794), .B(n_914), .Y(n_936) );
O2A1O1Ixp33_ASAP7_75t_L g940 ( .A1(n_794), .A2(n_941), .B(n_942), .C(n_943), .Y(n_940) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx3_ASAP7_75t_L g840 ( .A(n_795), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_795), .B(n_829), .Y(n_882) );
OR2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_801), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B1(n_799), .B2(n_800), .Y(n_796) );
OAI221xp5_ASAP7_75t_L g885 ( .A1(n_797), .A2(n_799), .B1(n_886), .B2(n_887), .C(n_888), .Y(n_885) );
INVx1_ASAP7_75t_L g994 ( .A(n_797), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_799), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_803), .B1(n_804), .B2(n_805), .Y(n_801) );
AND2x2_ASAP7_75t_L g828 ( .A(n_806), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g906 ( .A(n_806), .Y(n_906) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_814), .Y(n_806) );
CKINVDCx6p67_ASAP7_75t_R g825 ( .A(n_807), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_807), .B(n_819), .Y(n_843) );
INVx1_ASAP7_75t_L g850 ( .A(n_807), .Y(n_850) );
AND2x2_ASAP7_75t_L g862 ( .A(n_807), .B(n_863), .Y(n_862) );
OR2x2_ASAP7_75t_L g933 ( .A(n_807), .B(n_819), .Y(n_933) );
AND2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_811), .Y(n_807) );
INVx1_ASAP7_75t_L g831 ( .A(n_809), .Y(n_831) );
INVx1_ASAP7_75t_L g838 ( .A(n_812), .Y(n_838) );
INVx1_ASAP7_75t_L g836 ( .A(n_813), .Y(n_836) );
AND2x2_ASAP7_75t_SL g959 ( .A(n_814), .B(n_825), .Y(n_959) );
AND2x2_ASAP7_75t_L g966 ( .A(n_814), .B(n_895), .Y(n_966) );
OR2x2_ASAP7_75t_L g972 ( .A(n_814), .B(n_863), .Y(n_972) );
INVxp33_ASAP7_75t_L g979 ( .A(n_814), .Y(n_979) );
AND2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_818), .Y(n_814) );
INVx1_ASAP7_75t_L g827 ( .A(n_815), .Y(n_827) );
AND2x2_ASAP7_75t_L g855 ( .A(n_815), .B(n_819), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
AND2x2_ASAP7_75t_L g826 ( .A(n_818), .B(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_818), .B(n_849), .Y(n_930) );
OAI222xp33_ASAP7_75t_L g963 ( .A1(n_818), .A2(n_947), .B1(n_952), .B2(n_964), .C1(n_965), .C2(n_967), .Y(n_963) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
AND2x2_ASAP7_75t_L g863 ( .A(n_819), .B(n_827), .Y(n_863) );
AOI322xp5_ASAP7_75t_L g912 ( .A1(n_819), .A2(n_866), .A3(n_868), .B1(n_903), .B2(n_913), .C1(n_914), .C2(n_916), .Y(n_912) );
AND2x4_ASAP7_75t_SL g819 ( .A(n_820), .B(n_821), .Y(n_819) );
OAI21xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_828), .B(n_839), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
AND2x2_ASAP7_75t_L g856 ( .A(n_825), .B(n_857), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_825), .B(n_855), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_825), .B(n_829), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_825), .B(n_871), .Y(n_876) );
AND2x2_ASAP7_75t_L g899 ( .A(n_825), .B(n_827), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_825), .A2(n_905), .B1(n_906), .B2(n_907), .Y(n_904) );
AND2x2_ASAP7_75t_L g924 ( .A(n_825), .B(n_863), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_825), .B(n_902), .Y(n_944) );
AND2x2_ASAP7_75t_L g894 ( .A(n_826), .B(n_895), .Y(n_894) );
AND2x2_ASAP7_75t_L g902 ( .A(n_826), .B(n_829), .Y(n_902) );
INVx1_ASAP7_75t_L g917 ( .A(n_826), .Y(n_917) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_827), .B(n_849), .Y(n_848) );
AND2x2_ASAP7_75t_L g881 ( .A(n_827), .B(n_849), .Y(n_881) );
INVx1_ASAP7_75t_L g911 ( .A(n_827), .Y(n_911) );
INVx1_ASAP7_75t_L g846 ( .A(n_829), .Y(n_846) );
CKINVDCx6p67_ASAP7_75t_R g857 ( .A(n_829), .Y(n_857) );
AND2x2_ASAP7_75t_L g920 ( .A(n_829), .B(n_840), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_829), .B(n_848), .Y(n_952) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_829), .B(n_840), .Y(n_984) );
OR2x6_ASAP7_75t_SL g829 ( .A(n_830), .B(n_834), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_836), .B1(n_837), .B2(n_838), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_840), .B(n_852), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_840), .B(n_869), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_840), .B(n_955), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g990 ( .A(n_840), .B(n_857), .Y(n_990) );
O2A1O1Ixp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_844), .B(n_851), .C(n_853), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_847), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_845), .B(n_862), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_845), .B(n_908), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g978 ( .A(n_845), .B(n_979), .Y(n_978) );
INVx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g895 ( .A(n_849), .B(n_857), .Y(n_895) );
AND2x2_ASAP7_75t_L g901 ( .A(n_849), .B(n_902), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_849), .B(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
AOI221xp5_ASAP7_75t_L g935 ( .A1(n_851), .A2(n_884), .B1(n_936), .B2(n_937), .C(n_939), .Y(n_935) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
INVx1_ASAP7_75t_L g871 ( .A(n_855), .Y(n_871) );
AND2x2_ASAP7_75t_L g914 ( .A(n_855), .B(n_915), .Y(n_914) );
AND2x2_ASAP7_75t_L g955 ( .A(n_855), .B(n_895), .Y(n_955) );
INVxp67_ASAP7_75t_L g973 ( .A(n_856), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_857), .B(n_866), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_857), .B(n_877), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_857), .B(n_908), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_857), .B(n_924), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_857), .B(n_930), .Y(n_929) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_857), .B(n_918), .Y(n_934) );
OAI221xp5_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_865), .B1(n_867), .B2(n_871), .C(n_872), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_864), .Y(n_860) );
OAI221xp5_ASAP7_75t_L g980 ( .A1(n_861), .A2(n_974), .B1(n_981), .B2(n_985), .C(n_987), .Y(n_980) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
OAI21xp33_ASAP7_75t_L g931 ( .A1(n_862), .A2(n_932), .B(n_934), .Y(n_931) );
INVx1_ASAP7_75t_L g874 ( .A(n_863), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_863), .B(n_920), .Y(n_919) );
OAI321xp33_ASAP7_75t_L g970 ( .A1(n_864), .A2(n_971), .A3(n_973), .B1(n_974), .B2(n_975), .C(n_976), .Y(n_970) );
INVx3_ASAP7_75t_L g879 ( .A(n_866), .Y(n_879) );
INVx1_ASAP7_75t_L g967 ( .A(n_866), .Y(n_967) );
O2A1O1Ixp33_ASAP7_75t_SL g909 ( .A1(n_867), .A2(n_910), .B(n_912), .C(n_921), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_870), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_868), .B(n_958), .Y(n_957) );
INVx3_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g905 ( .A(n_870), .Y(n_905) );
NAND3xp33_ASAP7_75t_L g976 ( .A(n_870), .B(n_881), .C(n_913), .Y(n_976) );
O2A1O1Ixp33_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_876), .B(n_877), .C(n_878), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
INVx1_ASAP7_75t_L g915 ( .A(n_875), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_876), .B(n_894), .Y(n_893) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_879), .B(n_921), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_879), .B(n_884), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
CKINVDCx16_ASAP7_75t_R g991 ( .A(n_883), .Y(n_991) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
BUFx3_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx2_ASAP7_75t_L g921 ( .A(n_885), .Y(n_921) );
NAND5xp2_ASAP7_75t_L g889 ( .A(n_890), .B(n_935), .C(n_948), .D(n_960), .E(n_977), .Y(n_889) );
AOI211xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_892), .B(n_909), .C(n_922), .Y(n_890) );
OAI221xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_896), .B1(n_897), .B2(n_898), .C(n_900), .Y(n_892) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_903), .B(n_904), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_903), .B(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g947 ( .A(n_908), .Y(n_947) );
INVx1_ASAP7_75t_L g983 ( .A(n_911), .Y(n_983) );
OAI21xp33_ASAP7_75t_SL g916 ( .A1(n_917), .A2(n_918), .B(n_919), .Y(n_916) );
INVx1_ASAP7_75t_L g950 ( .A(n_918), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_920), .B(n_959), .Y(n_958) );
CKINVDCx16_ASAP7_75t_R g941 ( .A(n_921), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_921), .B(n_947), .Y(n_946) );
OAI221xp5_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_925), .B1(n_926), .B2(n_928), .C(n_931), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_924), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g961 ( .A(n_938), .Y(n_961) );
OAI21xp33_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_944), .B(n_945), .Y(n_939) );
AOI211xp5_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_951), .B(n_953), .C(n_957), .Y(n_948) );
A2O1A1Ixp33_ASAP7_75t_L g977 ( .A1(n_949), .A2(n_978), .B(n_980), .C(n_991), .Y(n_977) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g962 ( .A(n_956), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_962), .B1(n_963), .B2(n_968), .C(n_970), .Y(n_960) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVxp67_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_984), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g992 ( .A(n_993), .Y(n_992) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g997 ( .A(n_998), .B(n_1003), .C(n_1012), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1001), .Y(n_999) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1002), .Y(n_1040) );
NOR2x1_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1007), .Y(n_1003) );
OAI22x1_ASAP7_75t_SL g1007 ( .A1(n_1008), .A2(n_1009), .B1(n_1010), .B2(n_1011), .Y(n_1007) );
NOR3xp33_ASAP7_75t_SL g1012 ( .A(n_1013), .B(n_1018), .C(n_1022), .Y(n_1012) );
OAI22xp5_ASAP7_75t_SL g1013 ( .A1(n_1014), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1013) );
OAI21xp33_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1024), .B(n_1027), .Y(n_1022) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
HB1xp67_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1052), .Y(n_1037) );
NOR3xp33_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1045), .C(n_1048), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_1040), .A2(n_1041), .B1(n_1042), .B2(n_1044), .Y(n_1039) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
NAND2xp5_ASAP7_75t_SL g1045 ( .A(n_1046), .B(n_1047), .Y(n_1045) );
NOR3xp33_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1061), .C(n_1066), .Y(n_1052) );
NAND2xp5_ASAP7_75t_SL g1053 ( .A(n_1054), .B(n_1057), .Y(n_1053) );
BUFx3_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
NOR2xp33_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_1062), .A2(n_1063), .B1(n_1064), .B2(n_1065), .Y(n_1061) );
OAI21xp5_ASAP7_75t_L g1066 ( .A1(n_1067), .A2(n_1068), .B(n_1069), .Y(n_1066) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
endmodule