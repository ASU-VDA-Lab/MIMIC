module fake_jpeg_23328_n_290 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_41),
.B(n_47),
.Y(n_68)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_19),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_35),
.C(n_23),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_31),
.B1(n_27),
.B2(n_35),
.Y(n_66)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_35),
.B1(n_36),
.B2(n_20),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_42),
.B(n_36),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_33),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_48),
.B1(n_31),
.B2(n_27),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_67),
.B1(n_71),
.B2(n_75),
.Y(n_104)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_85),
.B(n_20),
.C(n_24),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_82),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_76),
.B(n_77),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_23),
.B1(n_26),
.B2(n_32),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_88),
.B1(n_36),
.B2(n_24),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_34),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_83),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_34),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_24),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_38),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_40),
.A2(n_23),
.B1(n_26),
.B2(n_18),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_42),
.B1(n_38),
.B2(n_37),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_89),
.B(n_84),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_108),
.Y(n_125)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_106),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_42),
.CI(n_36),
.CON(n_100),
.SN(n_100)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_69),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_42),
.B1(n_37),
.B2(n_18),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_112),
.B1(n_119),
.B2(n_121),
.Y(n_122)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_68),
.B(n_2),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_3),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_62),
.A2(n_24),
.B1(n_20),
.B2(n_6),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_126),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_15),
.C(n_5),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_133),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_67),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_131),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_73),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_132),
.A2(n_134),
.B(n_142),
.Y(n_184)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_56),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_146),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_56),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_137),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_138),
.B(n_140),
.Y(n_176)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_139),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_99),
.B(n_64),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_95),
.B(n_64),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_74),
.B1(n_69),
.B2(n_61),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_145),
.A2(n_94),
.B1(n_114),
.B2(n_93),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_81),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_63),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_61),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_50),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_179),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_104),
.B1(n_100),
.B2(n_119),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_164),
.B1(n_171),
.B2(n_181),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_104),
.B1(n_100),
.B2(n_119),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_103),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_167),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_150),
.B(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_173),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_123),
.A2(n_90),
.B1(n_93),
.B2(n_111),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_172),
.A2(n_178),
.B1(n_133),
.B2(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_123),
.A2(n_90),
.B1(n_93),
.B2(n_111),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_182),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_132),
.A2(n_50),
.B1(n_102),
.B2(n_108),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_142),
.B(n_117),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_130),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_195),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_135),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_192),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_134),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_154),
.C(n_157),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_131),
.C(n_137),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_198),
.C(n_202),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_191),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_124),
.B(n_145),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_152),
.C(n_134),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_197),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_136),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_127),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_124),
.B(n_125),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_203),
.B(n_180),
.C(n_173),
.D(n_154),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_102),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_147),
.B(n_143),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_106),
.B(n_96),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_172),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_139),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_209),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_164),
.B(n_168),
.C(n_158),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_223),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_160),
.C(n_183),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_186),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_178),
.Y(n_215)
);

NAND2x1_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_193),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_204),
.B1(n_192),
.B2(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_206),
.B1(n_203),
.B2(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_194),
.B(n_158),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_200),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_169),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_159),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_228),
.A2(n_212),
.B1(n_215),
.B2(n_214),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_238),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_233),
.B(n_227),
.Y(n_244)
);

FAx1_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_207),
.CI(n_198),
.CON(n_233),
.SN(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_191),
.B1(n_187),
.B2(n_188),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_194),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

OAI322xp33_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_226),
.A3(n_213),
.B1(n_219),
.B2(n_15),
.C1(n_10),
.C2(n_11),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_155),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_237),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_199),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_199),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_242),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_162),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_231),
.B(n_243),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_246),
.A2(n_247),
.B(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_228),
.A2(n_212),
.B1(n_211),
.B2(n_218),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_254),
.B1(n_229),
.B2(n_233),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_215),
.B(n_217),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_216),
.C(n_213),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_248),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_257),
.B(n_4),
.Y(n_260)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

OAI221xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.C(n_260),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_264),
.C(n_266),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_238),
.B1(n_239),
.B2(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_263),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_162),
.B1(n_156),
.B2(n_155),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_230),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_4),
.B(n_7),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_267),
.B(n_247),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_271),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_245),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_253),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_253),
.B(n_256),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_271),
.Y(n_279)
);

AO21x1_ASAP7_75t_SL g280 ( 
.A1(n_275),
.A2(n_279),
.B(n_272),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_269),
.A2(n_256),
.B1(n_8),
.B2(n_9),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_277),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_7),
.C(n_8),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_13),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_276),
.A2(n_10),
.B(n_12),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_283),
.Y(n_284)
);

OAI21x1_ASAP7_75t_L g285 ( 
.A1(n_280),
.A2(n_277),
.B(n_13),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_13),
.C(n_14),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_284),
.B(n_14),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_287),
.Y(n_290)
);


endmodule