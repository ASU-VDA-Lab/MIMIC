module fake_jpeg_15261_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_44),
.Y(n_57)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.C(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_54),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_19),
.B1(n_16),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_56),
.B1(n_63),
.B2(n_32),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_26),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_19),
.B1(n_16),
.B2(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_32),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_19),
.B1(n_31),
.B2(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_32),
.B1(n_26),
.B2(n_18),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_31),
.B1(n_25),
.B2(n_17),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_23),
.B1(n_27),
.B2(n_25),
.Y(n_87)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx2_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_74),
.A2(n_79),
.B1(n_104),
.B2(n_50),
.Y(n_117)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_78),
.B(n_93),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_80),
.B(n_102),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_88),
.B1(n_98),
.B2(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_95),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_27),
.B1(n_23),
.B2(n_15),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_89),
.B1(n_104),
.B2(n_105),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_45),
.B1(n_43),
.B2(n_40),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_86),
.A2(n_96),
.B1(n_106),
.B2(n_50),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_53),
.B1(n_50),
.B2(n_60),
.Y(n_113)
);

NAND2x1_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_25),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_25),
.C(n_54),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_27),
.B1(n_23),
.B2(n_15),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_48),
.B(n_21),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_21),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_45),
.B1(n_43),
.B2(n_35),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_45),
.B1(n_43),
.B2(n_35),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_71),
.B1(n_60),
.B2(n_67),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_49),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_13),
.B1(n_25),
.B2(n_34),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_40),
.B1(n_39),
.B2(n_34),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_129),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_115),
.B(n_93),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_78),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_123),
.B1(n_100),
.B2(n_79),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_65),
.B(n_62),
.C(n_69),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_117),
.B1(n_136),
.B2(n_91),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_71),
.B1(n_39),
.B2(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_59),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_131),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_41),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_137),
.C(n_74),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_76),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_72),
.Y(n_131)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_77),
.B(n_58),
.C(n_41),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_148),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_77),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_149),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_141),
.A2(n_151),
.B(n_153),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_106),
.B1(n_86),
.B2(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_82),
.B1(n_87),
.B2(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_82),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_111),
.B1(n_124),
.B2(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_160),
.B1(n_166),
.B2(n_132),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_102),
.B(n_101),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_80),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_109),
.A2(n_101),
.B(n_75),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_164),
.C(n_114),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_73),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_161),
.Y(n_174)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_126),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_165),
.Y(n_194)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_111),
.A2(n_107),
.B1(n_103),
.B2(n_85),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_0),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_162),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_0),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_123),
.B1(n_121),
.B2(n_132),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_30),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_72),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_115),
.A2(n_85),
.B1(n_39),
.B2(n_49),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_94),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_170),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_133),
.B(n_13),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_181),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_178),
.B(n_193),
.Y(n_220)
);

AOI22x1_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_117),
.B1(n_116),
.B2(n_125),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_183),
.B1(n_118),
.B2(n_139),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_129),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_150),
.B(n_151),
.C(n_153),
.D(n_164),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_120),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_185),
.C(n_138),
.Y(n_208)
);

OAI22x1_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_34),
.B1(n_30),
.B2(n_125),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_120),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_188),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_149),
.B(n_114),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_199),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_122),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_140),
.B(n_170),
.Y(n_219)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_144),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_142),
.A2(n_118),
.B1(n_49),
.B2(n_13),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_200),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_231)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_90),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_207),
.B1(n_223),
.B2(n_224),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_184),
.B1(n_179),
.B2(n_183),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_221),
.C(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_138),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_209),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_210),
.B(n_218),
.Y(n_247)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_222),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_234),
.B1(n_204),
.B2(n_203),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_174),
.B(n_148),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_219),
.B(n_194),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_153),
.C(n_163),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_184),
.A2(n_163),
.B1(n_162),
.B2(n_160),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_179),
.A2(n_162),
.B1(n_1),
.B2(n_2),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_227),
.A2(n_231),
.B1(n_186),
.B2(n_205),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_173),
.B(n_33),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_230),
.B(n_232),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_195),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_178),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_200),
.A2(n_33),
.B1(n_21),
.B2(n_30),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_241),
.C(n_248),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_238),
.A2(n_249),
.B1(n_251),
.B2(n_29),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_204),
.C(n_173),
.Y(n_240)
);

OAI21x1_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_224),
.B(n_212),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_198),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_250),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_233),
.A2(n_198),
.B1(n_202),
.B2(n_176),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_255),
.B1(n_232),
.B2(n_210),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_182),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_254),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_194),
.C(n_195),
.Y(n_248)
);

INVx3_ASAP7_75t_SL g251 ( 
.A(n_214),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_228),
.C(n_209),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_258),
.C(n_259),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_189),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_213),
.A2(n_189),
.B1(n_176),
.B2(n_201),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_197),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_216),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_29),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_187),
.C(n_33),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_33),
.C(n_29),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_259),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_207),
.B1(n_206),
.B2(n_225),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_262),
.A2(n_268),
.B1(n_271),
.B2(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_263),
.Y(n_296)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_264),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_234),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_277),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_243),
.A2(n_225),
.B1(n_217),
.B2(n_229),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_217),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_216),
.Y(n_270)
);

NOR2x1_ASAP7_75t_SL g271 ( 
.A(n_242),
.B(n_231),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_278),
.B1(n_245),
.B2(n_257),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_33),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_255),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_3),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_250),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_248),
.C(n_252),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_282),
.C(n_289),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_254),
.C(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_6),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_291),
.C(n_294),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_258),
.C(n_251),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_266),
.B(n_251),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_33),
.C(n_29),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_295),
.C(n_277),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_29),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_266),
.B(n_3),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_269),
.B1(n_275),
.B2(n_262),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_287),
.A2(n_264),
.B(n_279),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_298),
.A2(n_303),
.B(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_301),
.B(n_302),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_268),
.C(n_280),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_307),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_310),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_267),
.B(n_260),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_281),
.B(n_276),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_5),
.C(n_6),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_6),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_294),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_283),
.Y(n_312)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_282),
.C(n_283),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_302),
.A2(n_292),
.B1(n_291),
.B2(n_295),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_300),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_321),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_7),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_322),
.B(n_316),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_326),
.B(n_328),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_L g328 ( 
.A1(n_314),
.A2(n_303),
.B(n_309),
.C(n_304),
.D(n_11),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_12),
.B(n_8),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_312),
.A2(n_7),
.B(n_8),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_315),
.Y(n_334)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_334),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_324),
.A2(n_313),
.B(n_312),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_336),
.B(n_331),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_323),
.Y(n_336)
);

AOI321xp33_ASAP7_75t_L g340 ( 
.A1(n_337),
.A2(n_339),
.A3(n_333),
.B1(n_320),
.B2(n_11),
.C(n_12),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_329),
.Y(n_339)
);

NAND2x1p5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_7),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_338),
.B(n_10),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_12),
.B(n_317),
.Y(n_343)
);


endmodule