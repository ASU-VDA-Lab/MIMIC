module fake_jpeg_6419_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_6),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_1),
.B(n_0),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_18),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_2),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_23),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_8),
.B(n_13),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_13),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_25),
.B(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_15),
.A2(n_11),
.B1(n_7),
.B2(n_9),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_9),
.C(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_29),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_7),
.A3(n_9),
.B1(n_20),
.B2(n_22),
.C1(n_23),
.C2(n_31),
.Y(n_36)
);

AOI31xp67_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_24),
.A3(n_32),
.B(n_28),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_38),
.B(n_28),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_32),
.B(n_26),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_34),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_41),
.B(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AOI322xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_45),
.A3(n_24),
.B1(n_29),
.B2(n_34),
.C1(n_40),
.C2(n_44),
.Y(n_46)
);


endmodule