module fake_netlist_6_4746_n_104 (n_41, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_50, n_49, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_51, n_44, n_104);

input n_41;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_51;
input n_44;

output n_104;

wire n_52;
wire n_91;
wire n_88;
wire n_98;
wire n_63;
wire n_73;
wire n_68;
wire n_83;
wire n_101;
wire n_77;
wire n_92;
wire n_96;
wire n_90;
wire n_54;
wire n_102;
wire n_87;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_62;
wire n_75;
wire n_70;
wire n_67;
wire n_82;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_55;
wire n_97;
wire n_94;
wire n_58;
wire n_64;
wire n_65;
wire n_93;
wire n_80;
wire n_86;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_69;
wire n_79;
wire n_57;
wire n_53;
wire n_56;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

OA21x2_ASAP7_75t_L g58 ( 
.A1(n_0),
.A2(n_51),
.B(n_9),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_38),
.B(n_5),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_17),
.A2(n_15),
.B1(n_37),
.B2(n_40),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_32),
.B1(n_3),
.B2(n_20),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_18),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_21),
.A2(n_25),
.B1(n_12),
.B2(n_14),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_1),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_23),
.B(n_41),
.C(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_2),
.B1(n_8),
.B2(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_11),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_13),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_16),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_19),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_22),
.C(n_30),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_66),
.B(n_72),
.C(n_60),
.Y(n_83)
);

OAI21x1_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_58),
.B(n_59),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_81),
.B(n_78),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_54),
.B(n_68),
.Y(n_86)
);

OAI21x1_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_69),
.B(n_61),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_55),
.B(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_73),
.Y(n_92)
);

OR2x6_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_74),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_93),
.B(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

NAND4xp75_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_65),
.C(n_96),
.D(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_55),
.B1(n_35),
.B2(n_45),
.Y(n_103)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_34),
.B(n_49),
.Y(n_104)
);


endmodule