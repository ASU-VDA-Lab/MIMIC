module fake_jpeg_3502_n_201 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_1),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_66),
.B1(n_49),
.B2(n_57),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_57),
.B1(n_68),
.B2(n_54),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_66),
.B1(n_50),
.B2(n_64),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_82),
.B1(n_61),
.B2(n_63),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_64),
.B1(n_61),
.B2(n_49),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_65),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_88),
.C(n_87),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_106),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_103),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_107),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_57),
.B1(n_71),
.B2(n_52),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_2),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_47),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_101),
.Y(n_125)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_99),
.Y(n_116)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_62),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_54),
.B1(n_63),
.B2(n_68),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_83),
.B1(n_85),
.B2(n_55),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_93),
.B1(n_102),
.B2(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_62),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_103),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_58),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_1),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_25),
.B(n_39),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_46),
.C(n_45),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_7),
.C(n_8),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_3),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_138),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_95),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_143),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_42),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_137),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_4),
.B(n_5),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_41),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_4),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_142),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_9),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_11),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_147),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_116),
.B(n_108),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_12),
.B(n_13),
.Y(n_146)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_122),
.B(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_14),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_125),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_153),
.C(n_165),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_164),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_108),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_30),
.C(n_38),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_129),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_18),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_136),
.B(n_143),
.Y(n_168)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_160),
.B(n_157),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_145),
.B(n_139),
.Y(n_171)
);

NOR2xp67_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_150),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_28),
.B(n_36),
.C(n_34),
.D(n_33),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_179),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_27),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_165),
.C(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_184),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_182),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_154),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_176),
.B(n_152),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_167),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_170),
.B1(n_178),
.B2(n_171),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_188),
.A2(n_172),
.B(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_195),
.C(n_189),
.Y(n_196)
);

OAI321xp33_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_177),
.A3(n_184),
.B1(n_157),
.B2(n_175),
.C(n_159),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_191),
.B1(n_170),
.B2(n_21),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_32),
.B(n_40),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_19),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_20),
.Y(n_201)
);


endmodule