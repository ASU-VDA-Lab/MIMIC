module real_aes_1234_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g204 ( .A(n_0), .B(n_151), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_1), .B(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_2), .B(n_135), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_3), .B(n_153), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_4), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g142 ( .A(n_5), .Y(n_142) );
NAND2xp33_ASAP7_75t_SL g248 ( .A(n_6), .B(n_141), .Y(n_248) );
INVx1_ASAP7_75t_L g240 ( .A(n_7), .Y(n_240) );
CKINVDCx16_ASAP7_75t_R g780 ( .A(n_8), .Y(n_780) );
AND2x2_ASAP7_75t_L g129 ( .A(n_9), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g464 ( .A(n_10), .B(n_246), .Y(n_464) );
AND2x2_ASAP7_75t_L g528 ( .A(n_11), .B(n_180), .Y(n_528) );
INVx2_ASAP7_75t_L g131 ( .A(n_12), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_13), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_14), .B(n_153), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_15), .Y(n_115) );
AOI221x1_ASAP7_75t_L g243 ( .A1(n_16), .A2(n_144), .B1(n_244), .B2(n_246), .C(n_247), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_17), .B(n_135), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_18), .B(n_135), .Y(n_483) );
INVx1_ASAP7_75t_L g119 ( .A(n_19), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_20), .A2(n_66), .B1(n_771), .B2(n_772), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_20), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_21), .A2(n_90), .B1(n_135), .B2(n_184), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_22), .A2(n_144), .B(n_149), .Y(n_143) );
AOI221xp5_ASAP7_75t_SL g214 ( .A1(n_23), .A2(n_37), .B1(n_135), .B2(n_144), .C(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_24), .B(n_151), .Y(n_150) );
OR2x2_ASAP7_75t_L g132 ( .A(n_25), .B(n_89), .Y(n_132) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_25), .A2(n_89), .B(n_131), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_26), .B(n_153), .Y(n_231) );
INVxp67_ASAP7_75t_L g242 ( .A(n_27), .Y(n_242) );
AND2x2_ASAP7_75t_L g175 ( .A(n_28), .B(n_165), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_29), .A2(n_144), .B(n_203), .Y(n_202) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_30), .A2(n_246), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_31), .B(n_153), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_32), .A2(n_144), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_33), .B(n_153), .Y(n_499) );
AND2x2_ASAP7_75t_L g141 ( .A(n_34), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g145 ( .A(n_34), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g192 ( .A(n_34), .Y(n_192) );
OR2x6_ASAP7_75t_L g117 ( .A(n_35), .B(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_36), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_38), .B(n_135), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_39), .A2(n_82), .B1(n_144), .B2(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_40), .B(n_153), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_41), .B(n_135), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_42), .B(n_151), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_43), .A2(n_144), .B(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_44), .A2(n_51), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_44), .Y(n_751) );
AND2x2_ASAP7_75t_L g207 ( .A(n_45), .B(n_165), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_46), .B(n_151), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_47), .B(n_165), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_48), .B(n_135), .Y(n_507) );
INVx1_ASAP7_75t_L g138 ( .A(n_49), .Y(n_138) );
INVx1_ASAP7_75t_L g148 ( .A(n_49), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_50), .B(n_153), .Y(n_462) );
INVx1_ASAP7_75t_L g750 ( .A(n_51), .Y(n_750) );
AND2x2_ASAP7_75t_L g474 ( .A(n_52), .B(n_165), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_53), .B(n_135), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_54), .B(n_151), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_55), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_56), .B(n_151), .Y(n_498) );
AND2x2_ASAP7_75t_L g166 ( .A(n_57), .B(n_165), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_58), .B(n_135), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_59), .B(n_153), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_60), .B(n_135), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_61), .A2(n_144), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_62), .B(n_151), .Y(n_162) );
AND2x2_ASAP7_75t_SL g232 ( .A(n_63), .B(n_130), .Y(n_232) );
AND2x2_ASAP7_75t_L g489 ( .A(n_64), .B(n_130), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_65), .A2(n_144), .B(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_66), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_67), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_68), .B(n_180), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_69), .B(n_151), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_70), .B(n_151), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_71), .A2(n_92), .B1(n_144), .B2(n_190), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_72), .B(n_153), .Y(n_486) );
INVx1_ASAP7_75t_L g140 ( .A(n_73), .Y(n_140) );
INVx1_ASAP7_75t_L g146 ( .A(n_73), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_74), .B(n_151), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_75), .A2(n_144), .B(n_478), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_76), .A2(n_144), .B(n_452), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_77), .A2(n_144), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g501 ( .A(n_78), .B(n_130), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_79), .B(n_165), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_80), .B(n_135), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_81), .A2(n_84), .B1(n_135), .B2(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_85), .B(n_151), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_86), .B(n_151), .Y(n_217) );
AND2x2_ASAP7_75t_L g455 ( .A(n_87), .B(n_180), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_88), .A2(n_144), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_91), .B(n_153), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_93), .A2(n_144), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_94), .B(n_153), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_95), .B(n_135), .Y(n_206) );
INVxp67_ASAP7_75t_L g245 ( .A(n_96), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_97), .B(n_153), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_98), .A2(n_144), .B(n_229), .Y(n_228) );
BUFx2_ASAP7_75t_L g488 ( .A(n_99), .Y(n_488) );
BUFx2_ASAP7_75t_L g105 ( .A(n_100), .Y(n_105) );
AOI21xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_774), .B(n_781), .Y(n_101) );
AO21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_106), .B(n_763), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_105), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_121), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_108), .A2(n_768), .B(n_773), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
CKINVDCx11_ASAP7_75t_R g773 ( .A(n_112), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x6_ASAP7_75t_SL g440 ( .A(n_115), .B(n_117), .Y(n_440) );
OR2x6_ASAP7_75t_SL g748 ( .A(n_115), .B(n_116), .Y(n_748) );
OR2x2_ASAP7_75t_L g762 ( .A(n_115), .B(n_117), .Y(n_762) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AOI221xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_749), .B1(n_752), .B2(n_757), .C(n_758), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_439), .B1(n_441), .B2(n_746), .Y(n_122) );
INVx3_ASAP7_75t_SL g753 ( .A(n_123), .Y(n_753) );
XNOR2x1_ASAP7_75t_L g769 ( .A(n_123), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_369), .Y(n_123) );
NOR4xp25_ASAP7_75t_SL g124 ( .A(n_125), .B(n_262), .C(n_306), .D(n_333), .Y(n_124) );
OAI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_223), .B1(n_233), .B2(n_250), .C(n_252), .Y(n_125) );
AOI32xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_176), .A3(n_196), .B1(n_208), .B2(n_219), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_127), .B(n_405), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_127), .A2(n_375), .B1(n_433), .B2(n_436), .Y(n_432) );
AND2x4_ASAP7_75t_SL g127 ( .A(n_128), .B(n_156), .Y(n_127) );
INVx5_ASAP7_75t_L g222 ( .A(n_128), .Y(n_222) );
OR2x2_ASAP7_75t_L g251 ( .A(n_128), .B(n_221), .Y(n_251) );
AND2x4_ASAP7_75t_L g253 ( .A(n_128), .B(n_168), .Y(n_253) );
INVx2_ASAP7_75t_L g268 ( .A(n_128), .Y(n_268) );
OR2x2_ASAP7_75t_L g280 ( .A(n_128), .B(n_177), .Y(n_280) );
AND2x2_ASAP7_75t_L g287 ( .A(n_128), .B(n_167), .Y(n_287) );
AND2x2_ASAP7_75t_SL g329 ( .A(n_128), .B(n_210), .Y(n_329) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_128), .Y(n_386) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x4_ASAP7_75t_L g155 ( .A(n_131), .B(n_132), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_143), .B(n_155), .Y(n_133) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_141), .Y(n_135) );
INVx1_ASAP7_75t_L g249 ( .A(n_136), .Y(n_249) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
AND2x6_ASAP7_75t_L g151 ( .A(n_137), .B(n_146), .Y(n_151) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g153 ( .A(n_139), .B(n_148), .Y(n_153) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx5_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
AND2x2_ASAP7_75t_L g147 ( .A(n_142), .B(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
BUFx3_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
INVx2_ASAP7_75t_L g194 ( .A(n_146), .Y(n_194) );
AND2x4_ASAP7_75t_L g190 ( .A(n_147), .B(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_152), .B(n_154), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_151), .B(n_488), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_154), .A2(n_161), .B(n_162), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_154), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_154), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_154), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_154), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_154), .A2(n_453), .B(n_454), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_154), .A2(n_461), .B(n_462), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_154), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_154), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_154), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_154), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_154), .A2(n_525), .B(n_526), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_155), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_155), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_155), .B(n_245), .Y(n_244) );
NOR3xp33_ASAP7_75t_L g247 ( .A(n_155), .B(n_248), .C(n_249), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_155), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_155), .A2(n_507), .B(n_508), .Y(n_506) );
INVx3_ASAP7_75t_SL g281 ( .A(n_156), .Y(n_281) );
AND2x2_ASAP7_75t_L g300 ( .A(n_156), .B(n_222), .Y(n_300) );
AOI32xp33_ASAP7_75t_L g415 ( .A1(n_156), .A2(n_286), .A3(n_316), .B1(n_346), .B2(n_381), .Y(n_415) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_167), .Y(n_156) );
AND2x2_ASAP7_75t_L g255 ( .A(n_157), .B(n_177), .Y(n_255) );
OR2x2_ASAP7_75t_L g271 ( .A(n_157), .B(n_168), .Y(n_271) );
INVx1_ASAP7_75t_L g294 ( .A(n_157), .Y(n_294) );
INVx2_ASAP7_75t_L g310 ( .A(n_157), .Y(n_310) );
AND2x2_ASAP7_75t_L g347 ( .A(n_157), .B(n_210), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_157), .B(n_168), .Y(n_366) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_157), .Y(n_435) );
AO21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_164), .B(n_166), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_163), .Y(n_158) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_164), .A2(n_169), .B(n_175), .Y(n_168) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_164), .A2(n_169), .B(n_175), .Y(n_221) );
AOI21x1_ASAP7_75t_L g521 ( .A1(n_164), .A2(n_522), .B(n_528), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_165), .Y(n_164) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_165), .A2(n_214), .B(n_218), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_165), .A2(n_450), .B(n_451), .Y(n_449) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_165), .A2(n_468), .B(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g402 ( .A(n_168), .B(n_177), .Y(n_402) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_168), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_174), .Y(n_169) );
OR2x2_ASAP7_75t_L g250 ( .A(n_176), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g256 ( .A(n_176), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g269 ( .A(n_176), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g431 ( .A(n_176), .B(n_300), .Y(n_431) );
BUFx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g360 ( .A(n_177), .B(n_310), .Y(n_360) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_178), .Y(n_210) );
AOI21x1_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_195), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_180), .A2(n_227), .B(n_228), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_180), .A2(n_483), .B(n_484), .Y(n_482) );
BUFx4f_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx3_ASAP7_75t_L g200 ( .A(n_181), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_189), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_184), .A2(n_190), .B1(n_239), .B2(n_241), .Y(n_238) );
AND2x4_ASAP7_75t_L g184 ( .A(n_185), .B(n_188), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2x1p5_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_196), .B(n_327), .Y(n_429) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_197), .B(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g212 ( .A(n_198), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g234 ( .A(n_198), .Y(n_234) );
AND2x2_ASAP7_75t_L g260 ( .A(n_198), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_198), .B(n_236), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_198), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g318 ( .A(n_198), .Y(n_318) );
OR2x2_ASAP7_75t_L g337 ( .A(n_198), .B(n_264), .Y(n_337) );
INVx1_ASAP7_75t_L g344 ( .A(n_198), .Y(n_344) );
NOR2xp33_ASAP7_75t_R g396 ( .A(n_198), .B(n_225), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_198), .B(n_237), .Y(n_400) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AOI21x1_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_207), .Y(n_199) );
INVx4_ASAP7_75t_L g246 ( .A(n_200), .Y(n_246) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_200), .A2(n_458), .B(n_464), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_206), .Y(n_201) );
AOI32xp33_ASAP7_75t_L g423 ( .A1(n_208), .A2(n_259), .A3(n_424), .B1(n_425), .B2(n_426), .Y(n_423) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g290 ( .A(n_210), .Y(n_290) );
AND2x4_ASAP7_75t_L g309 ( .A(n_210), .B(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_210), .B(n_281), .Y(n_338) );
OR2x2_ASAP7_75t_L g392 ( .A(n_210), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g350 ( .A(n_211), .B(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g408 ( .A(n_211), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_212), .B(n_225), .Y(n_374) );
AND2x2_ASAP7_75t_L g411 ( .A(n_212), .B(n_377), .Y(n_411) );
INVx2_ASAP7_75t_L g261 ( .A(n_213), .Y(n_261) );
INVx2_ASAP7_75t_L g264 ( .A(n_213), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_213), .B(n_225), .Y(n_284) );
INVx1_ASAP7_75t_L g315 ( .A(n_213), .Y(n_315) );
OR2x2_ASAP7_75t_L g341 ( .A(n_213), .B(n_225), .Y(n_341) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_213), .Y(n_393) );
BUFx3_ASAP7_75t_L g422 ( .A(n_213), .Y(n_422) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g291 ( .A(n_220), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_220), .B(n_309), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_220), .B(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_221), .B(n_294), .Y(n_293) );
OAI21xp33_ASAP7_75t_L g323 ( .A1(n_221), .A2(n_290), .B(n_308), .Y(n_323) );
OAI32xp33_ASAP7_75t_L g345 ( .A1(n_222), .A2(n_346), .A3(n_348), .B1(n_350), .B2(n_352), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_222), .B(n_309), .Y(n_418) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g351 ( .A(n_224), .Y(n_351) );
NOR2x1p5_ASAP7_75t_L g421 ( .A(n_224), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_L g235 ( .A(n_225), .B(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_SL g259 ( .A(n_225), .B(n_237), .Y(n_259) );
OR2x2_ASAP7_75t_L g263 ( .A(n_225), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
AND2x2_ASAP7_75t_L g316 ( .A(n_225), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g327 ( .A(n_225), .B(n_237), .Y(n_327) );
OR2x2_ASAP7_75t_L g389 ( .A(n_225), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g406 ( .A(n_225), .B(n_337), .Y(n_406) );
INVx1_ASAP7_75t_L g438 ( .A(n_225), .Y(n_438) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_232), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_234), .B(n_315), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_235), .B(n_349), .Y(n_348) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_235), .A2(n_354), .B1(n_359), .B2(n_361), .C1(n_364), .C2(n_367), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_235), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g381 ( .A(n_235), .B(n_260), .Y(n_381) );
AND2x2_ASAP7_75t_L g343 ( .A(n_236), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g358 ( .A(n_236), .B(n_263), .Y(n_358) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_237), .B(n_264), .Y(n_296) );
AND2x4_ASAP7_75t_L g317 ( .A(n_237), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g377 ( .A(n_237), .B(n_298), .Y(n_377) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_243), .Y(n_237) );
INVx3_ASAP7_75t_L g494 ( .A(n_246), .Y(n_494) );
INVx1_ASAP7_75t_SL g257 ( .A(n_251), .Y(n_257) );
NAND2xp33_ASAP7_75t_SL g426 ( .A(n_251), .B(n_281), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_256), .C(n_258), .Y(n_252) );
INVx2_ASAP7_75t_SL g303 ( .A(n_253), .Y(n_303) );
AND2x2_ASAP7_75t_L g307 ( .A(n_254), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_255), .B(n_303), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_255), .A2(n_293), .B(n_329), .C(n_330), .Y(n_328) );
AND2x2_ASAP7_75t_L g405 ( .A(n_255), .B(n_386), .Y(n_405) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x4_ASAP7_75t_L g304 ( .A(n_259), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g409 ( .A(n_259), .Y(n_409) );
OAI211xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B(n_272), .C(n_299), .Y(n_262) );
INVx2_ASAP7_75t_L g274 ( .A(n_263), .Y(n_274) );
OR2x2_ASAP7_75t_L g321 ( .A(n_263), .B(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_264), .Y(n_305) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_267), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g359 ( .A(n_267), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_267), .B(n_347), .Y(n_413) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AOI222xp33_ASAP7_75t_L g371 ( .A1(n_269), .A2(n_372), .B1(n_373), .B2(n_375), .C1(n_378), .C2(n_381), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_270), .A2(n_335), .B1(n_338), .B2(n_339), .C(n_345), .Y(n_334) );
AND2x2_ASAP7_75t_L g372 ( .A(n_270), .B(n_329), .Y(n_372) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp33_ASAP7_75t_SL g285 ( .A(n_271), .B(n_286), .Y(n_285) );
AOI221x1_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_277), .B1(n_282), .B2(n_285), .C(n_288), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_L g425 ( .A(n_275), .B(n_363), .Y(n_425) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g283 ( .A(n_276), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
OAI32xp33_ASAP7_75t_L g391 ( .A1(n_281), .A2(n_322), .A3(n_392), .B1(n_394), .B2(n_398), .Y(n_391) );
OAI21xp33_ASAP7_75t_SL g410 ( .A1(n_282), .A2(n_411), .B(n_412), .Y(n_410) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AOI21xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_292), .B(n_295), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
OR2x2_ASAP7_75t_L g292 ( .A(n_290), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g365 ( .A(n_290), .B(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_294), .A2(n_320), .B1(n_323), .B2(n_324), .C(n_328), .Y(n_319) );
INVx1_ASAP7_75t_L g395 ( .A(n_294), .Y(n_395) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_294), .Y(n_401) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
OAI21xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B(n_304), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_303), .B(n_368), .Y(n_367) );
OAI21xp5_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_311), .B(n_319), .Y(n_306) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_310), .Y(n_380) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_313), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVxp67_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g332 ( .A(n_315), .Y(n_332) );
INVx1_ASAP7_75t_L g322 ( .A(n_317), .Y(n_322) );
AND2x2_ASAP7_75t_SL g331 ( .A(n_317), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_317), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_317), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g336 ( .A(n_327), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_332), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_334), .B(n_353), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g349 ( .A(n_337), .Y(n_349) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_SL g363 ( .A(n_341), .Y(n_363) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_343), .B(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_344), .Y(n_357) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_355), .B(n_358), .Y(n_354) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g368 ( .A(n_360), .Y(n_368) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g387 ( .A(n_366), .Y(n_387) );
NOR4xp25_ASAP7_75t_L g369 ( .A(n_370), .B(n_403), .C(n_414), .D(n_427), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_382), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_L g382 ( .A1(n_372), .A2(n_383), .B(n_388), .C(n_391), .Y(n_382) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_387), .Y(n_384) );
OAI211xp5_ASAP7_75t_L g394 ( .A1(n_385), .A2(n_395), .B(n_396), .C(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
OAI21xp33_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_401), .B(n_402), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_402), .B(n_434), .Y(n_433) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_406), .B1(n_407), .B2(n_408), .C(n_410), .Y(n_403) );
INVx1_ASAP7_75t_SL g407 ( .A(n_405), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND3xp33_ASAP7_75t_SL g414 ( .A(n_415), .B(n_416), .C(n_423), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B(n_432), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp33_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
CKINVDCx11_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_440), .Y(n_754) );
INVx2_ASAP7_75t_SL g755 ( .A(n_441), .Y(n_755) );
AND2x4_ASAP7_75t_L g441 ( .A(n_442), .B(n_671), .Y(n_441) );
NOR2xp67_ASAP7_75t_L g442 ( .A(n_443), .B(n_590), .Y(n_442) );
NAND5xp2_ASAP7_75t_L g443 ( .A(n_444), .B(n_534), .C(n_544), .D(n_561), .E(n_577), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_470), .B1(n_512), .B2(n_516), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_456), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g518 ( .A(n_448), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g536 ( .A(n_448), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g557 ( .A(n_448), .B(n_558), .Y(n_557) );
INVx4_ASAP7_75t_L g571 ( .A(n_448), .Y(n_571) );
AND2x2_ASAP7_75t_L g580 ( .A(n_448), .B(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_SL g602 ( .A(n_448), .B(n_520), .Y(n_602) );
BUFx2_ASAP7_75t_L g645 ( .A(n_448), .Y(n_645) );
AND2x2_ASAP7_75t_L g660 ( .A(n_448), .B(n_457), .Y(n_660) );
OR2x2_ASAP7_75t_L g692 ( .A(n_448), .B(n_693), .Y(n_692) );
NOR4xp25_ASAP7_75t_L g741 ( .A(n_448), .B(n_742), .C(n_743), .D(n_744), .Y(n_741) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_455), .Y(n_448) );
AOI31xp33_ASAP7_75t_L g609 ( .A1(n_456), .A2(n_610), .A3(n_612), .B(n_614), .Y(n_609) );
INVx2_ASAP7_75t_SL g726 ( .A(n_456), .Y(n_726) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_465), .Y(n_456) );
INVx2_ASAP7_75t_L g533 ( .A(n_457), .Y(n_533) );
AND2x2_ASAP7_75t_L g537 ( .A(n_457), .B(n_521), .Y(n_537) );
INVx2_ASAP7_75t_L g560 ( .A(n_457), .Y(n_560) );
AND2x2_ASAP7_75t_L g579 ( .A(n_457), .B(n_520), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_463), .Y(n_458) );
AND2x2_ASAP7_75t_L g531 ( .A(n_465), .B(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g538 ( .A(n_465), .Y(n_538) );
INVx2_ASAP7_75t_L g556 ( .A(n_465), .Y(n_556) );
AND2x2_ASAP7_75t_L g611 ( .A(n_465), .B(n_571), .Y(n_611) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AND2x4_ASAP7_75t_L g582 ( .A(n_466), .B(n_467), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_502), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_490), .Y(n_471) );
OR2x2_ASAP7_75t_L g512 ( .A(n_472), .B(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g663 ( .A(n_472), .Y(n_663) );
OR2x2_ASAP7_75t_L g711 ( .A(n_472), .B(n_712), .Y(n_711) );
NAND2x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_481), .Y(n_472) );
OR2x2_ASAP7_75t_SL g503 ( .A(n_473), .B(n_504), .Y(n_503) );
INVx4_ASAP7_75t_L g541 ( .A(n_473), .Y(n_541) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_473), .Y(n_585) );
INVx2_ASAP7_75t_L g593 ( .A(n_473), .Y(n_593) );
OR2x2_ASAP7_75t_L g628 ( .A(n_473), .B(n_492), .Y(n_628) );
AND2x2_ASAP7_75t_L g740 ( .A(n_473), .B(n_595), .Y(n_740) );
AND2x2_ASAP7_75t_L g745 ( .A(n_473), .B(n_505), .Y(n_745) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
OR2x2_ASAP7_75t_L g504 ( .A(n_481), .B(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g569 ( .A(n_481), .B(n_491), .Y(n_569) );
OR2x2_ASAP7_75t_L g576 ( .A(n_481), .B(n_541), .Y(n_576) );
NOR2x1_ASAP7_75t_SL g595 ( .A(n_481), .B(n_515), .Y(n_595) );
BUFx2_ASAP7_75t_L g627 ( .A(n_481), .Y(n_627) );
AND2x2_ASAP7_75t_L g636 ( .A(n_481), .B(n_541), .Y(n_636) );
AND2x2_ASAP7_75t_L g669 ( .A(n_481), .B(n_589), .Y(n_669) );
INVx2_ASAP7_75t_SL g678 ( .A(n_481), .Y(n_678) );
AND2x2_ASAP7_75t_L g681 ( .A(n_481), .B(n_492), .Y(n_681) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_489), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_490), .B(n_546), .C(n_631), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_490), .B(n_593), .Y(n_696) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_491), .B(n_678), .Y(n_699) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_492), .Y(n_543) );
AND2x2_ASAP7_75t_L g587 ( .A(n_492), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g652 ( .A(n_492), .B(n_653), .Y(n_652) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_501), .Y(n_493) );
AO21x1_ASAP7_75t_SL g515 ( .A1(n_494), .A2(n_495), .B(n_501), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_500), .Y(n_495) );
AND2x4_ASAP7_75t_L g547 ( .A(n_502), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g683 ( .A(n_504), .B(n_628), .Y(n_683) );
AND2x2_ASAP7_75t_L g514 ( .A(n_505), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g551 ( .A(n_505), .Y(n_551) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_505), .Y(n_568) );
INVx2_ASAP7_75t_L g589 ( .A(n_505), .Y(n_589) );
INVx1_ASAP7_75t_L g653 ( .A(n_505), .Y(n_653) );
INVx2_ASAP7_75t_L g735 ( .A(n_512), .Y(n_735) );
OR2x2_ASAP7_75t_L g599 ( .A(n_513), .B(n_576), .Y(n_599) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g739 ( .A(n_514), .B(n_636), .Y(n_739) );
AND2x2_ASAP7_75t_L g632 ( .A(n_515), .B(n_589), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_529), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_518), .A2(n_646), .B1(n_663), .B2(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g559 ( .A(n_520), .Y(n_559) );
AND2x2_ASAP7_75t_L g613 ( .A(n_520), .B(n_533), .Y(n_613) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_520), .Y(n_640) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_521), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
INVxp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_531), .B(n_645), .Y(n_644) );
OAI32xp33_ASAP7_75t_L g661 ( .A1(n_531), .A2(n_662), .A3(n_664), .B1(n_665), .B2(n_667), .Y(n_661) );
BUFx2_ASAP7_75t_L g546 ( .A(n_532), .Y(n_546) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g688 ( .A(n_533), .B(n_582), .Y(n_688) );
OR4x1_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .C(n_539), .D(n_542), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_535), .A2(n_626), .B1(n_720), .B2(n_721), .Y(n_719) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_536), .Y(n_728) );
AND2x2_ASAP7_75t_L g570 ( .A(n_537), .B(n_571), .Y(n_570) );
BUFx2_ASAP7_75t_L g650 ( .A(n_537), .Y(n_650) );
INVx1_ASAP7_75t_L g666 ( .A(n_537), .Y(n_666) );
INVx1_ASAP7_75t_L g701 ( .A(n_537), .Y(n_701) );
OR2x2_ASAP7_75t_L g658 ( .A(n_538), .B(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g702 ( .A(n_538), .B(n_703), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_539), .A2(n_576), .B1(n_620), .B2(n_639), .Y(n_641) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g685 ( .A(n_540), .B(n_594), .Y(n_685) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx2_ASAP7_75t_L g552 ( .A(n_541), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g567 ( .A(n_541), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g548 ( .A(n_542), .Y(n_548) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_542), .B(n_546), .C(n_627), .D(n_639), .Y(n_675) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g712 ( .A(n_543), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B1(n_549), .B2(n_553), .Y(n_544) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_545), .A2(n_546), .B1(n_696), .B2(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVxp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx3_ASAP7_75t_L g574 ( .A(n_551), .Y(n_574) );
AOI32xp33_ASAP7_75t_L g690 ( .A1(n_551), .A2(n_691), .A3(n_695), .B1(n_700), .B2(n_704), .Y(n_690) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_554), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g649 ( .A(n_554), .B(n_650), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_554), .A2(n_562), .B1(n_674), .B2(n_679), .C(n_682), .Y(n_673) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g606 ( .A(n_555), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g721 ( .A(n_555), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_556), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g563 ( .A(n_558), .Y(n_563) );
AND2x2_ASAP7_75t_L g581 ( .A(n_558), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_SL g621 ( .A(n_559), .Y(n_621) );
INVx1_ASAP7_75t_L g605 ( .A(n_560), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_564), .B1(n_570), .B2(n_572), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g707 ( .A(n_563), .B(n_637), .Y(n_707) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g647 ( .A(n_566), .Y(n_647) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
AND2x2_ASAP7_75t_L g578 ( .A(n_571), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_571), .B(n_608), .Y(n_607) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_571), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_571), .B(n_613), .Y(n_734) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_572), .A2(n_732), .B1(n_733), .B2(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
OR2x2_ASAP7_75t_L g614 ( .A(n_574), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g624 ( .A(n_574), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_574), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_574), .B(n_678), .Y(n_677) );
AND2x4_ASAP7_75t_SL g679 ( .A(n_574), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g655 ( .A(n_576), .B(n_656), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_580), .B(n_583), .Y(n_577) );
INVx1_ASAP7_75t_L g597 ( .A(n_579), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_580), .A2(n_617), .B1(n_624), .B2(n_629), .Y(n_616) );
INVx3_ASAP7_75t_L g619 ( .A(n_582), .Y(n_619) );
INVx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OAI32xp33_ASAP7_75t_SL g674 ( .A1(n_585), .A2(n_645), .A3(n_675), .B1(n_676), .B2(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g594 ( .A(n_588), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND4xp25_ASAP7_75t_SL g590 ( .A(n_591), .B(n_616), .C(n_633), .D(n_648), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_596), .B1(n_598), .B2(n_600), .C(n_609), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx2_ASAP7_75t_L g631 ( .A(n_593), .Y(n_631) );
AND2x2_ASAP7_75t_L g680 ( .A(n_593), .B(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_593), .B(n_632), .Y(n_718) );
AND2x2_ASAP7_75t_L g729 ( .A(n_593), .B(n_652), .Y(n_729) );
INVx2_ASAP7_75t_L g615 ( .A(n_595), .Y(n_615) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .B(n_606), .Y(n_600) );
AND2x2_ASAP7_75t_L g732 ( .A(n_601), .B(n_603), .Y(n_732) );
INVx2_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_602), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g709 ( .A(n_607), .Y(n_709) );
INVx1_ASAP7_75t_L g694 ( .A(n_608), .Y(n_694) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_611), .B(n_666), .Y(n_665) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_612), .B(n_619), .Y(n_623) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g722 ( .A(n_613), .Y(n_722) );
INVx1_ASAP7_75t_L g704 ( .A(n_615), .Y(n_704) );
OR2x2_ASAP7_75t_L g720 ( .A(n_615), .B(n_631), .Y(n_720) );
NAND2xp33_ASAP7_75t_SL g617 ( .A(n_618), .B(n_622), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_L g637 ( .A(n_619), .Y(n_637) );
AND2x2_ASAP7_75t_L g642 ( .A(n_619), .B(n_632), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_619), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g716 ( .A(n_620), .Y(n_716) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_625), .A2(n_706), .B1(n_708), .B2(n_710), .Y(n_705) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g670 ( .A(n_628), .Y(n_670) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g656 ( .A(n_632), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .A3(n_638), .B1(n_641), .B2(n_642), .C1(n_643), .C2(n_646), .Y(n_633) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_634), .A2(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g651 ( .A(n_636), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g708 ( .A(n_637), .B(n_709), .Y(n_708) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_644), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g664 ( .A(n_645), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_645), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B1(n_654), .B2(n_657), .C(n_661), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_650), .A2(n_737), .B1(n_739), .B2(n_740), .C(n_741), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_652), .B(n_663), .Y(n_662) );
BUFx2_ASAP7_75t_L g703 ( .A(n_653), .Y(n_703) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g727 ( .A1(n_657), .A2(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp33_ASAP7_75t_SL g737 ( .A(n_666), .B(n_738), .Y(n_737) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
NOR4xp75_ASAP7_75t_L g671 ( .A(n_672), .B(n_689), .C(n_713), .D(n_730), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_684), .Y(n_672) );
INVx1_ASAP7_75t_L g743 ( .A(n_681), .Y(n_743) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g715 ( .A(n_688), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g742 ( .A(n_688), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_690), .B(n_705), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_SL g738 ( .A(n_709), .Y(n_738) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND3x1_ASAP7_75t_L g713 ( .A(n_714), .B(n_723), .C(n_727), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B(n_719), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_736), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_747), .Y(n_756) );
CKINVDCx11_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g757 ( .A(n_749), .Y(n_757) );
OAI22x1_ASAP7_75t_SL g752 ( .A1(n_753), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx2_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_761), .B(n_778), .Y(n_777) );
INVx3_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_767), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g783 ( .A(n_775), .Y(n_783) );
INVx3_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
endmodule