module fake_netlist_6_2920_n_1350 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_105, n_227, n_132, n_102, n_204, n_261, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_41, n_134, n_273, n_95, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1350);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_41;
input n_134;
input n_273;
input n_95;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1350;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_1332;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_482;
wire n_934;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_859;
wire n_570;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_62),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_217),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_47),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_189),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_180),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_183),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_231),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_120),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_184),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_293),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_95),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_61),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_251),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_236),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_75),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_84),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_252),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_90),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_112),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_209),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_82),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_304),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_163),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_69),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_56),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_101),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_169),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_155),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_188),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_258),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_99),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_211),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_195),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_162),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_11),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_270),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_25),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_303),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_84),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_253),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_157),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_45),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_59),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_140),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_172),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_192),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_91),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g363 ( 
.A(n_168),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_171),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_44),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_266),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_28),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_170),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_254),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_263),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_104),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_144),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_69),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_62),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_80),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_237),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_182),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_296),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_7),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_299),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_265),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_17),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_176),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_165),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_135),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_93),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_45),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_30),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_92),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_194),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_70),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_60),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_119),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_77),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_178),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_282),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_285),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_158),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_161),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_92),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_152),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_235),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_36),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_294),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_91),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_216),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_255),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_37),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_115),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_190),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_43),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_103),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_256),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_116),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_159),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_250),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_136),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_207),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_23),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_109),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_89),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_43),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_259),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_21),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_244),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_227),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_226),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_47),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_240),
.Y(n_429)
);

BUFx10_ASAP7_75t_L g430 ( 
.A(n_286),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_262),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_249),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_41),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_257),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_151),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_123),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_133),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_279),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_203),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_52),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_283),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_64),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_153),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_191),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_204),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_185),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_292),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_137),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_60),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_96),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_15),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_26),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_143),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_56),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_241),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_243),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_132),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_181),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_93),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_160),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_79),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_86),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_219),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_228),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_290),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_139),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_187),
.Y(n_467)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_233),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_210),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_306),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_221),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_23),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_287),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_0),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_65),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_201),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_234),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_230),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_59),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_277),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_14),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_29),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_288),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_63),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_17),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_205),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_68),
.Y(n_487)
);

CKINVDCx14_ASAP7_75t_R g488 ( 
.A(n_215),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_82),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_238),
.Y(n_490)
);

BUFx10_ASAP7_75t_L g491 ( 
.A(n_229),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_232),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_224),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_71),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g495 ( 
.A(n_111),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_117),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_33),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_53),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_177),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_271),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_90),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_1),
.Y(n_502)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_51),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_245),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_124),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_1),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_193),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_122),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_35),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_48),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_106),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_154),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_200),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_301),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_208),
.Y(n_515)
);

BUFx10_ASAP7_75t_L g516 ( 
.A(n_305),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_127),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_46),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_206),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_75),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_0),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_134),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_298),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_87),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_4),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_7),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_239),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_278),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_218),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_300),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_242),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_54),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_98),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_150),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_400),
.B(n_472),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_312),
.B(n_2),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_314),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_346),
.B(n_3),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_314),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_503),
.B(n_3),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_400),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_356),
.B(n_4),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_400),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_438),
.B(n_5),
.Y(n_545)
);

BUFx8_ASAP7_75t_SL g546 ( 
.A(n_328),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_314),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_315),
.B(n_5),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_400),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_426),
.B(n_6),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_360),
.B(n_6),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_436),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_472),
.Y(n_553)
);

BUFx12f_ASAP7_75t_L g554 ( 
.A(n_532),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_472),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_360),
.B(n_8),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_472),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_436),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_436),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_374),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_430),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_383),
.B(n_8),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_382),
.Y(n_564)
);

BUFx8_ASAP7_75t_L g565 ( 
.A(n_485),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_430),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_356),
.B(n_9),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_443),
.B(n_9),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_492),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_492),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_443),
.B(n_10),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_485),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_492),
.B(n_94),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_507),
.Y(n_575)
);

CKINVDCx6p67_ASAP7_75t_R g576 ( 
.A(n_532),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_507),
.Y(n_577)
);

BUFx12f_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_507),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_485),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_491),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_383),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_447),
.B(n_11),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_507),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_513),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_393),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_513),
.Y(n_587)
);

BUFx12f_ASAP7_75t_L g588 ( 
.A(n_516),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_428),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_485),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_513),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_428),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_393),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_363),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_534),
.B(n_447),
.Y(n_595)
);

BUFx12f_ASAP7_75t_L g596 ( 
.A(n_516),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_465),
.B(n_12),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_469),
.B(n_12),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_469),
.B(n_471),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_459),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_534),
.B(n_13),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_363),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_363),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_459),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_520),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_527),
.B(n_97),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_471),
.B(n_13),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_519),
.B(n_14),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_519),
.B(n_15),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_530),
.B(n_16),
.Y(n_610)
);

BUFx12f_ASAP7_75t_L g611 ( 
.A(n_516),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_530),
.B(n_16),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_450),
.B(n_466),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_506),
.Y(n_614)
);

BUFx8_ASAP7_75t_L g615 ( 
.A(n_506),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_450),
.B(n_18),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_465),
.B(n_18),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_520),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_316),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_468),
.B(n_19),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_466),
.B(n_19),
.Y(n_621)
);

BUFx12f_ASAP7_75t_L g622 ( 
.A(n_310),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_351),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_461),
.B(n_20),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_324),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_527),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_363),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_311),
.B(n_20),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_407),
.B(n_21),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_527),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_329),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_318),
.B(n_22),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_527),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_320),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_410),
.B(n_24),
.Y(n_635)
);

XNOR2x1_ASAP7_75t_L g636 ( 
.A(n_334),
.B(n_24),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_353),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_325),
.B(n_25),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_362),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_365),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_330),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_441),
.B(n_26),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_480),
.B(n_27),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_479),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_317),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_363),
.Y(n_646)
);

BUFx8_ASAP7_75t_L g647 ( 
.A(n_387),
.Y(n_647)
);

BUFx12f_ASAP7_75t_L g648 ( 
.A(n_337),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_377),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_397),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_335),
.B(n_27),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_389),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_336),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_468),
.B(n_28),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_339),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_363),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_344),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_488),
.B(n_29),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_345),
.B(n_30),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_349),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_413),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_347),
.B(n_31),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_391),
.Y(n_663)
);

BUFx12f_ASAP7_75t_L g664 ( 
.A(n_357),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_408),
.B(n_31),
.Y(n_665)
);

CKINVDCx11_ASAP7_75t_R g666 ( 
.A(n_331),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_488),
.B(n_32),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_338),
.B(n_32),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_490),
.B(n_33),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_348),
.B(n_34),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_495),
.B(n_34),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_495),
.B(n_35),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_500),
.B(n_36),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_355),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_379),
.B(n_38),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_359),
.B(n_39),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_368),
.B(n_39),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_319),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_413),
.B(n_40),
.Y(n_679)
);

BUFx12f_ASAP7_75t_L g680 ( 
.A(n_358),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_413),
.B(n_40),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_411),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_413),
.B(n_41),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_378),
.B(n_42),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_380),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_386),
.B(n_42),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_388),
.B(n_44),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_413),
.B(n_46),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_619),
.B(n_381),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_542),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_549),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_597),
.A2(n_620),
.B1(n_654),
.B2(n_617),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_SL g693 ( 
.A1(n_623),
.A2(n_373),
.B1(n_375),
.B2(n_367),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_667),
.A2(n_321),
.B1(n_333),
.B2(n_313),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_SL g695 ( 
.A1(n_536),
.A2(n_403),
.B1(n_405),
.B2(n_392),
.Y(n_695)
);

AO22x2_ASAP7_75t_L g696 ( 
.A1(n_551),
.A2(n_422),
.B1(n_424),
.B2(n_421),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_622),
.B(n_433),
.Y(n_697)
);

AO22x2_ASAP7_75t_L g698 ( 
.A1(n_551),
.A2(n_474),
.B1(n_482),
.B2(n_442),
.Y(n_698)
);

AO22x2_ASAP7_75t_L g699 ( 
.A1(n_556),
.A2(n_487),
.B1(n_489),
.B2(n_484),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_671),
.A2(n_350),
.B1(n_366),
.B2(n_342),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_672),
.A2(n_384),
.B1(n_414),
.B2(n_369),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_649),
.B(n_522),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_580),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_549),
.Y(n_704)
);

NAND3x1_ASAP7_75t_L g705 ( 
.A(n_538),
.B(n_409),
.C(n_395),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_SL g706 ( 
.A1(n_541),
.A2(n_449),
.B1(n_451),
.B2(n_440),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_540),
.B(n_322),
.Y(n_707)
);

AO22x2_ASAP7_75t_L g708 ( 
.A1(n_556),
.A2(n_510),
.B1(n_416),
.B2(n_417),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_590),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_590),
.Y(n_710)
);

OA22x2_ASAP7_75t_L g711 ( 
.A1(n_623),
.A2(n_592),
.B1(n_605),
.B2(n_589),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_648),
.B(n_664),
.Y(n_712)
);

NAND3x1_ASAP7_75t_L g713 ( 
.A(n_545),
.B(n_431),
.C(n_412),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_544),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_L g715 ( 
.A1(n_668),
.A2(n_454),
.B1(n_462),
.B2(n_452),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_649),
.B(n_650),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_649),
.B(n_323),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_SL g718 ( 
.A1(n_668),
.A2(n_494),
.B1(n_497),
.B2(n_481),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_658),
.A2(n_529),
.B1(n_455),
.B2(n_501),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_SL g720 ( 
.A1(n_548),
.A2(n_419),
.B1(n_475),
.B2(n_394),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_567),
.Y(n_721)
);

AO22x2_ASAP7_75t_L g722 ( 
.A1(n_563),
.A2(n_457),
.B1(n_463),
.B2(n_448),
.Y(n_722)
);

AO22x2_ASAP7_75t_L g723 ( 
.A1(n_563),
.A2(n_477),
.B1(n_478),
.B2(n_476),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_547),
.Y(n_724)
);

AO22x2_ASAP7_75t_L g725 ( 
.A1(n_621),
.A2(n_499),
.B1(n_514),
.B2(n_486),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_650),
.B(n_326),
.Y(n_726)
);

NAND3x1_ASAP7_75t_L g727 ( 
.A(n_550),
.B(n_531),
.C(n_528),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_678),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_561),
.A2(n_502),
.B1(n_509),
.B2(n_498),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_547),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_650),
.B(n_327),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_629),
.A2(n_521),
.B1(n_524),
.B2(n_518),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_SL g733 ( 
.A1(n_686),
.A2(n_526),
.B1(n_525),
.B2(n_340),
.Y(n_733)
);

OR2x6_ASAP7_75t_L g734 ( 
.A(n_680),
.B(n_48),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_544),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_553),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_635),
.A2(n_341),
.B1(n_343),
.B2(n_332),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_642),
.A2(n_354),
.B1(n_361),
.B2(n_352),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_SL g739 ( 
.A1(n_687),
.A2(n_370),
.B1(n_371),
.B2(n_364),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_559),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_SL g741 ( 
.A1(n_616),
.A2(n_376),
.B1(n_385),
.B2(n_372),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_562),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_643),
.A2(n_396),
.B1(n_398),
.B2(n_390),
.Y(n_743)
);

AO22x2_ASAP7_75t_L g744 ( 
.A1(n_621),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_559),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_SL g746 ( 
.A(n_675),
.B(n_399),
.Y(n_746)
);

AND2x2_ASAP7_75t_SL g747 ( 
.A(n_669),
.B(n_49),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_660),
.B(n_401),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_666),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_673),
.A2(n_404),
.B1(n_406),
.B2(n_402),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_582),
.B(n_415),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_586),
.B(n_418),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_564),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_624),
.A2(n_423),
.B1(n_425),
.B2(n_420),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_581),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_593),
.B(n_427),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_559),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_613),
.B(n_429),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_613),
.B(n_432),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_553),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_SL g761 ( 
.A1(n_624),
.A2(n_533),
.B1(n_523),
.B2(n_517),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_555),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_665),
.A2(n_515),
.B1(n_512),
.B2(n_511),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_588),
.A2(n_508),
.B1(n_505),
.B2(n_504),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_554),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_L g766 ( 
.A1(n_543),
.A2(n_496),
.B1(n_493),
.B2(n_483),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_555),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_596),
.A2(n_473),
.B1(n_470),
.B2(n_467),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_546),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_645),
.B(n_464),
.Y(n_770)
);

OAI22xp33_ASAP7_75t_L g771 ( 
.A1(n_543),
.A2(n_460),
.B1(n_458),
.B2(n_456),
.Y(n_771)
);

OA22x2_ASAP7_75t_L g772 ( 
.A1(n_631),
.A2(n_453),
.B1(n_446),
.B2(n_445),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_583),
.B(n_610),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_644),
.B(n_434),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_611),
.A2(n_578),
.B1(n_576),
.B2(n_569),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_583),
.A2(n_444),
.B1(n_439),
.B2(n_437),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_636),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_615),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_566),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_557),
.Y(n_780)
);

OAI22xp33_ASAP7_75t_L g781 ( 
.A1(n_610),
.A2(n_435),
.B1(n_57),
.B2(n_58),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_566),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_557),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_644),
.B(n_100),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_573),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_572),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_SL g787 ( 
.A1(n_665),
.A2(n_55),
.B1(n_61),
.B2(n_63),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_L g788 ( 
.A1(n_568),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_598),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_773),
.B(n_594),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_753),
.B(n_732),
.Y(n_791)
);

AND2x6_ASAP7_75t_L g792 ( 
.A(n_784),
.B(n_628),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_724),
.Y(n_793)
);

XNOR2x2_ASAP7_75t_L g794 ( 
.A(n_777),
.B(n_608),
.Y(n_794)
);

INVxp67_ASAP7_75t_SL g795 ( 
.A(n_714),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_730),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_740),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_757),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_719),
.B(n_618),
.Y(n_799)
);

XNOR2x2_ASAP7_75t_L g800 ( 
.A(n_777),
.B(n_612),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_779),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_751),
.B(n_752),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_756),
.B(n_652),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_782),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_689),
.B(n_595),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_691),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_691),
.Y(n_807)
);

XNOR2xp5_ASAP7_75t_L g808 ( 
.A(n_749),
.B(n_628),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_709),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_770),
.B(n_599),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_709),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_710),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_710),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_715),
.B(n_601),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_692),
.A2(n_535),
.B(n_607),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_767),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_754),
.B(n_609),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_780),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_714),
.B(n_602),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_748),
.Y(n_820)
);

NOR2xp67_ASAP7_75t_L g821 ( 
.A(n_737),
.B(n_539),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_745),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_728),
.B(n_632),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_783),
.A2(n_573),
.B(n_679),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_745),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_742),
.B(n_625),
.Y(n_826)
);

BUFx5_ASAP7_75t_L g827 ( 
.A(n_735),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_694),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_755),
.B(n_707),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_R g830 ( 
.A(n_758),
.B(n_638),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_785),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_759),
.B(n_625),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_729),
.B(n_634),
.Y(n_833)
);

INVxp33_ASAP7_75t_L g834 ( 
.A(n_693),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_704),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_690),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_703),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_R g838 ( 
.A(n_697),
.B(n_638),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_735),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_736),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_736),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_760),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_760),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_762),
.B(n_603),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_774),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_738),
.B(n_565),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_762),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_696),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_696),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_698),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_698),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_744),
.B(n_651),
.Y(n_852)
);

BUFx6f_ASAP7_75t_SL g853 ( 
.A(n_712),
.Y(n_853)
);

XOR2xp5_ASAP7_75t_L g854 ( 
.A(n_700),
.B(n_102),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_717),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_699),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_747),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_699),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_722),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_722),
.Y(n_860)
);

INVx4_ASAP7_75t_SL g861 ( 
.A(n_763),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_726),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_702),
.B(n_663),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_723),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_731),
.B(n_627),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_723),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_725),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_766),
.B(n_634),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_725),
.Y(n_869)
);

BUFx6f_ASAP7_75t_SL g870 ( 
.A(n_712),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_772),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_708),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_746),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_786),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_727),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_744),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_721),
.B(n_663),
.Y(n_877)
);

NAND2x1p5_ASAP7_75t_L g878 ( 
.A(n_764),
.B(n_651),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_788),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_716),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_705),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_713),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_761),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_711),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_701),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_734),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_805),
.B(n_810),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_805),
.B(n_743),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_840),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_790),
.B(n_659),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_810),
.B(n_750),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_880),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_839),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_841),
.Y(n_894)
);

NAND2x1p5_ASAP7_75t_L g895 ( 
.A(n_855),
.B(n_659),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_855),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_865),
.B(n_771),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_855),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_826),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_795),
.B(n_776),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_842),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_843),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_863),
.B(n_662),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_847),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_827),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_862),
.B(n_871),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_795),
.B(n_662),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_806),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_832),
.B(n_670),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_792),
.B(n_670),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_827),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_803),
.B(n_814),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_819),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_814),
.A2(n_741),
.B(n_677),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_845),
.B(n_802),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_845),
.B(n_676),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_827),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_844),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_823),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_816),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_873),
.B(n_718),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_829),
.B(n_676),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_817),
.A2(n_684),
.B(n_683),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_853),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_820),
.B(n_684),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_792),
.B(n_646),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_818),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_799),
.Y(n_928)
);

OR2x6_ASAP7_75t_L g929 ( 
.A(n_867),
.B(n_734),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_831),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_817),
.B(n_637),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_792),
.B(n_815),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_792),
.B(n_656),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_823),
.B(n_637),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_857),
.B(n_720),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_875),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_807),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_859),
.B(n_697),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_792),
.B(n_739),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_809),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_868),
.B(n_733),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_811),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_812),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_877),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_852),
.B(n_639),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_813),
.Y(n_946)
);

INVxp67_ASAP7_75t_SL g947 ( 
.A(n_822),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_825),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_852),
.B(n_640),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_796),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_879),
.B(n_833),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_836),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_SL g953 ( 
.A(n_857),
.B(n_787),
.Y(n_953)
);

OR2x2_ASAP7_75t_SL g954 ( 
.A(n_791),
.B(n_681),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_878),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_860),
.B(n_688),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_837),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_879),
.B(n_640),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_878),
.Y(n_959)
);

AND2x2_ASAP7_75t_SL g960 ( 
.A(n_883),
.B(n_768),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_884),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_835),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_868),
.B(n_815),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_793),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_833),
.B(n_695),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_874),
.B(n_682),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_848),
.B(n_682),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_849),
.B(n_600),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_850),
.B(n_600),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_864),
.B(n_574),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_797),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_798),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_882),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_824),
.B(n_661),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_801),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_804),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_851),
.B(n_604),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_856),
.B(n_604),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_858),
.B(n_614),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_866),
.B(n_614),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_887),
.B(n_876),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_919),
.B(n_906),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_896),
.B(n_882),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_912),
.B(n_834),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_973),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_893),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_919),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_896),
.B(n_869),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_893),
.Y(n_989)
);

NOR2x1_ASAP7_75t_L g990 ( 
.A(n_959),
.B(n_846),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_892),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_901),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_951),
.Y(n_993)
);

AND2x2_ASAP7_75t_SL g994 ( 
.A(n_888),
.B(n_778),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_887),
.B(n_872),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_901),
.Y(n_996)
);

OR2x6_ASAP7_75t_L g997 ( 
.A(n_929),
.B(n_886),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_915),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_901),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_951),
.Y(n_1000)
);

NOR2x1_ASAP7_75t_L g1001 ( 
.A(n_959),
.B(n_821),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_L g1002 ( 
.A(n_923),
.B(n_881),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_954),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_891),
.B(n_824),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_928),
.B(n_808),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_919),
.B(n_861),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_906),
.B(n_861),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_929),
.B(n_886),
.Y(n_1008)
);

NAND2x1p5_ASAP7_75t_L g1009 ( 
.A(n_896),
.B(n_886),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_SL g1010 ( 
.A(n_959),
.B(n_769),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_896),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_902),
.Y(n_1012)
);

OR2x6_ASAP7_75t_L g1013 ( 
.A(n_929),
.B(n_765),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_915),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_906),
.B(n_861),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_906),
.B(n_828),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_944),
.B(n_885),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_902),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_928),
.B(n_794),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_920),
.Y(n_1020)
);

INVx5_ASAP7_75t_L g1021 ( 
.A(n_973),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_920),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_938),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_938),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_944),
.B(n_775),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_890),
.B(n_706),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_SL g1027 ( 
.A(n_959),
.B(n_853),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_890),
.B(n_854),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_931),
.B(n_789),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_966),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_898),
.B(n_537),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_958),
.B(n_966),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_913),
.B(n_781),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_929),
.B(n_870),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_898),
.B(n_537),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_958),
.B(n_641),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_898),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_898),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_940),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_923),
.B(n_870),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_922),
.B(n_641),
.Y(n_1041)
);

AND2x6_ASAP7_75t_L g1042 ( 
.A(n_932),
.B(n_970),
.Y(n_1042)
);

OR2x6_ASAP7_75t_L g1043 ( 
.A(n_929),
.B(n_838),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_937),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_920),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_937),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_937),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_940),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_973),
.B(n_800),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_938),
.Y(n_1050)
);

AO21x2_ASAP7_75t_L g1051 ( 
.A1(n_932),
.A2(n_830),
.B(n_838),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_899),
.B(n_105),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_943),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_938),
.B(n_653),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_948),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_943),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_899),
.B(n_107),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_930),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_991),
.Y(n_1059)
);

INVx6_ASAP7_75t_SL g1060 ( 
.A(n_997),
.Y(n_1060)
);

INVx8_ASAP7_75t_L g1061 ( 
.A(n_1042),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_1049),
.A2(n_941),
.B1(n_921),
.B2(n_960),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_986),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_982),
.B(n_955),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_1003),
.Y(n_1065)
);

BUFx12f_ASAP7_75t_L g1066 ( 
.A(n_1034),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_982),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_985),
.A2(n_911),
.B(n_905),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_1032),
.Y(n_1069)
);

INVx3_ASAP7_75t_SL g1070 ( 
.A(n_1034),
.Y(n_1070)
);

BUFx8_ASAP7_75t_SL g1071 ( 
.A(n_997),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_986),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_1007),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_1007),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1036),
.B(n_903),
.Y(n_1075)
);

BUFx12f_ASAP7_75t_L g1076 ( 
.A(n_1008),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_1015),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_993),
.B(n_1000),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_1030),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_1039),
.Y(n_1080)
);

BUFx4_ASAP7_75t_SL g1081 ( 
.A(n_1008),
.Y(n_1081)
);

BUFx12f_ASAP7_75t_L g1082 ( 
.A(n_1013),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_1005),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_989),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_992),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_1017),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_1015),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_1006),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_1038),
.B(n_955),
.Y(n_1089)
);

CKINVDCx8_ASAP7_75t_R g1090 ( 
.A(n_1016),
.Y(n_1090)
);

CKINVDCx16_ASAP7_75t_R g1091 ( 
.A(n_1010),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_1039),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_1038),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_1006),
.Y(n_1094)
);

BUFx2_ASAP7_75t_SL g1095 ( 
.A(n_1016),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_985),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_985),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_1011),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_996),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_1017),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_1023),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_1025),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_1039),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_1024),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_984),
.B(n_903),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1011),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_996),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1019),
.B(n_935),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1029),
.B(n_909),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1028),
.B(n_998),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_987),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_1050),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_999),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_1009),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1014),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1012),
.Y(n_1116)
);

AO21x1_ASAP7_75t_L g1117 ( 
.A1(n_1002),
.A2(n_963),
.B(n_965),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_1021),
.Y(n_1118)
);

INVxp67_ASAP7_75t_SL g1119 ( 
.A(n_1055),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1021),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_987),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1021),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1012),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_987),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_1037),
.B(n_955),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1111),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_1111),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1112),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1063),
.Y(n_1129)
);

INVx6_ASAP7_75t_L g1130 ( 
.A(n_1059),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1062),
.A2(n_981),
.B1(n_995),
.B2(n_1033),
.Y(n_1131)
);

INVx6_ASAP7_75t_L g1132 ( 
.A(n_1059),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1110),
.A2(n_960),
.B1(n_1040),
.B2(n_994),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1078),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_1083),
.Y(n_1135)
);

BUFx2_ASAP7_75t_SL g1136 ( 
.A(n_1112),
.Y(n_1136)
);

INVx5_ASAP7_75t_L g1137 ( 
.A(n_1120),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1072),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_1081),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1084),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1111),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1108),
.A2(n_960),
.B1(n_1040),
.B2(n_914),
.Y(n_1142)
);

INVx6_ASAP7_75t_L g1143 ( 
.A(n_1066),
.Y(n_1143)
);

OAI22xp33_ASAP7_75t_SL g1144 ( 
.A1(n_1091),
.A2(n_953),
.B1(n_1010),
.B2(n_914),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1085),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1083),
.A2(n_1025),
.B1(n_990),
.B2(n_1026),
.Y(n_1146)
);

NAND2x1p5_ASAP7_75t_L g1147 ( 
.A(n_1096),
.B(n_1037),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1071),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1115),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1095),
.A2(n_1027),
.B1(n_1043),
.B2(n_973),
.Y(n_1150)
);

AOI22x1_ASAP7_75t_SL g1151 ( 
.A1(n_1065),
.A2(n_924),
.B1(n_927),
.B2(n_894),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1109),
.A2(n_1004),
.B(n_897),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_SL g1153 ( 
.A1(n_1102),
.A2(n_1043),
.B1(n_1051),
.B2(n_939),
.Y(n_1153)
);

CKINVDCx11_ASAP7_75t_R g1154 ( 
.A(n_1070),
.Y(n_1154)
);

CKINVDCx11_ASAP7_75t_R g1155 ( 
.A(n_1066),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_SL g1156 ( 
.A(n_1060),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_SL g1157 ( 
.A1(n_1065),
.A2(n_954),
.B1(n_936),
.B2(n_1054),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_SL g1158 ( 
.A1(n_1102),
.A2(n_1057),
.B1(n_1052),
.B2(n_922),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1109),
.A2(n_1105),
.B1(n_1069),
.B2(n_1075),
.Y(n_1159)
);

BUFx10_ASAP7_75t_L g1160 ( 
.A(n_1079),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1105),
.A2(n_956),
.B1(n_945),
.B2(n_949),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1069),
.A2(n_907),
.B1(n_1107),
.B2(n_1099),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1111),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1086),
.B(n_1052),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_1120),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1075),
.A2(n_956),
.B1(n_945),
.B2(n_949),
.Y(n_1166)
);

OAI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_1090),
.A2(n_990),
.B1(n_900),
.B2(n_907),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1100),
.A2(n_1041),
.B1(n_1042),
.B2(n_1057),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1101),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1103),
.Y(n_1170)
);

INVx6_ASAP7_75t_L g1171 ( 
.A(n_1076),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1116),
.Y(n_1172)
);

CKINVDCx11_ASAP7_75t_R g1173 ( 
.A(n_1082),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1123),
.A2(n_918),
.B1(n_900),
.B2(n_983),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1104),
.B(n_934),
.Y(n_1175)
);

NAND2x1p5_ASAP7_75t_L g1176 ( 
.A(n_1096),
.B(n_1048),
.Y(n_1176)
);

OAI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1090),
.A2(n_1054),
.B1(n_927),
.B2(n_894),
.Y(n_1177)
);

CKINVDCx11_ASAP7_75t_R g1178 ( 
.A(n_1082),
.Y(n_1178)
);

CKINVDCx8_ASAP7_75t_R g1179 ( 
.A(n_1064),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1113),
.B(n_918),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1133),
.A2(n_1079),
.B1(n_988),
.B2(n_1089),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1144),
.A2(n_1117),
.B1(n_930),
.B2(n_1067),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1144),
.A2(n_1117),
.B1(n_930),
.B2(n_1067),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1157),
.A2(n_1061),
.B1(n_647),
.B2(n_916),
.Y(n_1184)
);

OAI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1146),
.A2(n_904),
.B1(n_1074),
.B2(n_1073),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1175),
.B(n_1073),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1140),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1142),
.A2(n_904),
.B1(n_957),
.B2(n_962),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1151),
.A2(n_1061),
.B1(n_647),
.B2(n_925),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_SL g1190 ( 
.A1(n_1167),
.A2(n_1061),
.B1(n_1077),
.B2(n_1074),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1145),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1167),
.A2(n_1136),
.B1(n_1131),
.B2(n_1135),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1158),
.A2(n_1001),
.B(n_910),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_1149),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1177),
.A2(n_910),
.B(n_967),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1153),
.A2(n_952),
.B1(n_942),
.B2(n_940),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1150),
.A2(n_1001),
.B(n_961),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1130),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1159),
.A2(n_952),
.B1(n_942),
.B2(n_940),
.Y(n_1199)
);

OAI21xp33_ASAP7_75t_L g1200 ( 
.A1(n_1161),
.A2(n_1166),
.B(n_1152),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1164),
.A2(n_940),
.B1(n_895),
.B2(n_943),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1172),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1168),
.A2(n_969),
.B(n_968),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1128),
.A2(n_1061),
.B1(n_1087),
.B2(n_1088),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1129),
.Y(n_1205)
);

CKINVDCx14_ASAP7_75t_R g1206 ( 
.A(n_1155),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1152),
.A2(n_946),
.B1(n_972),
.B2(n_971),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1143),
.A2(n_1094),
.B1(n_1114),
.B2(n_1125),
.Y(n_1208)
);

INVx5_ASAP7_75t_L g1209 ( 
.A(n_1137),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1134),
.B(n_968),
.Y(n_1210)
);

BUFx12f_ASAP7_75t_L g1211 ( 
.A(n_1173),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1162),
.A2(n_975),
.B1(n_976),
.B2(n_964),
.Y(n_1212)
);

INVx5_ASAP7_75t_SL g1213 ( 
.A(n_1141),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1138),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1169),
.B(n_969),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1179),
.A2(n_1089),
.B1(n_1125),
.B2(n_1060),
.Y(n_1216)
);

BUFx4f_ASAP7_75t_SL g1217 ( 
.A(n_1139),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1162),
.B(n_977),
.Y(n_1218)
);

INVx8_ASAP7_75t_L g1219 ( 
.A(n_1137),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1174),
.A2(n_979),
.B(n_978),
.Y(n_1220)
);

BUFx5_ASAP7_75t_L g1221 ( 
.A(n_1160),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1180),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1171),
.A2(n_1122),
.B1(n_1120),
.B2(n_1097),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1141),
.B(n_1121),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1154),
.A2(n_976),
.B1(n_889),
.B2(n_1020),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1132),
.B(n_980),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1192),
.A2(n_1178),
.B1(n_1132),
.B2(n_889),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1195),
.A2(n_1022),
.B1(n_1058),
.B2(n_1045),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1222),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1200),
.A2(n_889),
.B1(n_606),
.B2(n_574),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1181),
.A2(n_1156),
.B1(n_1137),
.B2(n_1148),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1185),
.A2(n_606),
.B1(n_574),
.B2(n_1060),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1182),
.B(n_1141),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1184),
.A2(n_606),
.B1(n_574),
.B2(n_908),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1190),
.A2(n_606),
.B1(n_908),
.B2(n_1124),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1189),
.A2(n_908),
.B1(n_1018),
.B2(n_1160),
.Y(n_1236)
);

AOI211xp5_ASAP7_75t_L g1237 ( 
.A1(n_1203),
.A2(n_980),
.B(n_655),
.C(n_657),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1187),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1225),
.A2(n_1147),
.B1(n_1176),
.B2(n_1165),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1210),
.B(n_1163),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1183),
.B(n_1163),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1196),
.A2(n_1093),
.B1(n_1119),
.B2(n_1118),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1191),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1188),
.A2(n_950),
.B1(n_1046),
.B2(n_1044),
.Y(n_1244)
);

OAI222xp33_ASAP7_75t_L g1245 ( 
.A1(n_1204),
.A2(n_1056),
.B1(n_1053),
.B2(n_1047),
.C1(n_1046),
.C2(n_1127),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1218),
.A2(n_1047),
.B1(n_1056),
.B2(n_1053),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1194),
.B(n_1205),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1216),
.A2(n_1122),
.B1(n_1098),
.B2(n_1106),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1209),
.A2(n_1122),
.B1(n_1098),
.B2(n_1106),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1214),
.B(n_1126),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1208),
.A2(n_1106),
.B1(n_1098),
.B2(n_1055),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1186),
.A2(n_970),
.B1(n_933),
.B2(n_926),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1197),
.A2(n_1048),
.B1(n_1080),
.B2(n_1092),
.Y(n_1253)
);

OAI222xp33_ASAP7_75t_L g1254 ( 
.A1(n_1223),
.A2(n_1092),
.B1(n_1080),
.B2(n_947),
.C1(n_1068),
.C2(n_974),
.Y(n_1254)
);

AOI222xp33_ASAP7_75t_L g1255 ( 
.A1(n_1220),
.A2(n_653),
.B1(n_655),
.B2(n_657),
.C1(n_674),
.C2(n_685),
.Y(n_1255)
);

OAI221xp5_ASAP7_75t_L g1256 ( 
.A1(n_1193),
.A2(n_974),
.B1(n_1035),
.B2(n_1031),
.C(n_685),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1226),
.A2(n_1170),
.B1(n_1103),
.B2(n_917),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1199),
.A2(n_1170),
.B1(n_1103),
.B2(n_917),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1207),
.A2(n_1211),
.B1(n_1201),
.B2(n_1215),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1202),
.A2(n_905),
.B1(n_560),
.B2(n_626),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1206),
.A2(n_579),
.B1(n_630),
.B2(n_571),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1221),
.A2(n_577),
.B1(n_571),
.B2(n_587),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1224),
.B(n_71),
.Y(n_1263)
);

NOR3xp33_ASAP7_75t_L g1264 ( 
.A(n_1198),
.B(n_72),
.C(n_73),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1221),
.Y(n_1265)
);

AOI221xp5_ASAP7_75t_L g1266 ( 
.A1(n_1212),
.A2(n_575),
.B1(n_577),
.B2(n_584),
.C(n_585),
.Y(n_1266)
);

OAI221xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1264),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.C(n_76),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1231),
.A2(n_1227),
.B(n_1255),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1255),
.A2(n_1217),
.B1(n_1219),
.B2(n_1209),
.Y(n_1269)
);

OAI21xp33_ASAP7_75t_L g1270 ( 
.A1(n_1259),
.A2(n_1263),
.B(n_1237),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1229),
.B(n_1213),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1237),
.B(n_1209),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1243),
.B(n_76),
.Y(n_1273)
);

AND2x2_ASAP7_75t_SL g1274 ( 
.A(n_1228),
.B(n_1219),
.Y(n_1274)
);

OAI221xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1236),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.C(n_80),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1228),
.A2(n_1256),
.B(n_1254),
.Y(n_1276)
);

OAI221xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1261),
.A2(n_78),
.B1(n_81),
.B2(n_83),
.C(n_85),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1247),
.B(n_1238),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1240),
.B(n_81),
.Y(n_1279)
);

AND2x2_ASAP7_75t_SL g1280 ( 
.A(n_1233),
.B(n_88),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_L g1281 ( 
.A(n_1248),
.B(n_633),
.C(n_591),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1241),
.B(n_108),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1250),
.B(n_110),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1265),
.B(n_113),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1234),
.A2(n_114),
.B(n_118),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1239),
.A2(n_633),
.B(n_591),
.Y(n_1286)
);

NAND3xp33_ASAP7_75t_L g1287 ( 
.A(n_1257),
.B(n_1232),
.C(n_1235),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1246),
.B(n_121),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1252),
.B(n_125),
.Y(n_1289)
);

OAI221xp5_ASAP7_75t_L g1290 ( 
.A1(n_1249),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.C(n_130),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1260),
.B(n_131),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1260),
.A2(n_1245),
.B(n_1230),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1251),
.B(n_552),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1244),
.A2(n_570),
.B1(n_558),
.B2(n_141),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1253),
.B(n_138),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1258),
.B(n_142),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1242),
.B(n_145),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1262),
.A2(n_570),
.B1(n_558),
.B2(n_147),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1278),
.B(n_1266),
.Y(n_1299)
);

OA211x2_ASAP7_75t_L g1300 ( 
.A1(n_1270),
.A2(n_1272),
.B(n_1286),
.C(n_1269),
.Y(n_1300)
);

NAND4xp75_ASAP7_75t_L g1301 ( 
.A(n_1280),
.B(n_146),
.C(n_148),
.D(n_149),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1273),
.B(n_156),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1268),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_1303)
);

OA211x2_ASAP7_75t_L g1304 ( 
.A1(n_1269),
.A2(n_1293),
.B(n_1281),
.C(n_1295),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1267),
.B(n_173),
.C(n_174),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1274),
.B(n_175),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1274),
.B(n_179),
.Y(n_1307)
);

NOR2x1_ASAP7_75t_L g1308 ( 
.A(n_1271),
.B(n_186),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1279),
.B(n_196),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1282),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1276),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1282),
.B(n_1276),
.Y(n_1312)
);

NAND3xp33_ASAP7_75t_L g1313 ( 
.A(n_1277),
.B(n_202),
.C(n_212),
.Y(n_1313)
);

AOI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1275),
.A2(n_307),
.B1(n_213),
.B2(n_214),
.C(n_220),
.Y(n_1314)
);

OAI211xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1283),
.A2(n_222),
.B(n_223),
.C(n_225),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1312),
.B(n_1276),
.Y(n_1316)
);

NAND4xp75_ASAP7_75t_L g1317 ( 
.A(n_1300),
.B(n_1291),
.C(n_1289),
.D(n_1292),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1305),
.B(n_1294),
.C(n_1297),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1310),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1306),
.B(n_1284),
.Y(n_1320)
);

XNOR2xp5_ASAP7_75t_L g1321 ( 
.A(n_1303),
.B(n_1287),
.Y(n_1321)
);

XOR2xp5_ASAP7_75t_L g1322 ( 
.A(n_1301),
.B(n_1298),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1299),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1313),
.A2(n_1289),
.B1(n_1285),
.B2(n_1290),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1302),
.Y(n_1325)
);

INVxp67_ASAP7_75t_SL g1326 ( 
.A(n_1308),
.Y(n_1326)
);

XOR2x2_ASAP7_75t_L g1327 ( 
.A(n_1321),
.B(n_1314),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1324),
.A2(n_1304),
.B1(n_1311),
.B2(n_1315),
.Y(n_1328)
);

XOR2x2_ASAP7_75t_L g1329 ( 
.A(n_1322),
.B(n_1307),
.Y(n_1329)
);

AOI22x1_ASAP7_75t_SL g1330 ( 
.A1(n_1327),
.A2(n_1326),
.B1(n_1323),
.B2(n_1325),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1328),
.A2(n_1317),
.B1(n_1324),
.B2(n_1318),
.Y(n_1331)
);

XOR2x2_ASAP7_75t_L g1332 ( 
.A(n_1329),
.B(n_1318),
.Y(n_1332)
);

OA22x2_ASAP7_75t_L g1333 ( 
.A1(n_1331),
.A2(n_1316),
.B1(n_1319),
.B2(n_1320),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1333),
.A2(n_1331),
.B1(n_1330),
.B2(n_1332),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_SL g1335 ( 
.A1(n_1334),
.A2(n_1309),
.B(n_1288),
.C(n_1296),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1335),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1336),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1337),
.Y(n_1338)
);

INVxp33_ASAP7_75t_SL g1339 ( 
.A(n_1338),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1339),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1340),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1341),
.A2(n_260),
.B1(n_264),
.B2(n_267),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1342),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1342),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1343),
.A2(n_268),
.B1(n_269),
.B2(n_272),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1344),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1346),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1345),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_L g1349 ( 
.A1(n_1348),
.A2(n_276),
.B1(n_280),
.B2(n_281),
.C(n_284),
.Y(n_1349)
);

AOI211xp5_ASAP7_75t_L g1350 ( 
.A1(n_1349),
.A2(n_1347),
.B(n_295),
.C(n_297),
.Y(n_1350)
);


endmodule