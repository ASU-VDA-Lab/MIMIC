module fake_jpeg_5696_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_32),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_21),
.B1(n_17),
.B2(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_0),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_17),
.B1(n_26),
.B2(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_58),
.Y(n_87)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_61),
.Y(n_94)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_30),
.B1(n_26),
.B2(n_21),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_47),
.B1(n_24),
.B2(n_39),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_70),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_16),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_47),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_19),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_40),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_45),
.B1(n_22),
.B2(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_88),
.B1(n_91),
.B2(n_99),
.Y(n_112)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_82),
.Y(n_117)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_29),
.B1(n_59),
.B2(n_73),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_36),
.B1(n_48),
.B2(n_24),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_90),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_39),
.B1(n_36),
.B2(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_66),
.Y(n_101)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g130 ( 
.A(n_98),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_47),
.B1(n_35),
.B2(n_34),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_101),
.B(n_126),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_44),
.C(n_41),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_68),
.B1(n_48),
.B2(n_54),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_109),
.B1(n_116),
.B2(n_82),
.Y(n_131)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_107),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_108),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_97),
.B1(n_52),
.B2(n_49),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_40),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_127),
.Y(n_138)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_118),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_119),
.B1(n_120),
.B2(n_125),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_59),
.B1(n_71),
.B2(n_53),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_92),
.B1(n_93),
.B2(n_80),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_80),
.B1(n_93),
.B2(n_78),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_65),
.B1(n_53),
.B2(n_67),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_65),
.B1(n_67),
.B2(n_73),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_124),
.Y(n_147)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_76),
.A2(n_65),
.B1(n_67),
.B2(n_63),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_33),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_65),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_44),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_33),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_35),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_115),
.B1(n_107),
.B2(n_124),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_137),
.B1(n_139),
.B2(n_157),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_92),
.B1(n_86),
.B2(n_41),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_98),
.B1(n_86),
.B2(n_34),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_98),
.B1(n_41),
.B2(n_46),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_111),
.B1(n_130),
.B2(n_118),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_141),
.A2(n_144),
.B1(n_150),
.B2(n_151),
.Y(n_185)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_117),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_46),
.A3(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_155),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_46),
.C(n_29),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_113),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_121),
.B(n_102),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_105),
.A2(n_32),
.B1(n_28),
.B2(n_27),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_29),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_128),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_163),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_165),
.A2(n_167),
.B1(n_180),
.B2(n_0),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_101),
.B(n_138),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_169),
.B(n_179),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_101),
.B1(n_129),
.B2(n_126),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_101),
.B1(n_129),
.B2(n_126),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_127),
.B(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_129),
.B1(n_126),
.B2(n_102),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_181),
.B1(n_184),
.B2(n_142),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_136),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_176),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_130),
.B(n_106),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_139),
.B1(n_157),
.B2(n_140),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_186),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_134),
.A2(n_32),
.B(n_28),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_0),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_150),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_145),
.C(n_149),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_189),
.C(n_199),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_133),
.C(n_152),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_194),
.B1(n_210),
.B2(n_213),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_147),
.B1(n_137),
.B2(n_151),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_183),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_200),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_147),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_205),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_166),
.C(n_169),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_207),
.C(n_215),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_182),
.B(n_177),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_146),
.C(n_28),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_173),
.Y(n_232)
);

AOI22x1_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_146),
.B1(n_27),
.B2(n_20),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_179),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_211),
.Y(n_235)
);

AO22x2_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_27),
.B1(n_20),
.B2(n_146),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_167),
.B(n_15),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_220),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_197),
.A2(n_210),
.B1(n_211),
.B2(n_209),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_231),
.B1(n_222),
.B2(n_242),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_159),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_226),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_168),
.B(n_163),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_165),
.C(n_178),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_SL g261 ( 
.A(n_227),
.B(n_236),
.C(n_241),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_181),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_230),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_164),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_170),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_189),
.B(n_170),
.C(n_164),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_239),
.C(n_206),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_207),
.C(n_215),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_186),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_179),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_201),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_197),
.A2(n_214),
.B1(n_193),
.B2(n_204),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_242),
.A2(n_213),
.B1(n_160),
.B2(n_190),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_249),
.B1(n_253),
.B2(n_265),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_251),
.C(n_263),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_213),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_259),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_160),
.B1(n_208),
.B2(n_213),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_206),
.C(n_190),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_205),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_226),
.C(n_219),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_176),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_260),
.B(n_232),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_162),
.B1(n_179),
.B2(n_184),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_257),
.A2(n_227),
.B1(n_5),
.B2(n_6),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_2),
.C(n_3),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_15),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_237),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_259),
.CI(n_261),
.CON(n_287),
.SN(n_287)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_218),
.B1(n_233),
.B2(n_236),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_280),
.B1(n_260),
.B2(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_271),
.A2(n_272),
.B(n_279),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_274),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_238),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_283),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_237),
.C(n_240),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_278),
.C(n_282),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_223),
.Y(n_277)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_217),
.C(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_252),
.B(n_15),
.Y(n_281)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_4),
.C(n_5),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_14),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_14),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_296),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_254),
.C(n_243),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_293),
.C(n_12),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_262),
.B1(n_255),
.B2(n_246),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_291),
.A2(n_298),
.B1(n_13),
.B2(n_12),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_275),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_5),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_267),
.C(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_273),
.A2(n_278),
.B1(n_267),
.B2(n_282),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_266),
.A2(n_270),
.B1(n_280),
.B2(n_283),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_270),
.B(n_264),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_12),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_14),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_302),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_294),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_314),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_313),
.C(n_289),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_307),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_11),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_4),
.Y(n_308)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_4),
.Y(n_309)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_311),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_6),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_6),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_298),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_285),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_321),
.B(n_322),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_307),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_305),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_329),
.C(n_318),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_311),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_327),
.B(n_330),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_306),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_331),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_291),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_287),
.B(n_286),
.C(n_313),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_286),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_299),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_7),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_336),
.B(n_337),
.Y(n_339)
);

OAI321xp33_ASAP7_75t_L g336 ( 
.A1(n_326),
.A2(n_318),
.A3(n_327),
.B1(n_324),
.B2(n_10),
.C(n_7),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_335),
.A2(n_7),
.B(n_8),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_338),
.A2(n_333),
.B(n_9),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_339),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_8),
.C(n_9),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_9),
.B(n_10),
.Y(n_344)
);


endmodule