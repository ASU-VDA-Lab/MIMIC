module fake_jpeg_4966_n_315 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_44),
.B(n_47),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_1),
.C(n_2),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_46),
.B(n_60),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_52),
.Y(n_93)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_26),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_2),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_54),
.B(n_59),
.Y(n_107)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_61),
.B1(n_66),
.B2(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_64),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_58),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_36),
.B(n_3),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_68),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_3),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_27),
.B(n_3),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_27),
.B(n_43),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_19),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_32),
.B1(n_42),
.B2(n_38),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_72),
.A2(n_82),
.B1(n_102),
.B2(n_111),
.Y(n_134)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_75),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_74),
.B(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_79),
.Y(n_130)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_87),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_33),
.B1(n_25),
.B2(n_40),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_32),
.Y(n_83)
);

OR2x2_ASAP7_75t_SL g136 ( 
.A(n_83),
.B(n_100),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_22),
.B(n_20),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_86),
.A2(n_110),
.B(n_34),
.C(n_55),
.Y(n_141)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

CKINVDCx9p33_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_31),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_61),
.B1(n_53),
.B2(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_56),
.A2(n_42),
.B1(n_20),
.B2(n_41),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_28),
.B1(n_39),
.B2(n_35),
.Y(n_124)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_49),
.B(n_59),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_43),
.B1(n_41),
.B2(n_28),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_39),
.C(n_35),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_54),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_131),
.Y(n_154)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_122),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_83),
.B(n_20),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_121),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_85),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_134),
.B1(n_100),
.B2(n_143),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_60),
.B1(n_40),
.B2(n_33),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_144),
.B1(n_102),
.B2(n_70),
.Y(n_169)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_128),
.Y(n_168)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_133),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_4),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_141),
.B(n_8),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_83),
.B(n_55),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_113),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_82),
.A2(n_34),
.B1(n_40),
.B2(n_33),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_86),
.A2(n_34),
.B1(n_25),
.B2(n_7),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_95),
.B1(n_77),
.B2(n_70),
.Y(n_151)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_5),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_6),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_155),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_111),
.A3(n_81),
.B1(n_72),
.B2(n_110),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_181),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_157),
.B1(n_178),
.B2(n_125),
.Y(n_185)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_95),
.B1(n_77),
.B2(n_74),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_166),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_105),
.B(n_90),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_165),
.B(n_171),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_164),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_93),
.B(n_84),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_184),
.B1(n_171),
.B2(n_181),
.Y(n_190)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_170),
.B(n_172),
.Y(n_187)
);

AO22x1_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_78),
.B1(n_89),
.B2(n_92),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_101),
.C(n_106),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_133),
.C(n_143),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_175),
.B(n_176),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_116),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_117),
.A2(n_25),
.B1(n_101),
.B2(n_16),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_8),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_117),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_184),
.B(n_10),
.C(n_11),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_192),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_212),
.B1(n_146),
.B2(n_115),
.Y(n_238)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_153),
.A2(n_157),
.B1(n_152),
.B2(n_162),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_194),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_121),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_132),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_202),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_126),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_201),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_175),
.A2(n_136),
.B1(n_149),
.B2(n_138),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_131),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_136),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_209),
.Y(n_233)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_170),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_211),
.B(n_146),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_128),
.B1(n_149),
.B2(n_138),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_156),
.B(n_183),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_226),
.B(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_220),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_178),
.B1(n_166),
.B2(n_160),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_198),
.B(n_188),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_221),
.B(n_196),
.Y(n_246)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_227),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_166),
.B(n_180),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_161),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_231),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_230),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_129),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_190),
.B(n_127),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_207),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_208),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_237),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_200),
.A2(n_114),
.B1(n_155),
.B2(n_179),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_191),
.B(n_199),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_187),
.Y(n_237)
);

AOI221xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_239),
.B1(n_210),
.B2(n_199),
.C(n_14),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_186),
.B(n_12),
.C(n_13),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_243),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_194),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_257),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_197),
.C(n_213),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_251),
.C(n_258),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_254),
.B1(n_232),
.B2(n_224),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_185),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_189),
.B(n_214),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_217),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_240),
.B1(n_224),
.B2(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_265),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_252),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_226),
.C(n_228),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_269),
.C(n_270),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_254),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_268),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_241),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_225),
.C(n_236),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_258),
.C(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_247),
.B1(n_255),
.B2(n_236),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_263),
.B1(n_283),
.B2(n_277),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_244),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_284),
.C(n_220),
.Y(n_296)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_280),
.A2(n_282),
.B(n_285),
.Y(n_290)
);

XOR2x2_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_240),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_229),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_269),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_216),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_222),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_291),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_281),
.B(n_275),
.Y(n_289)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_264),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_241),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_264),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_295),
.A3(n_250),
.B1(n_262),
.B2(n_227),
.C1(n_242),
.C2(n_234),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_273),
.B1(n_223),
.B2(n_248),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_245),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_300),
.C(n_287),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_237),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_292),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_289),
.B1(n_293),
.B2(n_296),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_305),
.B(n_303),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_308),
.B(n_297),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_207),
.Y(n_308)
);

A2O1A1O1Ixp25_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_310),
.B(n_308),
.C(n_205),
.D(n_204),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_SL g311 ( 
.A(n_307),
.B(n_291),
.C(n_298),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_204),
.A3(n_215),
.B1(n_164),
.B2(n_205),
.C1(n_12),
.C2(n_13),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_312),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_313),
.Y(n_315)
);


endmodule