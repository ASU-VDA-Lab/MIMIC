module real_jpeg_7758_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_17;
wire n_57;
wire n_43;
wire n_37;
wire n_21;
wire n_54;
wire n_65;
wire n_35;
wire n_33;
wire n_50;
wire n_38;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_10;
wire n_31;
wire n_52;
wire n_67;
wire n_58;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_14;
wire n_71;
wire n_51;
wire n_45;
wire n_25;
wire n_47;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_70;
wire n_41;
wire n_26;
wire n_56;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_32;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_0),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_1),
.A2(n_17),
.B1(n_19),
.B2(n_24),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_6),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

HAxp5_ASAP7_75t_SL g55 ( 
.A(n_4),
.B(n_56),
.CON(n_55),
.SN(n_55)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_49),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_8),
.A2(n_14),
.B1(n_15),
.B2(n_22),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_29),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_27),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_23),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_19),
.B(n_21),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_19),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_21),
.B(n_24),
.C(n_25),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_26),
.C(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_25),
.A2(n_26),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_67),
.B(n_72),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_51),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_42),
.B(n_50),
.Y(n_31)
);

NOR3xp33_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_52),
.C(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_38),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.C(n_37),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_47),
.C(n_49),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_62),
.B(n_66),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_55),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_60),
.B(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_56),
.B(n_60),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_70),
.Y(n_71)
);


endmodule