module fake_jpeg_30957_n_361 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_361);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_361;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_23),
.B(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_43),
.B(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_47),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_8),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_62),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_7),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_102),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_26),
.B1(n_30),
.B2(n_22),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_81),
.A2(n_85),
.B1(n_87),
.B2(n_105),
.Y(n_141)
);

HAxp5_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_39),
.CON(n_83),
.SN(n_83)
);

OR2x2_ASAP7_75t_SL g148 ( 
.A(n_83),
.B(n_118),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_36),
.B1(n_26),
.B2(n_24),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_30),
.B1(n_36),
.B2(n_19),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_36),
.C(n_24),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_94),
.B(n_106),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_36),
.B1(n_24),
.B2(n_20),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_97),
.B1(n_103),
.B2(n_104),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_13),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_38),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_49),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_57),
.A2(n_32),
.B1(n_37),
.B2(n_35),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_30),
.B1(n_28),
.B2(n_35),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_37),
.C(n_34),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_64),
.A2(n_19),
.B1(n_33),
.B2(n_38),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_107),
.A2(n_111),
.B1(n_114),
.B2(n_0),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_63),
.A2(n_33),
.B1(n_38),
.B2(n_3),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_10),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_116),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_65),
.A2(n_38),
.B1(n_10),
.B2(n_3),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_72),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_31),
.Y(n_118)
);

NAND2x1_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_31),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_124),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_12),
.B(n_15),
.C(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_123),
.B(n_150),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_79),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_125),
.B(n_133),
.Y(n_196)
);

OR2x4_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_13),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

AO22x1_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_58),
.B1(n_45),
.B2(n_31),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_132),
.A2(n_95),
.B1(n_108),
.B2(n_93),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_31),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_119),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_139),
.B(n_142),
.Y(n_197)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_75),
.B(n_31),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g144 ( 
.A(n_119),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_6),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_149),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_98),
.B(n_4),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_98),
.A2(n_15),
.B(n_4),
.C(n_5),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_153),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_90),
.B(n_84),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_155),
.Y(n_175)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_102),
.A2(n_9),
.B1(n_14),
.B2(n_1),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_160),
.B1(n_84),
.B2(n_88),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_94),
.B(n_1),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_117),
.Y(n_177)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_155),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_113),
.A2(n_1),
.B1(n_9),
.B2(n_117),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_118),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_126),
.B(n_9),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_168),
.B(n_182),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_174),
.Y(n_220)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_86),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_77),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_180),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_77),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_117),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_183),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_93),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_146),
.C(n_120),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_90),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_186),
.B(n_195),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_131),
.B1(n_147),
.B2(n_153),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_128),
.B(n_78),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_132),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_78),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_129),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_143),
.Y(n_201)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_88),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_180),
.A2(n_141),
.B1(n_143),
.B2(n_132),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_198),
.A2(n_200),
.B1(n_203),
.B2(n_206),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_SL g200 ( 
.A1(n_187),
.A2(n_150),
.B(n_136),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_201),
.B(n_222),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_202),
.A2(n_225),
.B(n_230),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_136),
.B(n_123),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_205),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_161),
.A2(n_188),
.B1(n_182),
.B2(n_177),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_161),
.A2(n_140),
.B1(n_89),
.B2(n_95),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_215),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_137),
.Y(n_212)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_154),
.B(n_121),
.C(n_159),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_213),
.Y(n_259)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_130),
.A3(n_89),
.B1(n_135),
.B2(n_138),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_130),
.C(n_197),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_218),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_130),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_224),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_162),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_223),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_184),
.B1(n_170),
.B2(n_167),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_169),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_170),
.B1(n_167),
.B2(n_196),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_165),
.A2(n_185),
.B1(n_178),
.B2(n_166),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_192),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_228),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_174),
.A2(n_192),
.B1(n_171),
.B2(n_196),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_227),
.A2(n_165),
.B1(n_166),
.B2(n_190),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_189),
.A2(n_171),
.B(n_178),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_185),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_250),
.C(n_231),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_260),
.B1(n_204),
.B2(n_218),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_229),
.Y(n_236)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_237),
.B(n_242),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_207),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_248),
.Y(n_269)
);

AOI22x1_ASAP7_75t_L g247 ( 
.A1(n_198),
.A2(n_165),
.B1(n_191),
.B2(n_176),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_208),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_191),
.C(n_190),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_173),
.B(n_176),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_211),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_259),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_220),
.A2(n_173),
.B(n_202),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_226),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_210),
.A2(n_173),
.B1(n_199),
.B2(n_212),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_249),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_275),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_220),
.B1(n_206),
.B2(n_199),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_278),
.B1(n_283),
.B2(n_232),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_271),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_267),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_274),
.B1(n_280),
.B2(n_253),
.Y(n_286)
);

NOR4xp25_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_221),
.C(n_217),
.D(n_204),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_227),
.C(n_233),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_243),
.C(n_266),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_256),
.B1(n_254),
.B2(n_246),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_241),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_238),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_251),
.A2(n_242),
.B1(n_245),
.B2(n_240),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_234),
.B(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_269),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_256),
.A2(n_239),
.B1(n_260),
.B2(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_251),
.A2(n_245),
.B1(n_240),
.B2(n_247),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_256),
.B1(n_247),
.B2(n_257),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_287),
.Y(n_303)
);

AOI221xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_267),
.B1(n_270),
.B2(n_271),
.C(n_261),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_298),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_258),
.B1(n_250),
.B2(n_243),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_300),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_294),
.Y(n_308)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_262),
.A2(n_272),
.B(n_281),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_287),
.B(n_285),
.Y(n_304)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_281),
.B1(n_278),
.B2(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_277),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_306),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_294),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_305),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_280),
.B(n_274),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_316),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_302),
.C(n_284),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_277),
.Y(n_310)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_284),
.A2(n_277),
.B(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_288),
.B(n_295),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_308),
.B(n_291),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_322),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_308),
.B(n_302),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_327),
.C(n_320),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_301),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_329),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_293),
.B1(n_296),
.B2(n_290),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_328),
.B(n_330),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_290),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_300),
.C(n_312),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_325),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_313),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_332),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_333),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_303),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_323),
.B(n_318),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_337),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_310),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_311),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_312),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_320),
.B1(n_304),
.B2(n_313),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_346),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_342),
.B(n_344),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_315),
.C(n_303),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g352 ( 
.A(n_347),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_343),
.A2(n_331),
.B(n_340),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_353),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_334),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g354 ( 
.A(n_350),
.B(n_345),
.C(n_348),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_355),
.Y(n_358)
);

OAI21x1_ASAP7_75t_L g355 ( 
.A1(n_351),
.A2(n_342),
.B(n_346),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_356),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_357),
.B(n_314),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_359),
.A2(n_314),
.B1(n_358),
.B2(n_352),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_360),
.Y(n_361)
);


endmodule