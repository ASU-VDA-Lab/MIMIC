module real_jpeg_12170_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_139;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_4),
.A2(n_38),
.B1(n_43),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_4),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_4),
.A2(n_24),
.B1(n_28),
.B2(n_65),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_38),
.B1(n_43),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_6),
.A2(n_40),
.B1(n_48),
.B2(n_56),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_6),
.A2(n_24),
.B1(n_28),
.B2(n_56),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_7),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_7),
.A2(n_27),
.B1(n_38),
.B2(n_43),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_9),
.B(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_9),
.B(n_24),
.C(n_62),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_9),
.A2(n_31),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_9),
.B(n_50),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_10),
.A2(n_40),
.B1(n_48),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_10),
.A2(n_38),
.B1(n_43),
.B2(n_52),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_10),
.A2(n_24),
.B1(n_28),
.B2(n_52),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_11),
.A2(n_24),
.B1(n_28),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_13),
.A2(n_24),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_95),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_94),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_66),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_66),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_45),
.C(n_53),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_19),
.A2(n_20),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_35),
.B2(n_36),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_21),
.B(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_32),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_30),
.Y(n_134)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_24),
.A2(n_28),
.B1(n_60),
.B2(n_62),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_28),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_29),
.B(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_29),
.A2(n_30),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_31),
.A2(n_77),
.B(n_79),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_31),
.B(n_41),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_31),
.A2(n_110),
.B1(n_118),
.B2(n_119),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B(n_39),
.C(n_42),
.Y(n_36)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_40),
.B1(n_44),
.B2(n_48),
.Y(n_47)
);

OA22x2_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_49)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_43),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_38),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_45)
);

HAxp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_41),
.CON(n_39),
.SN(n_39)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_43),
.C(n_44),
.Y(n_42)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_48),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_41),
.B(n_107),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_45),
.B(n_53),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_46),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_55),
.A2(n_58),
.B1(n_106),
.B2(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_SL g62 ( 
.A(n_60),
.Y(n_62)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_85),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_81),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_136),
.B(n_141),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_125),
.B(n_135),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_113),
.B(n_124),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_108),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_108),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_119),
.B(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_120),
.B(n_123),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_122),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_127),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_140),
.Y(n_141)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);


endmodule