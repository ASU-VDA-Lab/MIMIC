module fake_jpeg_14019_n_401 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_401);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_401;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_44),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_45),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_47),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_59),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_52),
.Y(n_139)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g105 ( 
.A(n_53),
.Y(n_105)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_55),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_17),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_74),
.Y(n_110)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g116 ( 
.A(n_65),
.Y(n_116)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_14),
.B(n_0),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_17),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_80),
.B(n_93),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_21),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_82),
.Y(n_112)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_90),
.Y(n_130)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_94),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_16),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_35),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_42),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_99),
.B(n_84),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_74),
.B1(n_48),
.B2(n_88),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_115),
.B1(n_30),
.B2(n_28),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_60),
.A2(n_23),
.B1(n_40),
.B2(n_32),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_44),
.B(n_23),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_119),
.B(n_93),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_59),
.A2(n_30),
.B1(n_40),
.B2(n_27),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_134),
.B1(n_28),
.B2(n_27),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_133),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_49),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_57),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_102),
.A2(n_55),
.B1(n_65),
.B2(n_33),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_147),
.A2(n_29),
.B1(n_26),
.B2(n_25),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_150),
.A2(n_47),
.B1(n_81),
.B2(n_92),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_153),
.A2(n_157),
.B1(n_169),
.B2(n_190),
.Y(n_213)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_95),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_185),
.C(n_191),
.Y(n_206)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_25),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_173),
.Y(n_198)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_168),
.Y(n_195)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_167),
.B(n_174),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_105),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_73),
.B1(n_77),
.B2(n_86),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_110),
.B(n_33),
.Y(n_173)
);

AOI32xp33_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_35),
.A3(n_19),
.B1(n_32),
.B2(n_29),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_26),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_178),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_105),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_19),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_136),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_183),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_99),
.B(n_87),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_98),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

OAI32xp33_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_133),
.A3(n_127),
.B1(n_145),
.B2(n_52),
.Y(n_194)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_140),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_185),
.Y(n_227)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_137),
.A3(n_103),
.B1(n_116),
.B2(n_146),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_158),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_173),
.B(n_103),
.CI(n_116),
.CON(n_199),
.SN(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_199),
.A2(n_130),
.B(n_105),
.C(n_112),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_135),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_130),
.C(n_154),
.Y(n_244)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_153),
.B1(n_213),
.B2(n_205),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_224),
.A2(n_225),
.B1(n_243),
.B2(n_116),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_185),
.B1(n_169),
.B2(n_156),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_234),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_227),
.A2(n_245),
.B(n_246),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_201),
.B(n_185),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_228),
.A2(n_237),
.B(n_241),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_206),
.A2(n_193),
.B1(n_157),
.B2(n_194),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_232),
.B1(n_242),
.B2(n_97),
.Y(n_263)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_156),
.B1(n_170),
.B2(n_141),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_198),
.B(n_199),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_209),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_166),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_239),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_166),
.B(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_178),
.B(n_155),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_212),
.A2(n_172),
.B1(n_164),
.B2(n_171),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_196),
.A2(n_158),
.B1(n_184),
.B2(n_182),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_219),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_192),
.A2(n_181),
.B1(n_136),
.B2(n_165),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_244),
.C(n_225),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_253),
.A2(n_246),
.B(n_224),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_256),
.B1(n_242),
.B2(n_262),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_227),
.A2(n_212),
.B1(n_203),
.B2(n_101),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_228),
.A2(n_230),
.B(n_233),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_261),
.B(n_246),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_203),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_260),
.B(n_268),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_222),
.A2(n_204),
.B(n_208),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_129),
.B1(n_101),
.B2(n_139),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_234),
.B1(n_192),
.B2(n_129),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_208),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_267),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_207),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_237),
.B(n_207),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_232),
.C(n_231),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_277),
.C(n_281),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_264),
.B(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_261),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_273),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_274),
.A2(n_253),
.B(n_257),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_250),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_275),
.Y(n_299)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_240),
.C(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_284),
.B1(n_272),
.B2(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_243),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_287),
.B1(n_261),
.B2(n_254),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_234),
.B1(n_204),
.B2(n_217),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_162),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_139),
.B1(n_218),
.B2(n_200),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_218),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_288),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_294),
.B(n_297),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_253),
.B1(n_256),
.B2(n_264),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_253),
.B(n_257),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_298),
.A2(n_308),
.B1(n_217),
.B2(n_210),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_305),
.B1(n_307),
.B2(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_249),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_266),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_262),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_279),
.A2(n_263),
.B1(n_265),
.B2(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_280),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_323),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_306),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_295),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_270),
.C(n_286),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_315),
.C(n_319),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_281),
.C(n_277),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_287),
.B1(n_285),
.B2(n_258),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_316),
.A2(n_326),
.B1(n_327),
.B2(n_292),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_275),
.B1(n_284),
.B2(n_265),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_318),
.A2(n_322),
.B1(n_304),
.B2(n_292),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_309),
.B(n_247),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_325),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_273),
.C(n_289),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_200),
.C(n_159),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_303),
.B1(n_300),
.B2(n_294),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_289),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_291),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_247),
.Y(n_324)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_324),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_297),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_308),
.A2(n_282),
.B1(n_258),
.B2(n_131),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_301),
.Y(n_328)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_328),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_329),
.B(n_337),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_330),
.A2(n_333),
.B1(n_191),
.B2(n_186),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_336),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_301),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_332),
.B(n_120),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_335),
.A2(n_311),
.B1(n_180),
.B2(n_189),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_210),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_112),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_339),
.Y(n_346)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_340),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_310),
.A2(n_321),
.B1(n_317),
.B2(n_314),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_343),
.A2(n_326),
.B1(n_327),
.B2(n_311),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_344),
.B(n_336),
.C(n_342),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_347),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_223),
.Y(n_348)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_350),
.A2(n_344),
.B1(n_329),
.B2(n_331),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_352),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_354),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_117),
.C(n_109),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_56),
.C(n_51),
.Y(n_369)
);

FAx1_ASAP7_75t_SL g357 ( 
.A(n_330),
.B(n_1),
.CI(n_2),
.CON(n_357),
.SN(n_357)
);

A2O1A1Ixp33_ASAP7_75t_L g364 ( 
.A1(n_357),
.A2(n_349),
.B(n_356),
.C(n_351),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_106),
.Y(n_358)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_358),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_346),
.B(n_343),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_6),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_363),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_364),
.A2(n_357),
.B1(n_353),
.B2(n_6),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_347),
.A2(n_121),
.B(n_137),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_367),
.A2(n_5),
.B(n_6),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_3),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_46),
.C(n_4),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_3),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_372),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_366),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_357),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_373),
.A2(n_376),
.B(n_365),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_355),
.C(n_350),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_375),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_353),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_378),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_373),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_382),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_372),
.A2(n_359),
.B1(n_368),
.B2(n_364),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_386),
.B(n_387),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_376),
.A2(n_370),
.B(n_369),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_384),
.B(n_380),
.C(n_363),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_392),
.C(n_7),
.Y(n_393)
);

NAND2x1_ASAP7_75t_SL g391 ( 
.A(n_383),
.B(n_371),
.Y(n_391)
);

OAI21x1_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_7),
.B(n_9),
.Y(n_395)
);

XOR2x2_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_381),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_393),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_390),
.B(n_7),
.C(n_8),
.Y(n_394)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_394),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_397),
.A2(n_389),
.B1(n_395),
.B2(n_10),
.Y(n_398)
);

OAI321xp33_ASAP7_75t_L g399 ( 
.A1(n_398),
.A2(n_396),
.A3(n_389),
.B1(n_10),
.B2(n_12),
.C(n_13),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_399),
.A2(n_7),
.B(n_9),
.Y(n_400)
);

NOR3xp33_ASAP7_75t_SL g401 ( 
.A(n_400),
.B(n_12),
.C(n_13),
.Y(n_401)
);


endmodule