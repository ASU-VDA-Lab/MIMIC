module real_aes_353_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_618;
wire n_778;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_555;
wire n_421;
wire n_852;
wire n_766;
wire n_1113;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_884;
wire n_666;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_816;
wire n_400;
wire n_539;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_1108;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_1078;
wire n_744;
wire n_938;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_1031;
wire n_432;
wire n_1103;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_1041;
wire n_501;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_957;
wire n_995;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_898;
wire n_734;
wire n_604;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1083;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_787;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1045;
wire n_465;
wire n_473;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_652;
wire n_1097;
wire n_703;
wire n_500;
wire n_601;
wire n_1101;
wire n_1076;
wire n_463;
wire n_661;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_1104;
wire n_842;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_0), .A2(n_349), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_1), .A2(n_232), .B1(n_522), .B2(n_523), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g915 ( .A1(n_2), .A2(n_176), .B1(n_456), .B2(n_721), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_3), .A2(n_128), .B1(n_445), .B2(n_565), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_4), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_5), .A2(n_94), .B1(n_482), .B2(n_584), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_6), .B(n_601), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_7), .A2(n_55), .B1(n_445), .B2(n_565), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_8), .A2(n_268), .B1(n_612), .B2(n_613), .Y(n_827) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_9), .A2(n_345), .B1(n_485), .B2(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_10), .A2(n_295), .B1(n_594), .B2(n_672), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_11), .A2(n_384), .B1(n_434), .B2(n_902), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_12), .A2(n_215), .B1(n_619), .B2(n_620), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_13), .A2(n_91), .B1(n_491), .B2(n_757), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g988 ( .A1(n_14), .A2(n_93), .B1(n_607), .B2(n_608), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_15), .A2(n_112), .B1(n_675), .B2(n_731), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_16), .A2(n_343), .B1(n_546), .B2(n_793), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_17), .A2(n_257), .B1(n_439), .B2(n_444), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_18), .A2(n_95), .B1(n_631), .B2(n_951), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_19), .A2(n_233), .B1(n_605), .B2(n_822), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_20), .A2(n_194), .B1(n_583), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_SL g831 ( .A1(n_21), .A2(n_192), .B1(n_523), .B2(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_22), .A2(n_368), .B1(n_674), .B2(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_23), .A2(n_157), .B1(n_510), .B2(n_700), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_24), .A2(n_68), .B1(n_506), .B2(n_507), .Y(n_788) );
AO222x2_ASAP7_75t_L g967 ( .A1(n_25), .A2(n_152), .B1(n_254), .B2(n_532), .C1(n_537), .C2(n_800), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_26), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_27), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_28), .A2(n_356), .B1(n_822), .B2(n_971), .Y(n_970) );
INVx1_ASAP7_75t_SL g417 ( .A(n_29), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g1047 ( .A(n_29), .B(n_45), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_30), .A2(n_364), .B1(n_476), .B2(n_546), .Y(n_1069) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_31), .Y(n_984) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_32), .A2(n_186), .B1(n_595), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_33), .A2(n_395), .B1(n_589), .B2(n_591), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_34), .A2(n_141), .B1(n_451), .B2(n_456), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g1087 ( .A(n_35), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_36), .B(n_410), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_37), .A2(n_304), .B1(n_619), .B2(n_620), .Y(n_618) );
AOI22x1_ASAP7_75t_L g995 ( .A1(n_38), .A2(n_208), .B1(n_484), .B2(n_619), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_39), .A2(n_308), .B1(n_570), .B2(n_654), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_40), .A2(n_228), .B1(n_434), .B2(n_510), .Y(n_1072) );
OA22x2_ASAP7_75t_L g850 ( .A1(n_41), .A2(n_851), .B1(n_852), .B2(n_880), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_41), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_42), .A2(n_292), .B1(n_683), .B2(n_686), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_43), .A2(n_202), .B1(n_607), .B2(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_44), .A2(n_347), .B1(n_467), .B2(n_731), .Y(n_894) );
AO22x2_ASAP7_75t_L g419 ( .A1(n_45), .A2(n_376), .B1(n_416), .B2(n_420), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_46), .A2(n_184), .B1(n_553), .B2(n_554), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_47), .A2(n_224), .B1(n_671), .B2(n_672), .Y(n_1002) );
CKINVDCx20_ASAP7_75t_R g1097 ( .A(n_48), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_49), .A2(n_378), .B1(n_674), .B2(n_675), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_50), .A2(n_58), .B1(n_506), .B2(n_574), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g926 ( .A1(n_51), .A2(n_346), .B1(n_671), .B2(n_672), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_52), .A2(n_159), .B1(n_462), .B2(n_467), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_53), .A2(n_197), .B1(n_445), .B2(n_500), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_54), .A2(n_296), .B1(n_551), .B2(n_731), .Y(n_1003) );
INVx1_ASAP7_75t_L g418 ( .A(n_56), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_57), .A2(n_327), .B1(n_617), .B2(n_620), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_59), .A2(n_250), .B1(n_471), .B2(n_474), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_60), .A2(n_312), .B1(n_510), .B2(n_679), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_61), .A2(n_310), .B1(n_474), .B2(n_546), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_62), .A2(n_324), .B1(n_619), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_63), .A2(n_150), .B1(n_515), .B2(n_519), .Y(n_629) );
AOI22xp33_ASAP7_75t_SL g922 ( .A1(n_64), .A2(n_332), .B1(n_731), .B2(n_923), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_65), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_66), .A2(n_372), .B1(n_479), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_67), .A2(n_319), .B1(n_519), .B2(n_520), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_69), .A2(n_262), .B1(n_565), .B2(n_718), .Y(n_717) );
AO21x1_ASAP7_75t_SL g1051 ( .A1(n_70), .A2(n_1052), .B(n_1060), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_71), .A2(n_367), .B1(n_734), .B2(n_898), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_72), .A2(n_227), .B1(n_675), .B2(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_73), .A2(n_363), .B1(n_476), .B2(n_546), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_74), .B(n_410), .Y(n_749) );
AO22x2_ASAP7_75t_L g426 ( .A1(n_75), .A2(n_203), .B1(n_416), .B2(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_76), .A2(n_210), .B1(n_583), .B2(n_585), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_77), .A2(n_328), .B1(n_583), .B2(n_672), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_78), .A2(n_149), .B1(n_620), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_79), .A2(n_253), .B1(n_474), .B2(n_546), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_80), .A2(n_154), .B1(n_780), .B2(n_923), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_81), .A2(n_120), .B1(n_535), .B2(n_538), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_82), .A2(n_369), .B1(n_451), .B2(n_574), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_83), .A2(n_172), .B1(n_607), .B2(n_608), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_84), .A2(n_302), .B1(n_487), .B2(n_707), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_85), .A2(n_339), .B1(n_484), .B2(n_487), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_86), .A2(n_177), .B1(n_620), .B2(n_829), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_87), .A2(n_213), .B1(n_467), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_88), .A2(n_350), .B1(n_631), .B2(n_634), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_89), .A2(n_167), .B1(n_484), .B2(n_553), .Y(n_614) );
AOI22xp33_ASAP7_75t_SL g974 ( .A1(n_90), .A2(n_126), .B1(n_612), .B2(n_613), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_92), .A2(n_211), .B1(n_510), .B2(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_96), .A2(n_265), .B1(n_537), .B2(n_538), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_97), .A2(n_377), .B1(n_585), .B2(n_874), .C(n_876), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_98), .A2(n_116), .B1(n_479), .B2(n_482), .Y(n_478) );
AOI222xp33_ASAP7_75t_L g687 ( .A1(n_99), .A2(n_158), .B1(n_248), .B2(n_444), .C1(n_503), .C2(n_688), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_100), .A2(n_204), .B1(n_507), .B2(n_653), .Y(n_945) );
OAI22x1_ASAP7_75t_L g624 ( .A1(n_101), .A2(n_625), .B1(n_626), .B2(n_659), .Y(n_624) );
INVx1_ASAP7_75t_L g659 ( .A(n_101), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_102), .A2(n_252), .B1(n_520), .B2(n_671), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_103), .A2(n_390), .B1(n_445), .B2(n_565), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_104), .A2(n_246), .B1(n_476), .B2(n_631), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g1009 ( .A1(n_105), .A2(n_321), .B1(n_658), .B2(n_902), .Y(n_1009) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_106), .A2(n_293), .B1(n_686), .B2(n_777), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_107), .A2(n_142), .B1(n_736), .B2(n_737), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_108), .A2(n_342), .B1(n_578), .B2(n_700), .Y(n_946) );
AO222x2_ASAP7_75t_L g819 ( .A1(n_109), .A2(n_223), .B1(n_381), .B2(n_532), .C1(n_605), .C2(n_608), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_110), .A2(n_249), .B1(n_570), .B2(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g856 ( .A(n_111), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_113), .A2(n_267), .B1(n_520), .B2(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_114), .A2(n_269), .B1(n_537), .B2(n_538), .Y(n_824) );
AOI222xp33_ASAP7_75t_L g1010 ( .A1(n_115), .A2(n_189), .B1(n_361), .B2(n_445), .C1(n_688), .C2(n_768), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_117), .A2(n_140), .B1(n_639), .B2(n_640), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g1019 ( .A1(n_118), .A2(n_205), .B1(n_874), .B2(n_1020), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_119), .A2(n_226), .B1(n_653), .B2(n_654), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_121), .A2(n_353), .B1(n_479), .B2(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_122), .B(n_409), .Y(n_408) );
AO22x2_ASAP7_75t_L g423 ( .A1(n_123), .A2(n_298), .B1(n_416), .B2(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_124), .A2(n_318), .B1(n_699), .B2(n_700), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_125), .Y(n_865) );
OAI22x1_ASAP7_75t_L g785 ( .A1(n_127), .A2(n_786), .B1(n_801), .B2(n_802), .Y(n_785) );
CKINVDCx16_ASAP7_75t_R g802 ( .A(n_127), .Y(n_802) );
AO21x2_ASAP7_75t_L g1013 ( .A1(n_129), .A2(n_1014), .B(n_1033), .Y(n_1013) );
NOR2xp33_ASAP7_75t_L g1033 ( .A(n_129), .B(n_1016), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_130), .A2(n_134), .B1(n_644), .B2(n_1027), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_131), .A2(n_283), .B1(n_589), .B2(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_132), .A2(n_240), .B1(n_463), .B2(n_551), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_133), .A2(n_151), .B1(n_594), .B2(n_595), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_135), .A2(n_259), .B1(n_456), .B2(n_721), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_136), .A2(n_281), .B1(n_450), .B2(n_455), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_137), .A2(n_261), .B1(n_467), .B2(n_875), .Y(n_949) );
INVx1_ASAP7_75t_L g1011 ( .A(n_138), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_139), .B(n_410), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_143), .A2(n_251), .B1(n_491), .B2(n_674), .Y(n_955) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_144), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_145), .A2(n_287), .B1(n_445), .B2(n_565), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_146), .A2(n_245), .B1(n_489), .B2(n_589), .Y(n_1068) );
OA22x2_ASAP7_75t_L g404 ( .A1(n_147), .A2(n_405), .B1(n_406), .B2(n_492), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_147), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_148), .Y(n_1100) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_153), .A2(n_181), .B1(n_510), .B2(n_726), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_155), .A2(n_165), .B1(n_829), .B2(n_832), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_156), .A2(n_351), .B1(n_456), .B2(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_160), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_161), .A2(n_190), .B1(n_657), .B2(n_658), .Y(n_1025) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_162), .A2(n_239), .B1(n_551), .B2(n_671), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_163), .A2(n_258), .B1(n_565), .B2(n_904), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_164), .B(n_859), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_166), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_168), .A2(n_234), .B1(n_551), .B2(n_637), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_169), .B(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_170), .A2(n_300), .B1(n_472), .B2(n_476), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_171), .A2(n_386), .B1(n_429), .B2(n_658), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_173), .B(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_174), .A2(n_200), .B1(n_487), .B2(n_489), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_175), .A2(n_338), .B1(n_546), .B2(n_547), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_178), .A2(n_303), .B1(n_671), .B2(n_672), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g924 ( .A1(n_179), .A2(n_320), .B1(n_474), .B2(n_546), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_180), .A2(n_217), .B1(n_657), .B2(n_658), .Y(n_1112) );
INVx1_ASAP7_75t_L g909 ( .A(n_182), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_183), .A2(n_371), .B1(n_553), .B2(n_954), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_185), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_187), .A2(n_284), .B1(n_578), .B2(n_679), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g1104 ( .A(n_188), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_191), .B(n_1089), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_193), .A2(n_362), .B1(n_484), .B2(n_519), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_195), .B(n_768), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_196), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_198), .A2(n_220), .B1(n_456), .B2(n_506), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_199), .A2(n_272), .B1(n_506), .B2(n_574), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_201), .A2(n_278), .B1(n_506), .B2(n_574), .Y(n_1074) );
INVx1_ASAP7_75t_L g1046 ( .A(n_203), .Y(n_1046) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_206), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_207), .A2(n_274), .B1(n_612), .B2(n_613), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_209), .A2(n_1062), .B1(n_1075), .B2(n_1076), .Y(n_1061) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_209), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_212), .A2(n_329), .B1(n_657), .B2(n_658), .Y(n_656) );
XNOR2xp5_ASAP7_75t_L g979 ( .A(n_214), .B(n_980), .Y(n_979) );
XNOR2xp5_ASAP7_75t_L g998 ( .A(n_214), .B(n_980), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_216), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_218), .A2(n_379), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g821 ( .A1(n_219), .A2(n_337), .B1(n_822), .B2(n_823), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_221), .A2(n_746), .B1(n_747), .B2(n_759), .Y(n_745) );
INVxp67_ASAP7_75t_L g759 ( .A(n_221), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_222), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g1107 ( .A(n_225), .Y(n_1107) );
CKINVDCx20_ASAP7_75t_R g1092 ( .A(n_229), .Y(n_1092) );
OA22x2_ASAP7_75t_L g889 ( .A1(n_230), .A2(n_890), .B1(n_891), .B2(n_906), .Y(n_889) );
INVxp67_ASAP7_75t_L g906 ( .A(n_230), .Y(n_906) );
OA22x2_ASAP7_75t_L g958 ( .A1(n_230), .A2(n_890), .B1(n_891), .B2(n_906), .Y(n_958) );
XNOR2x1_ASAP7_75t_L g560 ( .A(n_231), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g1057 ( .A(n_235), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g1085 ( .A(n_236), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_237), .A2(n_391), .B1(n_523), .B2(n_617), .Y(n_977) );
OA22x2_ASAP7_75t_L g713 ( .A1(n_238), .A2(n_714), .B1(n_739), .B2(n_740), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_238), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_241), .A2(n_288), .B1(n_585), .B2(n_589), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g1103 ( .A(n_242), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_243), .A2(n_260), .B1(n_554), .B2(n_734), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_244), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_247), .A2(n_266), .B1(n_451), .B2(n_456), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_255), .A2(n_294), .B1(n_472), .B2(n_686), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_256), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_263), .A2(n_816), .B1(n_817), .B2(n_834), .Y(n_815) );
INVx1_ASAP7_75t_L g834 ( .A(n_263), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_264), .A2(n_360), .B1(n_429), .B2(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g983 ( .A(n_270), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_271), .A2(n_317), .B1(n_506), .B2(n_507), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_273), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_275), .A2(n_285), .B1(n_445), .B2(n_565), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_276), .A2(n_335), .B1(n_429), .B2(n_434), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g969 ( .A1(n_277), .A2(n_297), .B1(n_608), .B2(n_823), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_279), .A2(n_397), .B1(n_522), .B2(n_523), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_280), .B(n_503), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_282), .A2(n_315), .B1(n_445), .B2(n_500), .Y(n_499) );
AOI22x1_ASAP7_75t_L g762 ( .A1(n_286), .A2(n_763), .B1(n_764), .B2(n_784), .Y(n_762) );
INVx1_ASAP7_75t_L g784 ( .A(n_286), .Y(n_784) );
XNOR2x1_ASAP7_75t_L g805 ( .A(n_286), .B(n_764), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_289), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_290), .A2(n_375), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_291), .A2(n_370), .B1(n_472), .B2(n_547), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g1044 ( .A(n_298), .B(n_1045), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_299), .A2(n_374), .B1(n_565), .B2(n_904), .Y(n_1073) );
AOI222xp33_ASAP7_75t_L g798 ( .A1(n_301), .A2(n_316), .B1(n_357), .B2(n_532), .C1(n_799), .C2(n_800), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_305), .A2(n_359), .B1(n_523), .B2(n_617), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_306), .B(n_410), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_307), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_309), .A2(n_396), .B1(n_546), .B2(n_547), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_311), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_313), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_314), .A2(n_352), .B1(n_1029), .B2(n_1031), .Y(n_1028) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_322), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g895 ( .A1(n_323), .A2(n_340), .B1(n_547), .B2(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g956 ( .A(n_325), .Y(n_956) );
INVx3_ASAP7_75t_L g416 ( .A(n_326), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_330), .A2(n_341), .B1(n_523), .B2(n_617), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g1109 ( .A(n_331), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_333), .A2(n_385), .B1(n_434), .B2(n_578), .Y(n_916) );
OAI22x1_ASAP7_75t_L g692 ( .A1(n_334), .A2(n_693), .B1(n_710), .B2(n_711), .Y(n_692) );
INVx1_ASAP7_75t_L g711 ( .A(n_334), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_336), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_344), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g1113 ( .A(n_348), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_354), .A2(n_387), .B1(n_672), .B2(n_731), .Y(n_1066) );
XNOR2x1_ASAP7_75t_L g836 ( .A(n_355), .B(n_837), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_358), .Y(n_533) );
INVx1_ASAP7_75t_L g527 ( .A(n_365), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_366), .A2(n_394), .B1(n_510), .B2(n_511), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_373), .A2(n_383), .B1(n_456), .B2(n_506), .Y(n_677) );
INVx1_ASAP7_75t_L g1041 ( .A(n_380), .Y(n_1041) );
NAND2xp5_ASAP7_75t_SL g1058 ( .A(n_380), .B(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1042 ( .A(n_382), .Y(n_1042) );
AND2x2_ASAP7_75t_R g1078 ( .A(n_382), .B(n_1041), .Y(n_1078) );
OA22x2_ASAP7_75t_L g666 ( .A1(n_388), .A2(n_667), .B1(n_668), .B2(n_689), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_388), .Y(n_667) );
INVxp67_ASAP7_75t_L g1059 ( .A(n_389), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_392), .B(n_503), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_393), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_1048), .B(n_1051), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_884), .B(n_1038), .Y(n_399) );
INVx1_ASAP7_75t_L g1050 ( .A(n_400), .Y(n_1050) );
XOR2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_661), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_556), .B1(n_557), .B2(n_660), .Y(n_401) );
INVx2_ASAP7_75t_L g660 ( .A(n_402), .Y(n_660) );
AOI22x1_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_404), .B1(n_493), .B2(n_555), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g492 ( .A(n_406), .Y(n_492) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_460), .Y(n_406) );
NAND4xp25_ASAP7_75t_SL g407 ( .A(n_408), .B(n_428), .C(n_438), .D(n_449), .Y(n_407) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g503 ( .A(n_411), .Y(n_503) );
INVx4_ASAP7_75t_SL g601 ( .A(n_411), .Y(n_601) );
BUFx2_ASAP7_75t_L g647 ( .A(n_411), .Y(n_647) );
INVx3_ASAP7_75t_SL g697 ( .A(n_411), .Y(n_697) );
INVx4_ASAP7_75t_SL g768 ( .A(n_411), .Y(n_768) );
INVx6_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_421), .Y(n_412) );
AND2x4_ASAP7_75t_L g436 ( .A(n_413), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g457 ( .A(n_413), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g532 ( .A(n_413), .B(n_421), .Y(n_532) );
AND2x2_ASAP7_75t_L g605 ( .A(n_413), .B(n_458), .Y(n_605) );
AND2x2_ASAP7_75t_L g608 ( .A(n_413), .B(n_437), .Y(n_608) );
AND2x2_ASAP7_75t_L g790 ( .A(n_413), .B(n_437), .Y(n_790) );
AND2x2_ASAP7_75t_L g971 ( .A(n_413), .B(n_458), .Y(n_971) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_419), .Y(n_413) );
INVx2_ASAP7_75t_L g433 ( .A(n_414), .Y(n_433) );
AND2x2_ASAP7_75t_L g442 ( .A(n_414), .B(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_414), .Y(n_448) );
OAI22x1_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_416), .Y(n_420) );
INVx2_ASAP7_75t_L g424 ( .A(n_416), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_416), .Y(n_427) );
AND2x2_ASAP7_75t_L g432 ( .A(n_419), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g443 ( .A(n_419), .Y(n_443) );
BUFx2_ASAP7_75t_L g477 ( .A(n_419), .Y(n_477) );
AND2x4_ASAP7_75t_L g465 ( .A(n_421), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g481 ( .A(n_421), .B(n_432), .Y(n_481) );
AND2x4_ASAP7_75t_L g488 ( .A(n_421), .B(n_442), .Y(n_488) );
AND2x2_ASAP7_75t_L g522 ( .A(n_421), .B(n_442), .Y(n_522) );
AND2x2_ASAP7_75t_L g617 ( .A(n_421), .B(n_442), .Y(n_617) );
AND2x6_ASAP7_75t_L g619 ( .A(n_421), .B(n_432), .Y(n_619) );
AND2x2_ASAP7_75t_L g829 ( .A(n_421), .B(n_466), .Y(n_829) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g431 ( .A(n_423), .B(n_425), .Y(n_431) );
AND2x2_ASAP7_75t_L g447 ( .A(n_423), .B(n_426), .Y(n_447) );
INVx1_ASAP7_75t_L g454 ( .A(n_423), .Y(n_454) );
INVxp67_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g453 ( .A(n_426), .B(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g510 ( .A(n_430), .Y(n_510) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_430), .Y(n_578) );
BUFx2_ASAP7_75t_L g902 ( .A(n_430), .Y(n_902) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AND2x2_ASAP7_75t_L g441 ( .A(n_431), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g485 ( .A(n_431), .B(n_466), .Y(n_485) );
AND2x4_ASAP7_75t_L g537 ( .A(n_431), .B(n_442), .Y(n_537) );
AND2x2_ASAP7_75t_L g607 ( .A(n_431), .B(n_432), .Y(n_607) );
AND2x2_ASAP7_75t_L g823 ( .A(n_431), .B(n_432), .Y(n_823) );
AND2x2_ASAP7_75t_L g832 ( .A(n_431), .B(n_466), .Y(n_832) );
AND2x2_ASAP7_75t_L g473 ( .A(n_432), .B(n_453), .Y(n_473) );
AND2x2_ASAP7_75t_SL g612 ( .A(n_432), .B(n_453), .Y(n_612) );
AND2x4_ASAP7_75t_L g466 ( .A(n_433), .B(n_443), .Y(n_466) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g511 ( .A(n_435), .Y(n_511) );
INVx2_ASAP7_75t_L g542 ( .A(n_435), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_435), .A2(n_576), .B1(n_577), .B2(n_579), .Y(n_575) );
INVx2_ASAP7_75t_L g658 ( .A(n_435), .Y(n_658) );
INVx2_ASAP7_75t_L g679 ( .A(n_435), .Y(n_679) );
INVx2_ASAP7_75t_SL g700 ( .A(n_435), .Y(n_700) );
INVx2_ASAP7_75t_SL g726 ( .A(n_435), .Y(n_726) );
INVx6_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g1086 ( .A(n_439), .Y(n_1086) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g501 ( .A(n_441), .Y(n_501) );
BUFx5_ASAP7_75t_L g565 ( .A(n_441), .Y(n_565) );
BUFx3_ASAP7_75t_L g645 ( .A(n_441), .Y(n_645) );
AND2x2_ASAP7_75t_L g452 ( .A(n_442), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g822 ( .A(n_442), .B(n_453), .Y(n_822) );
INVx1_ASAP7_75t_L g942 ( .A(n_444), .Y(n_942) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g650 ( .A(n_445), .Y(n_650) );
BUFx12f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx3_ASAP7_75t_L g719 ( .A(n_446), .Y(n_719) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
AND2x4_ASAP7_75t_L g476 ( .A(n_447), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g491 ( .A(n_447), .B(n_466), .Y(n_491) );
AND2x4_ASAP7_75t_L g523 ( .A(n_447), .B(n_466), .Y(n_523) );
AND2x2_ASAP7_75t_SL g538 ( .A(n_447), .B(n_448), .Y(n_538) );
AND2x4_ASAP7_75t_L g613 ( .A(n_447), .B(n_477), .Y(n_613) );
AND2x2_ASAP7_75t_SL g800 ( .A(n_447), .B(n_448), .Y(n_800) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_452), .Y(n_506) );
INVx3_ASAP7_75t_L g571 ( .A(n_452), .Y(n_571) );
AND2x4_ASAP7_75t_L g469 ( .A(n_453), .B(n_466), .Y(n_469) );
AND2x6_ASAP7_75t_L g620 ( .A(n_453), .B(n_466), .Y(n_620) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_454), .Y(n_459) );
BUFx2_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g508 ( .A(n_457), .Y(n_508) );
BUFx4f_ASAP7_75t_L g574 ( .A(n_457), .Y(n_574) );
INVx1_ASAP7_75t_L g655 ( .A(n_457), .Y(n_655) );
BUFx3_ASAP7_75t_L g1032 ( .A(n_457), .Y(n_1032) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND4xp25_ASAP7_75t_L g460 ( .A(n_461), .B(n_470), .C(n_478), .D(n_486), .Y(n_460) );
INVx1_ASAP7_75t_L g1108 ( .A(n_462), .Y(n_1108) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g519 ( .A(n_464), .Y(n_519) );
INVx3_ASAP7_75t_SL g553 ( .A(n_464), .Y(n_553) );
INVx4_ASAP7_75t_L g584 ( .A(n_464), .Y(n_584) );
INVx2_ASAP7_75t_SL g731 ( .A(n_464), .Y(n_731) );
INVx8_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g515 ( .A(n_468), .Y(n_515) );
INVx2_ASAP7_75t_L g551 ( .A(n_468), .Y(n_551) );
INVx2_ASAP7_75t_SL g595 ( .A(n_468), .Y(n_595) );
INVx2_ASAP7_75t_L g709 ( .A(n_468), .Y(n_709) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_468), .Y(n_879) );
INVx1_ASAP7_75t_SL g923 ( .A(n_468), .Y(n_923) );
INVx2_ASAP7_75t_L g1020 ( .A(n_468), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_468), .A2(n_1097), .B1(n_1098), .B2(n_1100), .Y(n_1096) );
INVx8_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_473), .Y(n_546) );
INVx2_ASAP7_75t_L g633 ( .A(n_473), .Y(n_633) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g634 ( .A(n_475), .Y(n_634) );
INVx3_ASAP7_75t_L g686 ( .A(n_475), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_475), .A2(n_865), .B1(n_866), .B2(n_868), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_475), .A2(n_1092), .B1(n_1093), .B2(n_1095), .Y(n_1091) );
INVx5_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g547 ( .A(n_476), .Y(n_547) );
BUFx2_ASAP7_75t_L g793 ( .A(n_476), .Y(n_793) );
BUFx3_ASAP7_75t_L g951 ( .A(n_476), .Y(n_951) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_SL g594 ( .A(n_480), .Y(n_594) );
INVx2_ASAP7_75t_L g671 ( .A(n_480), .Y(n_671) );
INVx2_ASAP7_75t_L g736 ( .A(n_480), .Y(n_736) );
INVx2_ASAP7_75t_SL g780 ( .A(n_480), .Y(n_780) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g637 ( .A(n_481), .Y(n_637) );
BUFx2_ASAP7_75t_L g875 ( .A(n_481), .Y(n_875) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g869 ( .A1(n_483), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g1106 ( .A1(n_483), .A2(n_1107), .B1(n_1108), .B2(n_1109), .Y(n_1106) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
BUFx3_ASAP7_75t_L g672 ( .A(n_485), .Y(n_672) );
INVx2_ASAP7_75t_L g738 ( .A(n_485), .Y(n_738) );
BUFx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx6_ASAP7_75t_L g590 ( .A(n_488), .Y(n_590) );
BUFx3_ASAP7_75t_L g757 ( .A(n_488), .Y(n_757) );
INVx2_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g898 ( .A(n_490), .Y(n_898) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g554 ( .A(n_491), .Y(n_554) );
BUFx2_ASAP7_75t_SL g585 ( .A(n_491), .Y(n_585) );
BUFx3_ASAP7_75t_L g675 ( .A(n_491), .Y(n_675) );
BUFx2_ASAP7_75t_SL g707 ( .A(n_491), .Y(n_707) );
INVx2_ASAP7_75t_L g555 ( .A(n_493), .Y(n_555) );
OA22x2_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_525), .B2(n_526), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
XOR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_524), .Y(n_495) );
NAND2x1p5_ASAP7_75t_L g496 ( .A(n_497), .B(n_512), .Y(n_496) );
NOR2x1_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_502), .Y(n_498) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_500), .Y(n_938) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g688 ( .A(n_501), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
BUFx6f_ASAP7_75t_SL g653 ( .A(n_506), .Y(n_653) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NOR2x1_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_521), .Y(n_517) );
INVx1_ASAP7_75t_L g592 ( .A(n_520), .Y(n_592) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_520), .Y(n_954) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
XNOR2x1_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
NAND2x1_ASAP7_75t_L g528 ( .A(n_529), .B(n_543), .Y(n_528) );
NOR2xp67_ASAP7_75t_L g529 ( .A(n_530), .B(n_539), .Y(n_529) );
OAI21xp5_ASAP7_75t_SL g530 ( .A1(n_531), .A2(n_533), .B(n_534), .Y(n_530) );
OAI222xp33_ASAP7_75t_L g982 ( .A1(n_531), .A2(n_536), .B1(n_983), .B2(n_984), .C1(n_985), .C2(n_986), .Y(n_982) );
INVx2_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_537), .Y(n_799) );
INVxp67_ASAP7_75t_L g986 ( .A(n_538), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_549), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_548), .Y(n_544) );
HB1xp67_ASAP7_75t_L g1094 ( .A(n_546), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_554), .Y(n_640) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI22xp5_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_559), .B1(n_622), .B2(n_623), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
XOR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_596), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_580), .Y(n_561) );
NOR3xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .C(n_575), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_564), .B(n_566), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_572), .B2(n_573), .Y(n_567) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
INVx4_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g721 ( .A(n_571), .Y(n_721) );
INVx1_ASAP7_75t_L g1030 ( .A(n_571), .Y(n_1030) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g657 ( .A(n_578), .Y(n_657) );
BUFx4f_ASAP7_75t_SL g699 ( .A(n_578), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_587), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .Y(n_581) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g871 ( .A(n_584), .Y(n_871) );
INVx1_ASAP7_75t_L g1105 ( .A(n_585), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_593), .Y(n_587) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g639 ( .A(n_590), .Y(n_639) );
INVx3_ASAP7_75t_L g674 ( .A(n_590), .Y(n_674) );
INVx2_ASAP7_75t_L g734 ( .A(n_590), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_590), .A2(n_877), .B1(n_878), .B2(n_879), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_590), .A2(n_1103), .B1(n_1104), .B2(n_1105), .Y(n_1102) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
XOR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_621), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_609), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_603), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVx1_ASAP7_75t_SL g855 ( .A(n_601), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_615), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g842 ( .A(n_619), .Y(n_842) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g626 ( .A(n_627), .B(n_641), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_628), .B(n_635), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g685 ( .A(n_633), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_642), .B(n_651), .Y(n_641) );
OAI222xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_647), .B2(n_648), .C1(n_649), .C2(n_650), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g854 ( .A1(n_643), .A2(n_855), .B1(n_856), .B2(n_857), .C(n_858), .Y(n_854) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx6f_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g1089 ( .A(n_650), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_656), .Y(n_651) );
INVx2_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_808), .B1(n_882), .B2(n_883), .Y(n_661) );
INVx1_ASAP7_75t_L g882 ( .A(n_662), .Y(n_882) );
XNOR2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_743), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_690), .B2(n_742), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g689 ( .A(n_668), .Y(n_689) );
NAND4xp75_ASAP7_75t_L g668 ( .A(n_669), .B(n_676), .C(n_680), .D(n_687), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .Y(n_669) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g778 ( .A(n_685), .Y(n_778) );
BUFx6f_ASAP7_75t_L g896 ( .A(n_685), .Y(n_896) );
INVx1_ASAP7_75t_L g742 ( .A(n_690), .Y(n_742) );
AO22x2_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B1(n_712), .B2(n_713), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g710 ( .A(n_693), .Y(n_710) );
OR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_703), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .C(n_701), .D(n_702), .Y(n_694) );
INVx3_ASAP7_75t_L g940 ( .A(n_696), .Y(n_940) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .C(n_706), .D(n_708), .Y(n_703) );
AO22x2_ASAP7_75t_SL g907 ( .A1(n_712), .A2(n_713), .B1(n_908), .B2(n_929), .Y(n_907) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_727), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_722), .C(n_724), .Y(n_715) );
NOR4xp25_ASAP7_75t_L g740 ( .A(n_716), .B(n_728), .C(n_732), .D(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_720), .Y(n_716) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx3_ASAP7_75t_L g859 ( .A(n_719), .Y(n_859) );
INVx2_ASAP7_75t_L g904 ( .A(n_719), .Y(n_904) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_723), .B(n_725), .Y(n_741) );
INVxp67_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_732), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_736), .Y(n_1099) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OA22x2_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_760), .B1(n_806), .B2(n_807), .Y(n_743) );
HB1xp67_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g806 ( .A(n_745), .Y(n_806) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NOR2xp67_ASAP7_75t_L g747 ( .A(n_748), .B(n_753), .Y(n_747) );
NAND4xp25_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .C(n_751), .D(n_752), .Y(n_748) );
NAND4xp25_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .C(n_756), .D(n_758), .Y(n_753) );
INVx2_ASAP7_75t_L g807 ( .A(n_760), .Y(n_807) );
AO22x2_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_785), .B1(n_803), .B2(n_804), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AND2x4_ASAP7_75t_L g764 ( .A(n_765), .B(n_774), .Y(n_764) );
NOR2xp67_ASAP7_75t_L g765 ( .A(n_766), .B(n_771), .Y(n_765) );
OAI21xp5_ASAP7_75t_SL g766 ( .A1(n_767), .A2(n_769), .B(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
NOR2x1_ASAP7_75t_L g774 ( .A(n_775), .B(n_781), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_779), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g867 ( .A(n_778), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVx2_ASAP7_75t_L g803 ( .A(n_785), .Y(n_803) );
NAND4xp25_ASAP7_75t_SL g786 ( .A(n_787), .B(n_791), .C(n_795), .D(n_798), .Y(n_786) );
AND4x1_ASAP7_75t_L g801 ( .A(n_787), .B(n_791), .C(n_795), .D(n_798), .Y(n_801) );
AND2x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_794), .Y(n_791) );
AND2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
AO22x2_ASAP7_75t_L g810 ( .A1(n_803), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_803), .Y(n_811) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g883 ( .A(n_808), .Y(n_883) );
AO22x1_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B1(n_850), .B2(n_881), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
OA22x2_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_835), .B2(n_836), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_818), .B(n_825), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_824), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_830), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_833), .Y(n_830) );
INVx1_ASAP7_75t_SL g835 ( .A(n_836), .Y(n_835) );
NOR2x1_ASAP7_75t_L g837 ( .A(n_838), .B(n_845), .Y(n_837) );
NAND4xp25_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .C(n_843), .D(n_844), .Y(n_838) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NAND4xp25_ASAP7_75t_SL g845 ( .A(n_846), .B(n_847), .C(n_848), .D(n_849), .Y(n_845) );
INVx1_ASAP7_75t_L g881 ( .A(n_850), .Y(n_881) );
INVx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
AND3x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_863), .C(n_873), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_860), .Y(n_853) );
OAI21xp33_ASAP7_75t_L g917 ( .A1(n_855), .A2(n_918), .B(n_919), .Y(n_917) );
BUFx6f_ASAP7_75t_L g1027 ( .A(n_859), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_864), .B(n_869), .Y(n_863) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx3_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g1049 ( .A(n_884), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_931), .B1(n_1036), .B2(n_1037), .Y(n_884) );
INVx1_ASAP7_75t_L g1036 ( .A(n_885), .Y(n_1036) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OA21x2_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_907), .B(n_930), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_887), .B(n_907), .Y(n_930) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_888), .A2(n_933), .B1(n_957), .B2(n_958), .Y(n_932) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
NOR2x1_ASAP7_75t_L g891 ( .A(n_892), .B(n_899), .Y(n_891) );
NAND4xp25_ASAP7_75t_SL g892 ( .A(n_893), .B(n_894), .C(n_895), .D(n_897), .Y(n_892) );
NAND4xp25_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .C(n_903), .D(n_905), .Y(n_899) );
INVx2_ASAP7_75t_L g929 ( .A(n_908), .Y(n_929) );
OAI21x1_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_910), .B(n_928), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_909), .B(n_912), .Y(n_928) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_920), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_914), .B(n_917), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_925), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_924), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
INVx1_ASAP7_75t_SL g1037 ( .A(n_931), .Y(n_1037) );
OA22x2_ASAP7_75t_L g931 ( .A1(n_932), .A2(n_959), .B1(n_960), .B2(n_1035), .Y(n_931) );
INVx1_ASAP7_75t_L g1035 ( .A(n_932), .Y(n_1035) );
INVx3_ASAP7_75t_L g957 ( .A(n_933), .Y(n_957) );
XOR2x2_ASAP7_75t_L g933 ( .A(n_934), .B(n_956), .Y(n_933) );
NAND2xp5_ASAP7_75t_SL g934 ( .A(n_935), .B(n_947), .Y(n_934) );
NOR2x1_ASAP7_75t_L g935 ( .A(n_936), .B(n_944), .Y(n_935) );
OAI222xp33_ASAP7_75t_L g936 ( .A1(n_937), .A2(n_939), .B1(n_940), .B2(n_941), .C1(n_942), .C2(n_943), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g1084 ( .A1(n_940), .A2(n_1085), .B1(n_1086), .B2(n_1087), .C(n_1088), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_948), .B(n_952), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_953), .B(n_955), .Y(n_952) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
AOI22x1_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_1012), .B1(n_1013), .B2(n_1034), .Y(n_960) );
INVx2_ASAP7_75t_L g1034 ( .A(n_961), .Y(n_1034) );
XNOR2x1_ASAP7_75t_L g961 ( .A(n_962), .B(n_999), .Y(n_961) );
OAI21xp5_ASAP7_75t_L g962 ( .A1(n_963), .A2(n_979), .B(n_997), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_963), .B(n_998), .Y(n_997) );
XNOR2x1_ASAP7_75t_L g963 ( .A(n_964), .B(n_965), .Y(n_963) );
AND2x2_ASAP7_75t_L g965 ( .A(n_966), .B(n_972), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_969), .B(n_970), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g972 ( .A(n_973), .B(n_976), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_977), .B(n_978), .Y(n_976) );
NAND2x1p5_ASAP7_75t_L g980 ( .A(n_981), .B(n_990), .Y(n_980) );
NOR2x1_ASAP7_75t_L g981 ( .A(n_982), .B(n_987), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_988), .B(n_989), .Y(n_987) );
NOR2x1_ASAP7_75t_L g990 ( .A(n_991), .B(n_994), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_993), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
XOR2x2_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1011), .Y(n_999) );
NAND4xp75_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1004), .C(n_1007), .D(n_1010), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
NOR2xp33_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1023), .Y(n_1016) );
NAND4xp25_ASAP7_75t_SL g1017 ( .A(n_1018), .B(n_1019), .C(n_1021), .D(n_1022), .Y(n_1017) );
NAND4xp25_ASAP7_75t_SL g1023 ( .A(n_1024), .B(n_1025), .C(n_1026), .D(n_1028), .Y(n_1023) );
BUFx3_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
BUFx6f_ASAP7_75t_SL g1031 ( .A(n_1032), .Y(n_1031) );
INVx2_ASAP7_75t_SL g1038 ( .A(n_1039), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1043), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1040), .B(n_1044), .Y(n_1116) );
NOR2xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1042), .Y(n_1054) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1047), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1050), .Y(n_1048) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
NOR2x1_ASAP7_75t_R g1053 ( .A(n_1054), .B(n_1055), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1054), .B(n_1056), .Y(n_1117) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
NOR2xp33_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1058), .Y(n_1056) );
OAI222xp33_ASAP7_75t_R g1060 ( .A1(n_1061), .A2(n_1077), .B1(n_1079), .B2(n_1113), .C1(n_1114), .C2(n_1117), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g1076 ( .A(n_1062), .Y(n_1076) );
INVxp33_ASAP7_75t_SL g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_SL g1063 ( .A(n_1064), .Y(n_1063) );
NOR2x1_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1070), .Y(n_1064) );
NAND4xp25_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .C(n_1068), .D(n_1069), .Y(n_1065) );
NAND4xp25_ASAP7_75t_SL g1070 ( .A(n_1071), .B(n_1072), .C(n_1073), .D(n_1074), .Y(n_1070) );
INVx1_ASAP7_75t_SL g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
XNOR2x1_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1113), .Y(n_1081) );
NAND4xp75_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1090), .C(n_1101), .D(n_1110), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
NOR2x1_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1096), .Y(n_1090) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
NOR2x1_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1106), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1112), .Y(n_1110) );
CKINVDCx20_ASAP7_75t_R g1114 ( .A(n_1115), .Y(n_1114) );
CKINVDCx6p67_ASAP7_75t_R g1115 ( .A(n_1116), .Y(n_1115) );
endmodule