module fake_netlist_6_3697_n_447 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_447);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_447;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_443;
wire n_246;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_383;
wire n_200;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_222;
wire n_248;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_235;
wire n_191;
wire n_340;
wire n_387;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_156;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_197;
wire n_343;
wire n_397;
wire n_155;
wire n_445;
wire n_425;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_417;
wire n_446;
wire n_374;
wire n_366;
wire n_407;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_265;
wire n_260;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_164;
wire n_292;
wire n_307;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_319;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_328;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_57),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_87),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_23),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_51),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_20),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_54),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_89),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_59),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_44),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_38),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_62),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_101),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_56),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_43),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_36),
.B(n_13),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_92),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_53),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_120),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_73),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_82),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_69),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_27),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_46),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_42),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_66),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_98),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_37),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_48),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_64),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_114),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_126),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_144),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_31),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_14),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_131),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_112),
.B(n_58),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_18),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_22),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_147),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_77),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_52),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_L g211 ( 
.A(n_61),
.B(n_41),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_138),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_45),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_35),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_17),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_119),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_9),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_117),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_28),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_108),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_12),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_151),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_55),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_10),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_21),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_1),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_6),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_29),
.B(n_4),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_96),
.B(n_80),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_47),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_88),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_85),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_1),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_140),
.B(n_102),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_134),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_145),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_7),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_97),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_146),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_72),
.B(n_127),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_128),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_2),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_109),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_91),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_11),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_2),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_75),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_130),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_16),
.B(n_94),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_33),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_8),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_121),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_71),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_122),
.Y(n_258)
);

INVxp33_ASAP7_75t_SL g259 ( 
.A(n_106),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_60),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_118),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_93),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_74),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_0),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_67),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_142),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_123),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_SL g268 ( 
.A(n_187),
.B(n_230),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_267),
.B(n_0),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_185),
.A2(n_5),
.B1(n_15),
.B2(n_19),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_24),
.Y(n_272)
);

AO22x2_ASAP7_75t_L g273 ( 
.A1(n_157),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_157),
.B(n_32),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_194),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_214),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

OR2x6_ASAP7_75t_L g280 ( 
.A(n_190),
.B(n_34),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_237),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_213),
.B(n_39),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_155),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_154),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_158),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_156),
.Y(n_288)
);

OR2x6_ASAP7_75t_L g289 ( 
.A(n_216),
.B(n_40),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_217),
.B(n_49),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_184),
.B(n_65),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_219),
.B(n_259),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_168),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_264),
.A2(n_68),
.B1(n_70),
.B2(n_79),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_172),
.B(n_84),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_160),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_162),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_164),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_165),
.Y(n_299)
);

BUFx4f_ASAP7_75t_L g300 ( 
.A(n_169),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_170),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_167),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_174),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_175),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_166),
.A2(n_86),
.B1(n_90),
.B2(n_99),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_177),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_161),
.B(n_100),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_188),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_163),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_207),
.B(n_103),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_171),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_201),
.B(n_104),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_178),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_179),
.B(n_110),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_186),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_227),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_173),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_189),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_261),
.B(n_111),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_191),
.Y(n_320)
);

OR2x6_ASAP7_75t_L g321 ( 
.A(n_211),
.B(n_116),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_242),
.B(n_124),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_293),
.A2(n_199),
.B(n_176),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_300),
.A2(n_210),
.B(n_215),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_192),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_317),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_292),
.A2(n_262),
.B1(n_257),
.B2(n_256),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_195),
.Y(n_329)
);

NOR2x1p5_ASAP7_75t_SL g330 ( 
.A(n_272),
.B(n_196),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_290),
.A2(n_253),
.B(n_244),
.C(n_232),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_243),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_270),
.A2(n_222),
.B(n_240),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_311),
.A2(n_159),
.B(n_180),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_282),
.A2(n_275),
.B(n_281),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_231),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_280),
.A2(n_289),
.B1(n_291),
.B2(n_294),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_225),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_284),
.A2(n_221),
.B(n_197),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_280),
.A2(n_255),
.B1(n_254),
.B2(n_252),
.Y(n_341)
);

AO22x1_ASAP7_75t_L g342 ( 
.A1(n_274),
.A2(n_220),
.B1(n_224),
.B2(n_202),
.Y(n_342)
);

AO22x1_ASAP7_75t_L g343 ( 
.A1(n_274),
.A2(n_238),
.B1(n_181),
.B2(n_266),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_319),
.A2(n_233),
.B(n_204),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_268),
.A2(n_218),
.B(n_263),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_285),
.A2(n_265),
.B(n_260),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_322),
.A2(n_209),
.B(n_247),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_299),
.A2(n_245),
.B(n_241),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_308),
.B(n_251),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_277),
.B(n_235),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_304),
.A2(n_234),
.B(n_229),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_279),
.B(n_228),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_306),
.A2(n_200),
.B(n_226),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_289),
.A2(n_249),
.B1(n_248),
.B2(n_239),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_314),
.B(n_193),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_316),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_341),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_357),
.B(n_269),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_315),
.Y(n_360)
);

O2A1O1Ixp33_ASAP7_75t_L g361 ( 
.A1(n_331),
.A2(n_298),
.B(n_287),
.C(n_318),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_339),
.A2(n_312),
.B(n_307),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_326),
.Y(n_364)
);

INVx3_ASAP7_75t_SL g365 ( 
.A(n_353),
.Y(n_365)
);

NAND2x1p5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_271),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_340),
.A2(n_274),
.B1(n_273),
.B2(n_321),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_323),
.A2(n_301),
.B(n_295),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_325),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_327),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_334),
.A2(n_310),
.B(n_277),
.Y(n_372)
);

OAI321xp33_ASAP7_75t_L g373 ( 
.A1(n_333),
.A2(n_337),
.A3(n_347),
.B1(n_321),
.B2(n_332),
.C(n_329),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_335),
.C(n_349),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_350),
.Y(n_375)
);

NAND2x1p5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_313),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_355),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_344),
.A2(n_320),
.B(n_297),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_316),
.Y(n_381)
);

O2A1O1Ixp33_ASAP7_75t_L g382 ( 
.A1(n_324),
.A2(n_303),
.B(n_345),
.C(n_354),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_342),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_203),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

OAI21x1_ASAP7_75t_L g386 ( 
.A1(n_382),
.A2(n_351),
.B(n_348),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_223),
.Y(n_388)
);

OR2x6_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_305),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_360),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_381),
.Y(n_393)
);

BUFx12f_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_379),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_212),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_380),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

NAND4xp25_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_358),
.C(n_374),
.D(n_367),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_397),
.B(n_371),
.Y(n_402)
);

OAI21xp33_ASAP7_75t_L g403 ( 
.A1(n_384),
.A2(n_366),
.B(n_383),
.Y(n_403)
);

OAI221xp5_ASAP7_75t_L g404 ( 
.A1(n_389),
.A2(n_393),
.B1(n_385),
.B2(n_390),
.C(n_396),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_399),
.A2(n_365),
.B1(n_362),
.B2(n_375),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_400),
.B(n_368),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_388),
.B(n_373),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_400),
.B(n_208),
.Y(n_408)
);

OAI21xp33_ASAP7_75t_SL g409 ( 
.A1(n_385),
.A2(n_372),
.B(n_205),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_395),
.A2(n_198),
.B1(n_206),
.B2(n_183),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_398),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_406),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_391),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_404),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_405),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_403),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_390),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_407),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_410),
.B(n_395),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_418),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_411),
.B(n_417),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_413),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_416),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_417),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_414),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_389),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_394),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_419),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_423),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_426),
.A2(n_409),
.B(n_415),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_425),
.B(n_386),
.Y(n_431)
);

NOR3xp33_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_422),
.C(n_424),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_431),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_432),
.A2(n_429),
.B1(n_428),
.B2(n_420),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_431),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_431),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_431),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_435),
.Y(n_438)
);

NAND3x1_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_387),
.C(n_136),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_436),
.Y(n_440)
);

OR2x6_ASAP7_75t_L g441 ( 
.A(n_439),
.B(n_437),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_125),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_441),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_442),
.A2(n_433),
.B(n_440),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_141),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_444),
.Y(n_446)
);

OAI221xp5_ASAP7_75t_R g447 ( 
.A1(n_445),
.A2(n_446),
.B1(n_153),
.B2(n_143),
.C(n_182),
.Y(n_447)
);


endmodule