module fake_jpeg_7055_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_1),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx14_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

AND2x2_ASAP7_75t_SL g13 ( 
.A(n_1),
.B(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_13),
.A2(n_0),
.B(n_1),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_16),
.A2(n_20),
.B(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g17 ( 
.A(n_13),
.Y(n_17)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_2),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_2),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_6),
.Y(n_23)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_17),
.B(n_24),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_11),
.A2(n_15),
.B(n_8),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_23),
.C(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_30),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.C(n_29),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_26),
.B1(n_17),
.B2(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_38),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_33),
.B1(n_30),
.B2(n_27),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_31),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_37),
.C(n_39),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_35),
.B(n_40),
.Y(n_43)
);


endmodule