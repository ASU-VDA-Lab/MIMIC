module fake_netlist_5_2145_n_20 (n_8, n_4, n_5, n_7, n_0, n_2, n_3, n_6, n_1, n_20);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_2;
input n_3;
input n_6;
input n_1;

output n_20;

wire n_16;
wire n_12;
wire n_9;
wire n_18;
wire n_10;
wire n_11;
wire n_17;
wire n_19;
wire n_15;
wire n_14;
wire n_13;

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

OAI22xp33_ASAP7_75t_L g10 ( 
.A1(n_4),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_10)
);

INVxp67_ASAP7_75t_SL g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

AO31x2_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_0),
.A3(n_1),
.B(n_2),
.Y(n_13)
);

NOR2x1_ASAP7_75t_L g14 ( 
.A(n_13),
.B(n_12),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NAND3xp33_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_15),
.C(n_9),
.Y(n_17)
);

AOI221xp5_ASAP7_75t_SL g18 ( 
.A1(n_16),
.A2(n_10),
.B1(n_13),
.B2(n_2),
.C(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

OR2x6_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_18),
.Y(n_20)
);


endmodule