module fake_jpeg_18062_n_355 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_47),
.Y(n_81)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_63),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_57),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_24),
.B1(n_30),
.B2(n_34),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_32),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_61),
.Y(n_88)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx2_ASAP7_75t_SL g97 ( 
.A(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_35),
.B1(n_26),
.B2(n_33),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_23),
.C(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_68),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_23),
.C(n_32),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_82),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_35),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_95),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_26),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_27),
.B1(n_77),
.B2(n_66),
.Y(n_129)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_33),
.Y(n_106)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_71),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_31),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_31),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp33_ASAP7_75t_R g111 ( 
.A(n_57),
.B(n_18),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_65),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_85),
.B1(n_111),
.B2(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_113),
.A2(n_139),
.B1(n_108),
.B2(n_91),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_123),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_127),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_124),
.B(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_97),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_68),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_74),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_31),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_85),
.C(n_100),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_17),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_92),
.B(n_72),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_86),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_138),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_86),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_85),
.A2(n_79),
.B1(n_66),
.B2(n_45),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_95),
.A2(n_77),
.B1(n_62),
.B2(n_79),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_84),
.B1(n_110),
.B2(n_103),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_90),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_94),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_153),
.B1(n_156),
.B2(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_90),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_98),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_154),
.B(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_106),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_17),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_105),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_161),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_122),
.B1(n_127),
.B2(n_124),
.Y(n_169)
);

AO22x2_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_78),
.B1(n_102),
.B2(n_104),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_103),
.B1(n_142),
.B2(n_126),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_99),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_67),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_81),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_136),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_170),
.B1(n_175),
.B2(n_176),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_122),
.B1(n_132),
.B2(n_113),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_145),
.B1(n_149),
.B2(n_148),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_167),
.B1(n_164),
.B2(n_144),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_116),
.B1(n_121),
.B2(n_133),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_165),
.A2(n_117),
.B1(n_130),
.B2(n_84),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_182),
.B1(n_183),
.B2(n_188),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_186),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_130),
.B1(n_118),
.B2(n_131),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_118),
.B1(n_126),
.B2(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_158),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_87),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_156),
.C(n_67),
.Y(n_216)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_93),
.B1(n_87),
.B2(n_128),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_146),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_27),
.B(n_18),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_191),
.B(n_166),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_152),
.A2(n_34),
.B1(n_36),
.B2(n_40),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_145),
.B1(n_154),
.B2(n_159),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_199),
.B1(n_204),
.B2(n_208),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_155),
.Y(n_196)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_176),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_198),
.B(n_209),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_173),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_169),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_216),
.C(n_191),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_152),
.B1(n_150),
.B2(n_157),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_180),
.B(n_143),
.Y(n_209)
);

AND2x6_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_183),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_214),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_174),
.A2(n_147),
.B1(n_151),
.B2(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_162),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_221),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_162),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_163),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_230),
.C(n_200),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_224),
.B(n_236),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_182),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_194),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_239),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_206),
.A2(n_189),
.B(n_184),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_238),
.A2(n_212),
.B(n_214),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_194),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_199),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_231),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_192),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_246),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_208),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_268),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_258),
.B(n_260),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_205),
.B(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_201),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_256),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_243),
.A2(n_206),
.B(n_210),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_225),
.A2(n_200),
.B(n_184),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_226),
.A2(n_204),
.B1(n_216),
.B2(n_193),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_249),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_193),
.B(n_101),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_226),
.A2(n_125),
.B1(n_101),
.B2(n_36),
.Y(n_264)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_236),
.B(n_19),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_41),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_244),
.B1(n_231),
.B2(n_239),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_223),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_270),
.A2(n_223),
.B1(n_240),
.B2(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

AOI21x1_ASAP7_75t_SL g305 ( 
.A1(n_274),
.A2(n_6),
.B(n_8),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_222),
.C(n_230),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_286),
.C(n_290),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_278),
.B1(n_284),
.B2(n_285),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_260),
.A2(n_227),
.B1(n_238),
.B2(n_233),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_242),
.B1(n_224),
.B2(n_247),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_288),
.B1(n_289),
.B2(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_228),
.B1(n_36),
.B2(n_3),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_59),
.C(n_49),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_41),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_259),
.C(n_254),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_262),
.C(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_294),
.B(n_296),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_261),
.C(n_266),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_273),
.A2(n_251),
.B(n_250),
.C(n_269),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_301),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_279),
.A2(n_248),
.B1(n_250),
.B2(n_264),
.Y(n_299)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_59),
.C(n_25),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_286),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_282),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_303),
.A2(n_305),
.B1(n_288),
.B2(n_281),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_19),
.C(n_25),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_306),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_8),
.B(n_10),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_304),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_273),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_316),
.C(n_318),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_278),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_315),
.B(n_319),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_274),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_317),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_271),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_305),
.A2(n_287),
.B1(n_10),
.B2(n_11),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_292),
.A2(n_8),
.B(n_10),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_293),
.Y(n_321)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_316),
.Y(n_322)
);

AND2x2_ASAP7_75t_SL g340 ( 
.A(n_322),
.B(n_326),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_325),
.Y(n_336)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_297),
.B(n_298),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_327),
.A2(n_332),
.B(n_20),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_300),
.Y(n_329)
);

AOI21xp33_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_11),
.B(n_12),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_313),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_331),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_302),
.C(n_300),
.Y(n_332)
);

AOI221xp5_ASAP7_75t_L g333 ( 
.A1(n_323),
.A2(n_311),
.B1(n_309),
.B2(n_314),
.C(n_15),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_333),
.A2(n_334),
.B1(n_14),
.B2(n_18),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_20),
.C(n_18),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_330),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_339),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_324),
.B(n_322),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_341),
.A2(n_342),
.B(n_336),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_340),
.A2(n_328),
.B(n_331),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_344),
.Y(n_348)
);

O2A1O1Ixp5_ASAP7_75t_L g345 ( 
.A1(n_333),
.A2(n_21),
.B(n_28),
.C(n_337),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_345),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_347),
.Y(n_350)
);

NAND4xp25_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_349),
.C(n_348),
.D(n_346),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_351),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_21),
.B(n_28),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_21),
.C(n_28),
.Y(n_354)
);

AO21x1_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_21),
.B(n_28),
.Y(n_355)
);


endmodule