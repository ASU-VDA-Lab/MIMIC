module fake_jpeg_22484_n_220 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_31),
.B1(n_27),
.B2(n_29),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_1),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_61),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_64),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_29),
.B1(n_27),
.B2(n_33),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_62),
.B1(n_25),
.B2(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_31),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_57),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_31),
.B1(n_27),
.B2(n_19),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_59),
.B1(n_32),
.B2(n_28),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_33),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_25),
.B1(n_23),
.B2(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_25),
.B1(n_20),
.B2(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_33),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_67),
.Y(n_89)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_16),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_76),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_78),
.A2(n_90),
.B1(n_101),
.B2(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_21),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_80),
.B(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_21),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_23),
.C(n_19),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_79),
.Y(n_106)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_94),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

BUFx4f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_98),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_21),
.B1(n_20),
.B2(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_30),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_32),
.B1(n_26),
.B2(n_17),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_30),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_1),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_26),
.B(n_16),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_24),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_16),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_16),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_107),
.Y(n_140)
);

XNOR2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_81),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_97),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_1),
.Y(n_147)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_114),
.B1(n_124),
.B2(n_97),
.Y(n_145)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_92),
.Y(n_133)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_120),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_78),
.B1(n_76),
.B2(n_80),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_83),
.Y(n_134)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_46),
.B1(n_65),
.B2(n_52),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_89),
.A2(n_65),
.B1(n_16),
.B2(n_14),
.Y(n_127)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_133),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_81),
.C(n_72),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_149),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_114),
.B1(n_122),
.B2(n_126),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_88),
.C(n_87),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_88),
.B(n_77),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_118),
.B1(n_117),
.B2(n_116),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_145),
.B1(n_127),
.B2(n_134),
.C(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_112),
.B(n_98),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_148),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_146),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_128),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_112),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_158),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_131),
.B(n_117),
.C(n_12),
.D(n_84),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_131),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_147),
.A3(n_138),
.B1(n_144),
.B2(n_143),
.C1(n_148),
.C2(n_150),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_74),
.B1(n_103),
.B2(n_90),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_173),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_143),
.B1(n_136),
.B2(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_154),
.A2(n_147),
.B(n_135),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_177),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_180),
.C(n_139),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_149),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_135),
.B(n_113),
.Y(n_181)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_153),
.C(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_178),
.C(n_175),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_153),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_187),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_159),
.A3(n_161),
.B1(n_155),
.B2(n_160),
.C1(n_156),
.C2(n_12),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_185),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_191),
.B(n_176),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_199),
.B1(n_189),
.B2(n_184),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_196),
.C(n_201),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_188),
.A2(n_174),
.B1(n_175),
.B2(n_163),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_192),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_190),
.B(n_120),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_129),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_187),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_206),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_204),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_182),
.C(n_183),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_207),
.C(n_2),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_123),
.C(n_3),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_197),
.A3(n_198),
.B1(n_199),
.B2(n_5),
.C1(n_7),
.C2(n_2),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_2),
.B(n_3),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_214),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_3),
.B(n_4),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_213),
.A2(n_209),
.B(n_8),
.C(n_9),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_215),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_9),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_9),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_218),
.Y(n_220)
);


endmodule