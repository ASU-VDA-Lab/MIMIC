module fake_netlist_6_3353_n_1776 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1776);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1776;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_39),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_29),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_57),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_61),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_39),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_12),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_123),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_29),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_58),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_54),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_71),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_20),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_1),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_21),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_24),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_161),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_77),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_31),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_5),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_27),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_128),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_115),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_84),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_31),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_43),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_26),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_34),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_7),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_42),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_40),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_73),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_109),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_69),
.Y(n_203)
);

BUFx8_ASAP7_75t_SL g204 ( 
.A(n_59),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_129),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_116),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_145),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_82),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_2),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_0),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_24),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_138),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_94),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_64),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_86),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_4),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_33),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_12),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_18),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_50),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_105),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_30),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_97),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_87),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_99),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_112),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_139),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_41),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_108),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_66),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_18),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_41),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_16),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_133),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_49),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_22),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_16),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_72),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_38),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_151),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_36),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_23),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_2),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_65),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_19),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_154),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_44),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_78),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_101),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_22),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_30),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_79),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_91),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_159),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_141),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_48),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_140),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_149),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_137),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_0),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_21),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_132),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_98),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_38),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_150),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_134),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_60),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_135),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_63),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_15),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_81),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_40),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_23),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_74),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_131),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_158),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_100),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_26),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_51),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_52),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_120),
.Y(n_288)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_146),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_62),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_55),
.Y(n_291)
);

BUFx8_ASAP7_75t_SL g292 ( 
.A(n_126),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_14),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_36),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_117),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_4),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_37),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_142),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_8),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_34),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_5),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_144),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_1),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_122),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_6),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_19),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_43),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_68),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_14),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_111),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_56),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_92),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_28),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_136),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_17),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_127),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_44),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_110),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_130),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_162),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_35),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_11),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_46),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_171),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_170),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_170),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_170),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_168),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_204),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_170),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_292),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_164),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_166),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_170),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_252),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_215),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_252),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_252),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_172),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_180),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_252),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_188),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_173),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_180),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_280),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_280),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_187),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_258),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_187),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_189),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_260),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_244),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_168),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_181),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_235),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_182),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_232),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_296),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_260),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_193),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_190),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_195),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_182),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_198),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_211),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_258),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_219),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_220),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_191),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_225),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_238),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_241),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_232),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_272),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_272),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_242),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_185),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_247),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_169),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_201),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_202),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_169),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_203),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_299),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_299),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_281),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_289),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_281),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_214),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_214),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_283),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_295),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_205),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_259),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_353),
.B(n_231),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_325),
.B(n_206),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_231),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_327),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_333),
.B(n_206),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_336),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_R g416 ( 
.A(n_329),
.B(n_283),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_328),
.A2(n_199),
.B1(n_297),
.B2(n_294),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_334),
.B(n_249),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_341),
.B(n_249),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_359),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_339),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_340),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_354),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_347),
.B(n_262),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_343),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_356),
.B(n_262),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_367),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_348),
.A2(n_256),
.B1(n_199),
.B2(n_297),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_396),
.A2(n_308),
.B(n_295),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_324),
.A2(n_256),
.B1(n_279),
.B2(n_294),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_344),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_363),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_345),
.B(n_346),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_345),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_346),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_372),
.B(n_231),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_375),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_350),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_350),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_351),
.B(n_287),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_351),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_396),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_397),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_337),
.A2(n_279),
.B1(n_304),
.B2(n_185),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_399),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_388),
.B(n_287),
.Y(n_460)
);

CKINVDCx6p67_ASAP7_75t_R g461 ( 
.A(n_381),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_379),
.A2(n_321),
.B1(n_322),
.B2(n_304),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_390),
.B(n_308),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_372),
.B(n_175),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_366),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_366),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_330),
.B(n_364),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_400),
.B(n_167),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_361),
.B(n_178),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_380),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_332),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_330),
.B(n_174),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_342),
.B(n_300),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_352),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_409),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_409),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_468),
.Y(n_478)
);

OR2x6_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_177),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_445),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_428),
.B(n_401),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

INVx6_ASAP7_75t_L g483 ( 
.A(n_417),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_464),
.A2(n_383),
.B1(n_349),
.B2(n_378),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_445),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_404),
.A2(n_374),
.B1(n_376),
.B2(n_377),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_411),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_207),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_404),
.B(n_370),
.C(n_368),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_425),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_417),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

INVx8_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_417),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_428),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_425),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

BUFx6f_ASAP7_75t_SL g500 ( 
.A(n_404),
.Y(n_500)
);

INVxp33_ASAP7_75t_SL g501 ( 
.A(n_416),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_473),
.B(n_398),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_419),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_402),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_435),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_425),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_412),
.B(n_208),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_404),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_473),
.B(n_352),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_402),
.B(n_355),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_442),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_474),
.B(n_437),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_442),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_461),
.Y(n_516)
);

OAI22xp33_ASAP7_75t_L g517 ( 
.A1(n_458),
.A2(n_237),
.B1(n_268),
.B2(n_267),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_425),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_420),
.B(n_212),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_403),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_444),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_403),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_452),
.A2(n_360),
.B1(n_228),
.B2(n_265),
.Y(n_524)
);

INVxp33_ASAP7_75t_SL g525 ( 
.A(n_463),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_405),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_407),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_406),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_423),
.B(n_434),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

AND3x2_ASAP7_75t_L g532 ( 
.A(n_431),
.B(n_217),
.C(n_213),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_408),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_436),
.B(n_216),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_460),
.B(n_223),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_407),
.B(n_355),
.Y(n_536)
);

AND3x2_ASAP7_75t_L g537 ( 
.A(n_441),
.B(n_453),
.C(n_432),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_451),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_461),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_405),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_452),
.A2(n_228),
.B1(n_175),
.B2(n_265),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_448),
.B(n_224),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_451),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_405),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_410),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_452),
.B(n_370),
.C(n_368),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_449),
.B(n_393),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_405),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_410),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_448),
.B(n_395),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_405),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_454),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_454),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_452),
.A2(n_175),
.B1(n_265),
.B2(n_228),
.Y(n_554)
);

CKINVDCx6p67_ASAP7_75t_R g555 ( 
.A(n_443),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_458),
.B(n_386),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_415),
.B(n_229),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_405),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_463),
.B(n_163),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_413),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_443),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_415),
.Y(n_563)
);

BUFx8_ASAP7_75t_SL g564 ( 
.A(n_472),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_427),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_427),
.B(n_230),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_424),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_440),
.B(n_176),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_430),
.B(n_240),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_455),
.B(n_386),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_430),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_413),
.Y(n_572)
);

CKINVDCx6p67_ASAP7_75t_R g573 ( 
.A(n_465),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_433),
.B(n_245),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_433),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_447),
.B(n_253),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_440),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_447),
.B(n_254),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_438),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_439),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_439),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_413),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_413),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_439),
.A2(n_175),
.B1(n_228),
.B2(n_265),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_438),
.B(n_176),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_466),
.B(n_392),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_466),
.B(n_371),
.C(n_385),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_413),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_418),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_413),
.B(n_257),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_455),
.B(n_357),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_414),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_414),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_465),
.B(n_175),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_467),
.Y(n_595)
);

BUFx8_ASAP7_75t_SL g596 ( 
.A(n_418),
.Y(n_596)
);

INVxp67_ASAP7_75t_SL g597 ( 
.A(n_414),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_414),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_456),
.B(n_389),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_467),
.B(n_183),
.Y(n_600)
);

AO22x2_ASAP7_75t_L g601 ( 
.A1(n_456),
.A2(n_234),
.B1(n_222),
.B2(n_226),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_465),
.B(n_300),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_414),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_459),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_457),
.B(n_389),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_457),
.B(n_183),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_459),
.B(n_184),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_465),
.B(n_184),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_414),
.B(n_261),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_421),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_421),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_475),
.B(n_462),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_475),
.B(n_391),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_421),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_462),
.A2(n_236),
.B1(n_165),
.B2(n_323),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_421),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_421),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_421),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_465),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_422),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_422),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_422),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_422),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_422),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_529),
.B(n_422),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_481),
.B(n_179),
.Y(n_626)
);

BUFx6f_ASAP7_75t_SL g627 ( 
.A(n_479),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_511),
.B(n_391),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_510),
.A2(n_286),
.B1(n_273),
.B2(n_263),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_511),
.B(n_392),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_581),
.Y(n_631)
);

O2A1O1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_586),
.A2(n_371),
.B(n_385),
.C(n_384),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_481),
.B(n_186),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_497),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_480),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_510),
.B(n_227),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_483),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_595),
.B(n_426),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_595),
.B(n_426),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_571),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_480),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_482),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_581),
.A2(n_465),
.B1(n_265),
.B2(n_228),
.Y(n_643)
);

O2A1O1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_586),
.A2(n_373),
.B(n_384),
.C(n_382),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_497),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_491),
.B(n_426),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_512),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_478),
.B(n_373),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_491),
.B(n_426),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_525),
.A2(n_239),
.B1(n_310),
.B2(n_243),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_575),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_494),
.B(n_496),
.Y(n_652)
);

XNOR2x2_ASAP7_75t_SL g653 ( 
.A(n_556),
.B(n_382),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_482),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_512),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_494),
.B(n_426),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_575),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_478),
.B(n_192),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_567),
.B(n_251),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_L g660 ( 
.A(n_584),
.B(n_289),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_485),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_567),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_499),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_485),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_505),
.B(n_426),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_536),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_505),
.B(n_289),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_612),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_619),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_502),
.B(n_194),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_536),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_499),
.B(n_365),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_527),
.B(n_196),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_527),
.B(n_429),
.Y(n_674)
);

AOI221xp5_ASAP7_75t_L g675 ( 
.A1(n_517),
.A2(n_218),
.B1(n_210),
.B2(n_209),
.C(n_200),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_L g676 ( 
.A(n_495),
.B(n_289),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_604),
.B(n_429),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_619),
.B(n_289),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_532),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_591),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_479),
.A2(n_500),
.B1(n_503),
.B2(n_488),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_580),
.B(n_289),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_604),
.B(n_429),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_490),
.B(n_429),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_580),
.B(n_602),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_602),
.B(n_289),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_498),
.B(n_429),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_521),
.B(n_429),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_556),
.B(n_577),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_541),
.B(n_276),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_479),
.A2(n_290),
.B1(n_319),
.B2(n_221),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_550),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_568),
.B(n_197),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_591),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_479),
.A2(n_312),
.B1(n_288),
.B2(n_264),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_612),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_518),
.B(n_266),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_518),
.B(n_269),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_521),
.B(n_446),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_523),
.B(n_446),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_523),
.B(n_446),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_518),
.B(n_270),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_528),
.B(n_446),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_542),
.Y(n_704)
);

AND2x2_ASAP7_75t_SL g705 ( 
.A(n_524),
.B(n_446),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_585),
.B(n_271),
.C(n_255),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_530),
.B(n_446),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_479),
.B(n_233),
.Y(n_708)
);

OR2x2_ASAP7_75t_SL g709 ( 
.A(n_525),
.B(n_365),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_SL g710 ( 
.A(n_589),
.B(n_315),
.C(n_250),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_509),
.B(n_274),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_519),
.B(n_275),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_500),
.A2(n_302),
.B1(n_320),
.B2(n_318),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_530),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_531),
.B(n_450),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_483),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_579),
.B(n_317),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_495),
.B(n_298),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_531),
.B(n_450),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_533),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_495),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_534),
.B(n_301),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_533),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_545),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_545),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_535),
.B(n_311),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_483),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_500),
.A2(n_316),
.B1(n_314),
.B2(n_278),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_547),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_562),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_615),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_L g732 ( 
.A(n_495),
.B(n_291),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_549),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_549),
.B(n_450),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_563),
.B(n_450),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_565),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_L g737 ( 
.A(n_561),
.B(n_282),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_565),
.B(n_450),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_483),
.B(n_284),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_557),
.B(n_313),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_484),
.B(n_293),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_562),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_476),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_477),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_514),
.B(n_309),
.Y(n_745)
);

O2A1O1Ixp5_ASAP7_75t_L g746 ( 
.A1(n_566),
.A2(n_307),
.B(n_306),
.C(n_303),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_608),
.B(n_285),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_569),
.B(n_277),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_582),
.B(n_248),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_477),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_487),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_564),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_574),
.B(n_246),
.Y(n_753)
);

O2A1O1Ixp5_ASAP7_75t_L g754 ( 
.A1(n_576),
.A2(n_75),
.B(n_153),
.C(n_152),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_582),
.B(n_67),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_487),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_588),
.B(n_70),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_578),
.B(n_597),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_600),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_570),
.B(n_3),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_588),
.B(n_156),
.Y(n_761)
);

AO221x1_ASAP7_75t_L g762 ( 
.A1(n_601),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_561),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_508),
.B(n_76),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_606),
.B(n_9),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_607),
.B(n_10),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_492),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_508),
.B(n_80),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_590),
.B(n_609),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_495),
.B(n_83),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_555),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_492),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_526),
.B(n_148),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_555),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_493),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_493),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_SL g777 ( 
.A(n_501),
.B(n_11),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_592),
.B(n_143),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_615),
.B(n_489),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_501),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_579),
.B(n_559),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_504),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_599),
.B(n_13),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_504),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_526),
.B(n_124),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_506),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_605),
.A2(n_13),
.B(n_17),
.C(n_20),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_506),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_635),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_662),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_668),
.B(n_554),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_672),
.B(n_516),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_641),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_637),
.B(n_592),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_642),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_662),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_669),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_669),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_668),
.B(n_489),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_654),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_696),
.B(n_546),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_634),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_692),
.B(n_537),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_689),
.B(n_589),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_645),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_661),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_637),
.B(n_598),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_664),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_727),
.B(n_598),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_R g810 ( 
.A(n_780),
.B(n_539),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_696),
.B(n_546),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_727),
.B(n_614),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_714),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_625),
.B(n_551),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_647),
.B(n_587),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_714),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_722),
.B(n_551),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_655),
.B(n_587),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_730),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_720),
.Y(n_820)
);

BUFx4f_ASAP7_75t_SL g821 ( 
.A(n_771),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_628),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_742),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_722),
.B(n_560),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_669),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_630),
.Y(n_826)
);

AND2x4_ASAP7_75t_SL g827 ( 
.A(n_669),
.B(n_573),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_725),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_771),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_631),
.B(n_560),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_721),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_721),
.B(n_614),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_626),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_640),
.Y(n_834)
);

NAND2x1p5_ASAP7_75t_L g835 ( 
.A(n_721),
.B(n_593),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_704),
.B(n_560),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_752),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_723),
.B(n_526),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_721),
.B(n_643),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_724),
.B(n_572),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_733),
.B(n_572),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_779),
.A2(n_624),
.B1(n_623),
.B2(n_620),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_736),
.B(n_572),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_643),
.B(n_610),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_SL g845 ( 
.A1(n_779),
.A2(n_522),
.B(n_507),
.C(n_513),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_648),
.B(n_558),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_626),
.B(n_516),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_717),
.B(n_539),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_716),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_763),
.Y(n_850)
);

AND2x6_ASAP7_75t_L g851 ( 
.A(n_769),
.B(n_611),
.Y(n_851)
);

BUFx12f_ASAP7_75t_L g852 ( 
.A(n_679),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_663),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_636),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_681),
.B(n_610),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_666),
.B(n_486),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_680),
.B(n_694),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_758),
.A2(n_544),
.B(n_548),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_716),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_651),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_671),
.B(n_613),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_751),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_651),
.B(n_611),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_657),
.B(n_622),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_SL g865 ( 
.A(n_710),
.B(n_596),
.C(n_601),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_781),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_759),
.B(n_622),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_685),
.A2(n_573),
.B1(n_601),
.B2(n_624),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_744),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_633),
.B(n_558),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_731),
.B(n_621),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_729),
.B(n_709),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_633),
.B(n_623),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_659),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_743),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_760),
.B(n_783),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_765),
.A2(n_507),
.B(n_513),
.C(n_553),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_762),
.A2(n_601),
.B1(n_515),
.B2(n_552),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_746),
.B(n_621),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_650),
.A2(n_552),
.B1(n_520),
.B2(n_522),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_743),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_705),
.B(n_620),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_659),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_658),
.Y(n_884)
);

NAND2x1p5_ASAP7_75t_L g885 ( 
.A(n_784),
.B(n_544),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_659),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_784),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_750),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_745),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_705),
.B(n_616),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_740),
.B(n_616),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_748),
.B(n_551),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_756),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_776),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_636),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_658),
.B(n_515),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_753),
.B(n_540),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_670),
.B(n_673),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_767),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_652),
.B(n_540),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_782),
.Y(n_901)
);

NOR2x1_ASAP7_75t_R g902 ( 
.A(n_741),
.B(n_520),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_650),
.A2(n_553),
.B1(n_543),
.B2(n_538),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_670),
.B(n_540),
.Y(n_904)
);

AND2x2_ASAP7_75t_SL g905 ( 
.A(n_770),
.B(n_594),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_772),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_636),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_665),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_674),
.Y(n_909)
);

BUFx12f_ASAP7_75t_L g910 ( 
.A(n_653),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_764),
.B(n_618),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_693),
.B(n_538),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_768),
.B(n_772),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_775),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_775),
.B(n_618),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_673),
.B(n_543),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_749),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_693),
.B(n_593),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_711),
.B(n_593),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_786),
.Y(n_920)
);

OAI22xp33_ASAP7_75t_L g921 ( 
.A1(n_777),
.A2(n_593),
.B1(n_548),
.B2(n_544),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_711),
.B(n_548),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_786),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_706),
.B(n_548),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_708),
.B(n_25),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_685),
.A2(n_544),
.B1(n_617),
.B2(n_603),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_712),
.B(n_618),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_712),
.B(n_618),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_788),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_788),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_677),
.Y(n_931)
);

NAND2x1p5_ASAP7_75t_L g932 ( 
.A(n_755),
.B(n_757),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_646),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_688),
.B(n_618),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_699),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_726),
.B(n_617),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_766),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_774),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_765),
.A2(n_603),
.B1(n_583),
.B2(n_617),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_683),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_700),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_726),
.B(n_617),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_638),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_639),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_649),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_773),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_749),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_656),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_701),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_785),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_703),
.B(n_617),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_667),
.B(n_682),
.Y(n_952)
);

INVx5_ASAP7_75t_L g953 ( 
.A(n_754),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_707),
.Y(n_954)
);

NAND2x1_ASAP7_75t_L g955 ( 
.A(n_715),
.B(n_603),
.Y(n_955)
);

AND2x6_ASAP7_75t_SL g956 ( 
.A(n_708),
.B(n_25),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_719),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_667),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_SL g959 ( 
.A1(n_766),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_SL g960 ( 
.A1(n_695),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_734),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_735),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_737),
.B(n_603),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_SL g964 ( 
.A(n_627),
.B(n_603),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_831),
.A2(n_732),
.B(n_718),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_831),
.A2(n_676),
.B(n_739),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_797),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_823),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_831),
.A2(n_687),
.B(n_684),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_898),
.B(n_738),
.Y(n_970)
);

INVx3_ASAP7_75t_SL g971 ( 
.A(n_837),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_937),
.A2(n_691),
.B(n_747),
.C(n_787),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_816),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_872),
.B(n_747),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_813),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_876),
.B(n_678),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_797),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_820),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_810),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_823),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_853),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_SL g982 ( 
.A(n_847),
.B(n_675),
.C(n_728),
.Y(n_982)
);

OAI22xp33_ASAP7_75t_L g983 ( 
.A1(n_833),
.A2(n_713),
.B1(n_629),
.B2(n_697),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_906),
.Y(n_984)
);

OAI22xp33_ASAP7_75t_L g985 ( 
.A1(n_884),
.A2(n_698),
.B1(n_697),
.B2(n_702),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_882),
.A2(n_678),
.B(n_686),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_945),
.B(n_698),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_945),
.B(n_702),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_918),
.A2(n_627),
.B1(n_761),
.B2(n_757),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_792),
.B(n_632),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_831),
.A2(n_778),
.B(n_761),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_SL g992 ( 
.A1(n_910),
.A2(n_644),
.B1(n_686),
.B2(n_660),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_822),
.B(n_778),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_873),
.B(n_755),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_804),
.B(n_690),
.Y(n_995)
);

AOI221x1_ASAP7_75t_L g996 ( 
.A1(n_918),
.A2(n_583),
.B1(n_690),
.B2(n_45),
.C(n_46),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_839),
.A2(n_583),
.B(n_93),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_810),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_873),
.B(n_583),
.Y(n_999)
);

OA21x2_ASAP7_75t_L g1000 ( 
.A1(n_877),
.A2(n_583),
.B(n_90),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_819),
.B(n_37),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_832),
.A2(n_96),
.B(n_118),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_826),
.B(n_89),
.Y(n_1003)
);

NOR3xp33_ASAP7_75t_SL g1004 ( 
.A(n_959),
.B(n_804),
.C(n_960),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_R g1005 ( 
.A(n_938),
.B(n_88),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_850),
.Y(n_1006)
);

NAND2x1p5_ASAP7_75t_L g1007 ( 
.A(n_797),
.B(n_102),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_889),
.B(n_85),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_937),
.B(n_42),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_805),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_866),
.B(n_45),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_850),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_925),
.A2(n_47),
.B1(n_104),
.B2(n_106),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_832),
.A2(n_119),
.B(n_47),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_839),
.A2(n_858),
.B(n_835),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_853),
.B(n_790),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_871),
.A2(n_857),
.B(n_855),
.C(n_947),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_828),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_933),
.B(n_948),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_854),
.B(n_796),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_935),
.B(n_941),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_949),
.B(n_957),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_896),
.B(n_962),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_802),
.B(n_848),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_912),
.B(n_916),
.Y(n_1025)
);

AOI221xp5_ASAP7_75t_L g1026 ( 
.A1(n_815),
.A2(n_818),
.B1(n_865),
.B2(n_871),
.C(n_800),
.Y(n_1026)
);

OAI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_856),
.A2(n_907),
.B1(n_895),
.B2(n_861),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_802),
.B(n_803),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_803),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_912),
.A2(n_917),
.B(n_958),
.C(n_952),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_815),
.B(n_818),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_875),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_908),
.B(n_909),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_835),
.A2(n_824),
.B(n_817),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_908),
.B(n_909),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_955),
.A2(n_926),
.B(n_913),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_902),
.B(n_907),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_874),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_789),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_855),
.A2(n_882),
.B(n_890),
.C(n_845),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_919),
.A2(n_922),
.B(n_892),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_793),
.B(n_795),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_814),
.A2(n_904),
.B(n_891),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_891),
.A2(n_846),
.B(n_897),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_852),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_854),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_890),
.A2(n_877),
.B(n_844),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_799),
.B(n_801),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_862),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_829),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_821),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_L g1052 ( 
.A1(n_879),
.A2(n_911),
.B(n_913),
.C(n_870),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_854),
.B(n_825),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_867),
.B(n_829),
.Y(n_1054)
);

CKINVDCx11_ASAP7_75t_R g1055 ( 
.A(n_956),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_806),
.B(n_808),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_811),
.B(n_954),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_825),
.B(n_867),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_963),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_954),
.B(n_961),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_834),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_961),
.B(n_943),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_830),
.A2(n_844),
.B(n_900),
.Y(n_1063)
);

OR2x6_ASAP7_75t_L g1064 ( 
.A(n_883),
.B(n_886),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_900),
.A2(n_812),
.B(n_794),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_794),
.A2(n_812),
.B(n_809),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_836),
.B(n_821),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_869),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_888),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_924),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_963),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_827),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_943),
.B(n_940),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_845),
.A2(n_894),
.B(n_893),
.C(n_901),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_860),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_931),
.B(n_940),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_807),
.A2(n_809),
.B(n_936),
.Y(n_1077)
);

XOR2xp5_ASAP7_75t_L g1078 ( 
.A(n_924),
.B(n_842),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_921),
.B(n_964),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_899),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_868),
.A2(n_843),
.B(n_841),
.C(n_840),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_827),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_931),
.B(n_944),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_914),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_798),
.B(n_944),
.Y(n_1085)
);

O2A1O1Ixp5_ASAP7_75t_SL g1086 ( 
.A1(n_879),
.A2(n_911),
.B(n_934),
.C(n_951),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_875),
.B(n_881),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_865),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_881),
.B(n_887),
.Y(n_1089)
);

INVx5_ASAP7_75t_L g1090 ( 
.A(n_851),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_927),
.A2(n_928),
.B(n_942),
.C(n_791),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_920),
.B(n_929),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_921),
.B(n_887),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_939),
.A2(n_905),
.B1(n_932),
.B2(n_953),
.Y(n_1094)
);

INVx5_ASAP7_75t_L g1095 ( 
.A(n_851),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_SL g1096 ( 
.A1(n_950),
.A2(n_849),
.B(n_859),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_849),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_923),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_807),
.A2(n_905),
.B(n_951),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_930),
.B(n_851),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_851),
.B(n_903),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1028),
.B(n_932),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1039),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1041),
.A2(n_1034),
.B(n_1015),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1054),
.B(n_859),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_973),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1036),
.A2(n_1077),
.B(n_1065),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1054),
.B(n_838),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1043),
.A2(n_953),
.B(n_950),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_L g1110 ( 
.A1(n_1079),
.A2(n_934),
.B(n_915),
.C(n_864),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_SL g1111 ( 
.A(n_1050),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_982),
.A2(n_851),
.B1(n_946),
.B2(n_880),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_1012),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1061),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_984),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1093),
.A2(n_953),
.B(n_946),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1046),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_966),
.A2(n_953),
.B(n_946),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_994),
.A2(n_946),
.B(n_939),
.Y(n_1119)
);

INVx3_ASAP7_75t_SL g1120 ( 
.A(n_1006),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1031),
.B(n_878),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1040),
.A2(n_863),
.B(n_864),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1025),
.A2(n_1021),
.B1(n_1022),
.B2(n_1023),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1066),
.A2(n_863),
.B(n_915),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_994),
.A2(n_885),
.B(n_880),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1063),
.A2(n_885),
.B(n_903),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1099),
.A2(n_1044),
.B(n_1086),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_979),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1097),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_997),
.A2(n_1052),
.B(n_965),
.Y(n_1131)
);

AOI211x1_ASAP7_75t_L g1132 ( 
.A1(n_1009),
.A2(n_1027),
.B(n_983),
.C(n_1021),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_998),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1048),
.A2(n_1094),
.B(n_970),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_974),
.B(n_1010),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1022),
.B(n_1048),
.Y(n_1136)
);

NOR2x1_ASAP7_75t_SL g1137 ( 
.A(n_1090),
.B(n_1095),
.Y(n_1137)
);

OAI22x1_ASAP7_75t_L g1138 ( 
.A1(n_1078),
.A2(n_1088),
.B1(n_1004),
.B2(n_1024),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_972),
.A2(n_1017),
.B(n_1026),
.C(n_995),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1047),
.A2(n_1100),
.B(n_969),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_968),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_970),
.B(n_1019),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1091),
.A2(n_1101),
.B(n_1030),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1042),
.A2(n_1056),
.B1(n_1019),
.B2(n_1026),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1098),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_975),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1057),
.B(n_976),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_999),
.A2(n_1096),
.B(n_1081),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1100),
.A2(n_991),
.B(n_1002),
.Y(n_1149)
);

AOI221x1_ASAP7_75t_L g1150 ( 
.A1(n_989),
.A2(n_1101),
.B1(n_986),
.B2(n_992),
.C(n_988),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1060),
.B(n_987),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1060),
.B(n_987),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1074),
.A2(n_1014),
.B(n_1092),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_978),
.Y(n_1154)
);

AOI221x1_ASAP7_75t_L g1155 ( 
.A1(n_988),
.A2(n_1085),
.B1(n_1011),
.B2(n_996),
.C(n_1033),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_990),
.B(n_980),
.Y(n_1156)
);

AOI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1000),
.A2(n_1092),
.B(n_993),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1051),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1089),
.A2(n_985),
.B(n_1076),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_981),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1037),
.B(n_1016),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1073),
.A2(n_1076),
.B(n_1062),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1000),
.A2(n_1073),
.B(n_1062),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1075),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1087),
.A2(n_1083),
.B(n_1097),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_1072),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_1008),
.A2(n_1003),
.B(n_1083),
.C(n_1053),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1005),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1068),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1087),
.A2(n_1035),
.B(n_1032),
.Y(n_1170)
);

INVx6_ASAP7_75t_SL g1171 ( 
.A(n_1064),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_L g1172 ( 
.A(n_1067),
.B(n_1055),
.C(n_1045),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1082),
.B(n_1072),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_SL g1174 ( 
.A1(n_1013),
.A2(n_967),
.B(n_1018),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1032),
.A2(n_1095),
.B(n_1090),
.Y(n_1175)
);

AO22x1_ASAP7_75t_L g1176 ( 
.A1(n_1069),
.A2(n_1038),
.B1(n_1046),
.B2(n_1071),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1001),
.A2(n_1058),
.B(n_1020),
.C(n_1064),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1064),
.Y(n_1178)
);

NAND2xp33_ASAP7_75t_L g1179 ( 
.A(n_1059),
.B(n_1071),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1029),
.B(n_1070),
.Y(n_1180)
);

AOI22x1_ASAP7_75t_L g1181 ( 
.A1(n_1049),
.A2(n_1080),
.B1(n_1084),
.B2(n_1007),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1084),
.B(n_1071),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1046),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1084),
.B(n_1059),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1090),
.A2(n_1095),
.B(n_977),
.C(n_1029),
.Y(n_1185)
);

AOI21xp33_ASAP7_75t_L g1186 ( 
.A1(n_1090),
.A2(n_1095),
.B(n_967),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1007),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1039),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1052),
.A2(n_1047),
.B(n_1041),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1054),
.B(n_1031),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1015),
.A2(n_1036),
.B(n_1077),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1039),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_1052),
.A2(n_1047),
.B(n_1041),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1015),
.A2(n_1036),
.B(n_1077),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1041),
.A2(n_727),
.B(n_637),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1040),
.A2(n_994),
.B(n_1063),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1199)
);

AOI221xp5_ASAP7_75t_L g1200 ( 
.A1(n_1004),
.A2(n_517),
.B1(n_525),
.B2(n_577),
.C(n_559),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1015),
.A2(n_1036),
.B(n_1077),
.Y(n_1201)
);

OAI22x1_ASAP7_75t_L g1202 ( 
.A1(n_1078),
.A2(n_589),
.B1(n_438),
.B2(n_440),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_1085),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1016),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1016),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1094),
.A2(n_996),
.A3(n_877),
.B(n_1034),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1040),
.A2(n_994),
.B(n_1063),
.Y(n_1209)
);

INVx6_ASAP7_75t_SL g1210 ( 
.A(n_1064),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1041),
.A2(n_727),
.B(n_637),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1054),
.B(n_1031),
.Y(n_1212)
);

INVx3_ASAP7_75t_SL g1213 ( 
.A(n_1006),
.Y(n_1213)
);

NOR3xp33_ASAP7_75t_SL g1214 ( 
.A(n_982),
.B(n_589),
.C(n_561),
.Y(n_1214)
);

OAI22x1_ASAP7_75t_L g1215 ( 
.A1(n_1078),
.A2(n_589),
.B1(n_438),
.B2(n_440),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1039),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1040),
.A2(n_994),
.B(n_1063),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1052),
.A2(n_1047),
.B(n_1041),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1017),
.A2(n_1074),
.B(n_1047),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_973),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1015),
.A2(n_1036),
.B(n_1077),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1050),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1025),
.B(n_1023),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1015),
.A2(n_1036),
.B(n_1077),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_999),
.A2(n_879),
.B(n_1034),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1010),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_SL g1228 ( 
.A1(n_1017),
.A2(n_1074),
.B(n_1047),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1015),
.A2(n_1036),
.B(n_1077),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_973),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1041),
.A2(n_727),
.B(n_637),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_999),
.A2(n_879),
.B(n_1034),
.Y(n_1232)
);

BUFx2_ASAP7_75t_R g1233 ( 
.A(n_971),
.Y(n_1233)
);

INVx6_ASAP7_75t_SL g1234 ( 
.A(n_1064),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1106),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1204),
.B(n_1156),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1202),
.A2(n_1215),
.B1(n_1144),
.B2(n_1200),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1103),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1115),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1201),
.A2(n_1225),
.B(n_1221),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1223),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1229),
.A2(n_1107),
.B(n_1118),
.Y(n_1243)
);

OR3x4_ASAP7_75t_SL g1244 ( 
.A(n_1160),
.B(n_1214),
.C(n_1138),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1223),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1136),
.B(n_1130),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1136),
.A2(n_1144),
.B1(n_1190),
.B2(n_1207),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1127),
.A2(n_1150),
.B(n_1148),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1104),
.A2(n_1211),
.B(n_1197),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1139),
.A2(n_1134),
.B(n_1217),
.C(n_1198),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1231),
.A2(n_1109),
.B(n_1198),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1205),
.B(n_1206),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1123),
.A2(n_1102),
.B1(n_1121),
.B2(n_1199),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1130),
.B(n_1190),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1209),
.A2(n_1217),
.B(n_1116),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1105),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_SL g1257 ( 
.A1(n_1137),
.A2(n_1174),
.B(n_1123),
.Y(n_1257)
);

AOI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1209),
.A2(n_1177),
.B(n_1219),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1131),
.A2(n_1140),
.B(n_1124),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1191),
.B(n_1212),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1188),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1143),
.A2(n_1153),
.B(n_1228),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1226),
.A2(n_1232),
.B(n_1126),
.Y(n_1263)
);

BUFx4f_ASAP7_75t_L g1264 ( 
.A(n_1120),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1165),
.A2(n_1170),
.B(n_1157),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1195),
.A2(n_1207),
.B1(n_1203),
.B2(n_1199),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1113),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1155),
.A2(n_1159),
.A3(n_1125),
.B(n_1119),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1227),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1132),
.B(n_1143),
.C(n_1161),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1175),
.A2(n_1122),
.B(n_1163),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1195),
.B(n_1203),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1117),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1122),
.A2(n_1163),
.B(n_1162),
.Y(n_1274)
);

NOR3xp33_ASAP7_75t_L g1275 ( 
.A(n_1222),
.B(n_1224),
.C(n_1176),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1189),
.A2(n_1218),
.B(n_1194),
.Y(n_1276)
);

NAND2x1p5_ASAP7_75t_L g1277 ( 
.A(n_1187),
.B(n_1129),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1110),
.A2(n_1112),
.B(n_1147),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1181),
.A2(n_1218),
.B(n_1194),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1220),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1230),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1117),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1222),
.A2(n_1224),
.B1(n_1142),
.B2(n_1135),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1142),
.A2(n_1152),
.B(n_1151),
.C(n_1114),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1169),
.B(n_1227),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1178),
.B(n_1173),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1128),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1164),
.B(n_1141),
.Y(n_1288)
);

CKINVDCx16_ASAP7_75t_R g1289 ( 
.A(n_1111),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1108),
.B(n_1216),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_1133),
.B(n_1180),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1193),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1108),
.B(n_1213),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_SL g1294 ( 
.A1(n_1186),
.A2(n_1184),
.B(n_1182),
.Y(n_1294)
);

NOR2x1_ASAP7_75t_SL g1295 ( 
.A(n_1166),
.B(n_1146),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1167),
.A2(n_1185),
.B(n_1179),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1223),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1186),
.A2(n_1145),
.B(n_1154),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1168),
.B(n_1158),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1172),
.A2(n_1173),
.B1(n_1111),
.B2(n_1166),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1184),
.B(n_1117),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1171),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1233),
.B(n_1183),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1183),
.Y(n_1304)
);

BUFx10_ASAP7_75t_L g1305 ( 
.A(n_1183),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1208),
.A2(n_1171),
.B(n_1210),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_SL g1307 ( 
.A1(n_1208),
.A2(n_1079),
.B(n_1139),
.C(n_1093),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1234),
.A2(n_1149),
.B(n_1192),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1135),
.B(n_1156),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1202),
.A2(n_959),
.B1(n_960),
.B2(n_898),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1113),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1202),
.A2(n_959),
.B1(n_960),
.B2(n_898),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1204),
.B(n_833),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1103),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_R g1317 ( 
.A(n_1128),
.B(n_837),
.Y(n_1317)
);

INVx4_ASAP7_75t_L g1318 ( 
.A(n_1223),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1159),
.A2(n_898),
.B(n_833),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1127),
.A2(n_1150),
.B(n_1148),
.Y(n_1321)
);

AND2x6_ASAP7_75t_L g1322 ( 
.A(n_1112),
.B(n_1187),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1191),
.B(n_1212),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1113),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1132),
.B(n_1176),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1204),
.A2(n_804),
.B1(n_1004),
.B2(n_692),
.Y(n_1329)
);

NAND3xp33_ASAP7_75t_L g1330 ( 
.A(n_1200),
.B(n_898),
.C(n_692),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1187),
.B(n_797),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1128),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1106),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1202),
.A2(n_959),
.B1(n_960),
.B2(n_898),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1156),
.B(n_1161),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1106),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1136),
.B(n_1130),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1139),
.A2(n_898),
.B(n_779),
.C(n_972),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1204),
.A2(n_804),
.B1(n_1004),
.B2(n_692),
.Y(n_1339)
);

INVxp33_ASAP7_75t_L g1340 ( 
.A(n_1156),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1191),
.B(n_1212),
.Y(n_1343)
);

BUFx5_ASAP7_75t_L g1344 ( 
.A(n_1187),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1103),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1144),
.B(n_898),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1136),
.B(n_1130),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1136),
.B(n_1130),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1227),
.Y(n_1349)
);

NAND2x1p5_ASAP7_75t_L g1350 ( 
.A(n_1187),
.B(n_797),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1149),
.A2(n_1196),
.B(n_1192),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1159),
.A2(n_898),
.B(n_833),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1136),
.B(n_1130),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1204),
.B(n_833),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1310),
.A2(n_1314),
.B1(n_1334),
.B2(n_1237),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1335),
.B(n_1340),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1286),
.B(n_1301),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1340),
.B(n_1237),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1279),
.A2(n_1276),
.B(n_1274),
.Y(n_1359)
);

AOI21x1_ASAP7_75t_SL g1360 ( 
.A1(n_1303),
.A2(n_1272),
.B(n_1254),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1285),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1266),
.B(n_1283),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1266),
.B(n_1283),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1276),
.A2(n_1255),
.B(n_1263),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1310),
.A2(n_1314),
.B1(n_1334),
.B2(n_1338),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1261),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1338),
.A2(n_1250),
.B(n_1319),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1346),
.A2(n_1329),
.B(n_1339),
.C(n_1352),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1330),
.A2(n_1253),
.B1(n_1353),
.B2(n_1348),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1286),
.B(n_1256),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1250),
.A2(n_1251),
.B(n_1346),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1280),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1317),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1246),
.B(n_1337),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1258),
.A2(n_1247),
.B(n_1307),
.C(n_1354),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1292),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1271),
.A2(n_1259),
.B(n_1265),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1267),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1293),
.B(n_1315),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1315),
.B(n_1354),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1284),
.A2(n_1295),
.B(n_1347),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1247),
.A2(n_1307),
.B(n_1275),
.C(n_1284),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1296),
.A2(n_1300),
.B(n_1270),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1238),
.A2(n_1351),
.B(n_1342),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1253),
.B(n_1275),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1290),
.B(n_1260),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1269),
.B(n_1349),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1242),
.B(n_1297),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1316),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_1288),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1288),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1306),
.B(n_1327),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1323),
.B(n_1343),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1317),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1249),
.A2(n_1278),
.B(n_1243),
.Y(n_1395)
);

AOI21x1_ASAP7_75t_SL g1396 ( 
.A1(n_1244),
.A2(n_1289),
.B(n_1264),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1278),
.B(n_1322),
.Y(n_1397)
);

AOI21x1_ASAP7_75t_SL g1398 ( 
.A1(n_1244),
.A2(n_1264),
.B(n_1257),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1327),
.A2(n_1252),
.B(n_1294),
.C(n_1345),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1235),
.B(n_1240),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1322),
.B(n_1268),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1322),
.B(n_1268),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1322),
.B(n_1268),
.Y(n_1403)
);

AOI21x1_ASAP7_75t_SL g1404 ( 
.A1(n_1308),
.A2(n_1291),
.B(n_1248),
.Y(n_1404)
);

AOI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1248),
.A2(n_1321),
.B(n_1298),
.Y(n_1405)
);

AND2x2_ASAP7_75t_SL g1406 ( 
.A(n_1313),
.B(n_1325),
.Y(n_1406)
);

OA22x2_ASAP7_75t_L g1407 ( 
.A1(n_1245),
.A2(n_1336),
.B1(n_1281),
.B2(n_1333),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1318),
.B(n_1302),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1287),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1322),
.B(n_1268),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1277),
.B(n_1282),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1318),
.B(n_1282),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1331),
.A2(n_1350),
.B1(n_1248),
.B2(n_1321),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1331),
.A2(n_1299),
.B(n_1332),
.Y(n_1414)
);

A2O1A1Ixp33_ASAP7_75t_SL g1415 ( 
.A1(n_1298),
.A2(n_1262),
.B(n_1344),
.C(n_1305),
.Y(n_1415)
);

AOI221x1_ASAP7_75t_SL g1416 ( 
.A1(n_1262),
.A2(n_1287),
.B1(n_1305),
.B2(n_1344),
.C(n_1304),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1273),
.B(n_1344),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1344),
.A2(n_1273),
.B(n_1324),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1344),
.B(n_1326),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1311),
.B(n_1312),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1320),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1328),
.B(n_1341),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1241),
.B(n_1335),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1239),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1242),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1266),
.B(n_1283),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1250),
.A2(n_1104),
.B(n_1197),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1330),
.B(n_898),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1309),
.B(n_1285),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1279),
.A2(n_1276),
.B(n_1274),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1335),
.B(n_1340),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1266),
.B(n_1283),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1285),
.Y(n_1433)
);

AOI21x1_ASAP7_75t_SL g1434 ( 
.A1(n_1303),
.A2(n_847),
.B(n_898),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1286),
.B(n_1301),
.Y(n_1435)
);

AOI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1310),
.A2(n_1314),
.B1(n_1334),
.B2(n_1237),
.C(n_1247),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1338),
.A2(n_1204),
.B(n_1144),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1338),
.A2(n_1204),
.B(n_1144),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1335),
.B(n_1340),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1279),
.A2(n_1276),
.B(n_1274),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1310),
.A2(n_1314),
.B1(n_1334),
.B2(n_1004),
.Y(n_1441)
);

OAI22x1_ASAP7_75t_L g1442 ( 
.A1(n_1270),
.A2(n_1346),
.B1(n_1300),
.B2(n_1236),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1239),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1401),
.B(n_1402),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1392),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1395),
.A2(n_1371),
.B(n_1427),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1359),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_SL g1448 ( 
.A1(n_1428),
.A2(n_1382),
.B(n_1368),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1443),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1420),
.B(n_1419),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1430),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1440),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1403),
.B(n_1410),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1420),
.B(n_1421),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1392),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1369),
.B(n_1362),
.Y(n_1456)
);

INVx4_ASAP7_75t_L g1457 ( 
.A(n_1392),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1440),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1423),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1366),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_SL g1461 ( 
.A(n_1416),
.Y(n_1461)
);

INVx4_ASAP7_75t_L g1462 ( 
.A(n_1407),
.Y(n_1462)
);

AO21x1_ASAP7_75t_SL g1463 ( 
.A1(n_1397),
.A2(n_1385),
.B(n_1419),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1407),
.Y(n_1464)
);

BUFx12f_ASAP7_75t_L g1465 ( 
.A(n_1373),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1364),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1376),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1364),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1422),
.B(n_1377),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1413),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1394),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1384),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1389),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1406),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1365),
.B(n_1355),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1413),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1369),
.B(n_1362),
.Y(n_1477)
);

CKINVDCx11_ASAP7_75t_R g1478 ( 
.A(n_1409),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1424),
.B(n_1367),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1355),
.A2(n_1365),
.B1(n_1441),
.B2(n_1436),
.Y(n_1480)
);

XNOR2xp5_ASAP7_75t_L g1481 ( 
.A(n_1441),
.B(n_1436),
.Y(n_1481)
);

OR2x6_ASAP7_75t_L g1482 ( 
.A(n_1381),
.B(n_1437),
.Y(n_1482)
);

AO21x2_ASAP7_75t_L g1483 ( 
.A1(n_1415),
.A2(n_1385),
.B(n_1426),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1405),
.A2(n_1404),
.B(n_1418),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1361),
.B(n_1433),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1363),
.A2(n_1426),
.B(n_1432),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1358),
.B(n_1356),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1363),
.A2(n_1432),
.B(n_1438),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1391),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1431),
.B(n_1439),
.Y(n_1490)
);

OA21x2_ASAP7_75t_L g1491 ( 
.A1(n_1374),
.A2(n_1400),
.B(n_1372),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1383),
.B(n_1399),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1375),
.B(n_1417),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1442),
.A2(n_1380),
.B1(n_1429),
.B2(n_1390),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1386),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1449),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1463),
.B(n_1379),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1445),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1470),
.B(n_1387),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1463),
.B(n_1435),
.Y(n_1500)
);

AO21x2_ASAP7_75t_L g1501 ( 
.A1(n_1446),
.A2(n_1411),
.B(n_1414),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1470),
.B(n_1378),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1449),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1491),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_L g1505 ( 
.A(n_1482),
.B(n_1425),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1444),
.B(n_1357),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1486),
.B(n_1435),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1482),
.A2(n_1370),
.B(n_1393),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1491),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1454),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1450),
.Y(n_1511)
);

INVxp67_ASAP7_75t_SL g1512 ( 
.A(n_1469),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1486),
.B(n_1388),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1450),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1491),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1484),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1476),
.B(n_1469),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1453),
.B(n_1388),
.Y(n_1518)
);

OAI211xp5_ASAP7_75t_L g1519 ( 
.A1(n_1448),
.A2(n_1396),
.B(n_1360),
.C(n_1434),
.Y(n_1519)
);

AO21x2_ASAP7_75t_L g1520 ( 
.A1(n_1446),
.A2(n_1451),
.B(n_1458),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1507),
.A2(n_1480),
.B1(n_1475),
.B2(n_1481),
.C(n_1456),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1511),
.B(n_1514),
.Y(n_1522)
);

AOI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1507),
.A2(n_1480),
.B1(n_1475),
.B2(n_1481),
.C(n_1456),
.Y(n_1523)
);

AOI33xp33_ASAP7_75t_L g1524 ( 
.A1(n_1497),
.A2(n_1494),
.A3(n_1479),
.B1(n_1487),
.B2(n_1495),
.B3(n_1453),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1505),
.B(n_1492),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1520),
.A2(n_1451),
.B(n_1447),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1496),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1498),
.Y(n_1528)
);

AOI31xp33_ASAP7_75t_L g1529 ( 
.A1(n_1505),
.A2(n_1481),
.A3(n_1492),
.B(n_1494),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1519),
.A2(n_1482),
.B(n_1477),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1496),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1499),
.B(n_1486),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1497),
.A2(n_1482),
.B1(n_1477),
.B2(n_1488),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1499),
.B(n_1486),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1496),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1497),
.A2(n_1482),
.B1(n_1488),
.B2(n_1486),
.Y(n_1536)
);

AOI211xp5_ASAP7_75t_L g1537 ( 
.A1(n_1519),
.A2(n_1479),
.B(n_1461),
.C(n_1474),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1499),
.Y(n_1538)
);

AO21x2_ASAP7_75t_L g1539 ( 
.A1(n_1520),
.A2(n_1458),
.B(n_1452),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1503),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1497),
.A2(n_1461),
.B1(n_1482),
.B2(n_1488),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1498),
.Y(n_1542)
);

AND4x1_ASAP7_75t_L g1543 ( 
.A(n_1505),
.B(n_1479),
.C(n_1398),
.D(n_1465),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1506),
.B(n_1465),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1502),
.A2(n_1474),
.B1(n_1465),
.B2(n_1462),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1500),
.A2(n_1488),
.B1(n_1474),
.B2(n_1455),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1500),
.A2(n_1488),
.B1(n_1474),
.B2(n_1493),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1508),
.A2(n_1493),
.B(n_1484),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1506),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1500),
.A2(n_1493),
.B1(n_1455),
.B2(n_1445),
.Y(n_1550)
);

OA21x2_ASAP7_75t_L g1551 ( 
.A1(n_1504),
.A2(n_1468),
.B(n_1466),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1511),
.B(n_1450),
.Y(n_1552)
);

AOI222xp33_ASAP7_75t_L g1553 ( 
.A1(n_1512),
.A2(n_1478),
.B1(n_1489),
.B2(n_1465),
.C1(n_1464),
.C2(n_1490),
.Y(n_1553)
);

OAI33xp33_ASAP7_75t_L g1554 ( 
.A1(n_1517),
.A2(n_1489),
.A3(n_1485),
.B1(n_1460),
.B2(n_1473),
.B3(n_1467),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1511),
.B(n_1459),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1503),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1511),
.B(n_1459),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1508),
.A2(n_1493),
.B(n_1484),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1548),
.A2(n_1472),
.B(n_1468),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1527),
.Y(n_1560)
);

NOR3xp33_ASAP7_75t_L g1561 ( 
.A(n_1529),
.B(n_1478),
.C(n_1513),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1551),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1538),
.B(n_1512),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1532),
.B(n_1517),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1525),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1527),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1531),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1551),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1551),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1551),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1526),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1526),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1548),
.A2(n_1472),
.B(n_1466),
.Y(n_1573)
);

INVx5_ASAP7_75t_L g1574 ( 
.A(n_1522),
.Y(n_1574)
);

INVx4_ASAP7_75t_L g1575 ( 
.A(n_1528),
.Y(n_1575)
);

AND2x6_ASAP7_75t_SL g1576 ( 
.A(n_1544),
.B(n_1408),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1552),
.B(n_1514),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1531),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1535),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1552),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1526),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1535),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1526),
.Y(n_1583)
);

INVx3_ASAP7_75t_SL g1584 ( 
.A(n_1528),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1540),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1528),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1552),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1558),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1552),
.B(n_1514),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1534),
.B(n_1517),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1540),
.B(n_1483),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_L g1592 ( 
.A(n_1521),
.B(n_1516),
.C(n_1509),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1556),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1539),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1565),
.B(n_1523),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1575),
.B(n_1558),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1560),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1560),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1566),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1566),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1567),
.Y(n_1603)
);

AOI33xp33_ASAP7_75t_L g1604 ( 
.A1(n_1592),
.A2(n_1546),
.A3(n_1536),
.B1(n_1541),
.B2(n_1533),
.B3(n_1537),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1567),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1578),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1574),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1575),
.B(n_1542),
.Y(n_1608)
);

O2A1O1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1592),
.A2(n_1529),
.B(n_1537),
.C(n_1530),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1565),
.B(n_1524),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1588),
.B(n_1557),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1584),
.B(n_1557),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1578),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1584),
.B(n_1542),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1584),
.B(n_1542),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1579),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1579),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1584),
.B(n_1549),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1564),
.B(n_1513),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1582),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1586),
.B(n_1541),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1586),
.B(n_1510),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1586),
.B(n_1510),
.Y(n_1623)
);

NAND3xp33_ASAP7_75t_SL g1624 ( 
.A(n_1561),
.B(n_1553),
.C(n_1543),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1561),
.B(n_1506),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1586),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1582),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1575),
.B(n_1510),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_L g1629 ( 
.A(n_1591),
.B(n_1553),
.C(n_1547),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1585),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1585),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1568),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1590),
.B(n_1518),
.Y(n_1633)
);

AOI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1590),
.A2(n_1554),
.B1(n_1509),
.B2(n_1504),
.C(n_1515),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1576),
.B(n_1471),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1575),
.B(n_1501),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1564),
.B(n_1563),
.Y(n_1637)
);

NOR3x1_ASAP7_75t_L g1638 ( 
.A(n_1624),
.B(n_1595),
.C(n_1610),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1609),
.B(n_1575),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1604),
.B(n_1563),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1598),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1598),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1637),
.B(n_1564),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1599),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1626),
.B(n_1621),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1599),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1637),
.B(n_1502),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1614),
.B(n_1615),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1605),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1632),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1607),
.B(n_1574),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1633),
.B(n_1591),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1605),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1606),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1606),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1613),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1613),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1625),
.B(n_1502),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1616),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1616),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1617),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1617),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1627),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1619),
.B(n_1593),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1621),
.B(n_1490),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1618),
.A2(n_1559),
.B(n_1573),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1596),
.B(n_1490),
.Y(n_1668)
);

AND2x4_ASAP7_75t_SL g1669 ( 
.A(n_1608),
.B(n_1580),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1627),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1615),
.B(n_1580),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1635),
.A2(n_1573),
.B(n_1559),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1630),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1653),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1651),
.B(n_1607),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1648),
.B(n_1608),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1648),
.B(n_1608),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1645),
.B(n_1596),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1669),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1669),
.B(n_1612),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1639),
.A2(n_1629),
.B(n_1634),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1656),
.B(n_1612),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1656),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1653),
.Y(n_1685)
);

OAI31xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1639),
.A2(n_1597),
.A3(n_1601),
.B(n_1611),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1671),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1641),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1666),
.B(n_1600),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1642),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1671),
.A2(n_1597),
.B1(n_1611),
.B2(n_1601),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1668),
.B(n_1622),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1644),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1659),
.A2(n_1597),
.B1(n_1545),
.B2(n_1457),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1643),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1646),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1654),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1672),
.A2(n_1607),
.B(n_1636),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1685),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1682),
.A2(n_1667),
.B1(n_1545),
.B2(n_1559),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1679),
.B(n_1647),
.Y(n_1703)
);

NOR4xp25_ASAP7_75t_L g1704 ( 
.A(n_1678),
.B(n_1670),
.C(n_1655),
.D(n_1664),
.Y(n_1704)
);

OAI21xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1686),
.A2(n_1658),
.B(n_1657),
.Y(n_1705)
);

AOI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1685),
.A2(n_1573),
.B(n_1636),
.C(n_1663),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1687),
.B(n_1660),
.Y(n_1707)
);

NAND4xp25_ASAP7_75t_L g1708 ( 
.A(n_1695),
.B(n_1662),
.C(n_1661),
.D(n_1550),
.Y(n_1708)
);

OAI31xp33_ASAP7_75t_L g1709 ( 
.A1(n_1685),
.A2(n_1623),
.A3(n_1628),
.B(n_1665),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1691),
.A2(n_1680),
.B1(n_1684),
.B2(n_1694),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1699),
.A2(n_1628),
.B(n_1650),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1680),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1674),
.Y(n_1713)
);

OAI21xp33_ASAP7_75t_L g1714 ( 
.A1(n_1676),
.A2(n_1652),
.B(n_1665),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1680),
.A2(n_1574),
.B1(n_1587),
.B2(n_1623),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1674),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1676),
.B(n_1577),
.Y(n_1717)
);

NAND2x1p5_ASAP7_75t_L g1718 ( 
.A(n_1681),
.B(n_1543),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1693),
.A2(n_1650),
.B1(n_1652),
.B2(n_1602),
.C(n_1620),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1700),
.B(n_1674),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1712),
.B(n_1677),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1713),
.B(n_1677),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1718),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1710),
.B(n_1683),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_SL g1726 ( 
.A(n_1709),
.B(n_1681),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1705),
.B(n_1708),
.Y(n_1727)
);

OAI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1701),
.A2(n_1697),
.B1(n_1693),
.B2(n_1692),
.C(n_1689),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1716),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1709),
.B(n_1714),
.Y(n_1730)
);

O2A1O1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1723),
.A2(n_1702),
.B(n_1707),
.C(n_1711),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1727),
.A2(n_1719),
.B1(n_1706),
.B2(n_1698),
.C(n_1690),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1730),
.A2(n_1706),
.B(n_1715),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1725),
.A2(n_1703),
.B(n_1675),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1726),
.A2(n_1698),
.B(n_1696),
.C(n_1690),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1728),
.A2(n_1696),
.B1(n_1688),
.B2(n_1675),
.C(n_1717),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1721),
.B(n_1688),
.Y(n_1737)
);

NOR3x1_ASAP7_75t_L g1738 ( 
.A(n_1729),
.B(n_1689),
.C(n_1587),
.Y(n_1738)
);

AOI322xp5_ASAP7_75t_L g1739 ( 
.A1(n_1720),
.A2(n_1724),
.A3(n_1722),
.B1(n_1568),
.B2(n_1675),
.C1(n_1572),
.C2(n_1571),
.Y(n_1739)
);

OAI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1722),
.A2(n_1574),
.B(n_1583),
.C(n_1572),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1727),
.A2(n_1675),
.B1(n_1571),
.B2(n_1583),
.C(n_1572),
.Y(n_1741)
);

O2A1O1Ixp5_ASAP7_75t_SL g1742 ( 
.A1(n_1740),
.A2(n_1631),
.B(n_1630),
.C(n_1603),
.Y(n_1742)
);

AOI221x1_ASAP7_75t_L g1743 ( 
.A1(n_1733),
.A2(n_1631),
.B1(n_1632),
.B2(n_1572),
.C(n_1571),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1731),
.A2(n_1571),
.B1(n_1583),
.B2(n_1594),
.C(n_1581),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_R g1745 ( 
.A(n_1737),
.B(n_1576),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1732),
.A2(n_1583),
.B(n_1568),
.C(n_1587),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1735),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1747),
.B(n_1734),
.Y(n_1748)
);

NAND3xp33_ASAP7_75t_L g1749 ( 
.A(n_1746),
.B(n_1743),
.C(n_1736),
.Y(n_1749)
);

INVxp67_ASAP7_75t_L g1750 ( 
.A(n_1744),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1742),
.B(n_1739),
.C(n_1741),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1745),
.B(n_1738),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1747),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1752),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1753),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1749),
.A2(n_1574),
.B1(n_1619),
.B2(n_1589),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1748),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1750),
.B(n_1574),
.Y(n_1758)
);

NAND4xp25_ASAP7_75t_L g1759 ( 
.A(n_1756),
.B(n_1758),
.C(n_1757),
.D(n_1755),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1754),
.Y(n_1760)
);

NOR2xp67_ASAP7_75t_R g1761 ( 
.A(n_1755),
.B(n_1751),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1760),
.B(n_1568),
.Y(n_1762)
);

NOR2x1_ASAP7_75t_L g1763 ( 
.A(n_1762),
.B(n_1759),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1763),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1763),
.Y(n_1765)
);

AOI22x1_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1761),
.B1(n_1594),
.B2(n_1581),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1765),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1767),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1766),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1768),
.A2(n_1764),
.B1(n_1765),
.B2(n_1574),
.Y(n_1770)
);

AOI222xp33_ASAP7_75t_SL g1771 ( 
.A1(n_1769),
.A2(n_1581),
.B1(n_1594),
.B2(n_1568),
.C1(n_1569),
.C2(n_1562),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1770),
.B(n_1574),
.Y(n_1772)
);

AOI222xp33_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1771),
.B1(n_1562),
.B2(n_1569),
.C1(n_1570),
.C2(n_1593),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1569),
.B1(n_1562),
.B2(n_1570),
.Y(n_1774)
);

AOI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1569),
.B1(n_1562),
.B2(n_1570),
.Y(n_1775)
);

AOI211xp5_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1412),
.B(n_1485),
.C(n_1516),
.Y(n_1776)
);


endmodule