module fake_jpeg_29973_n_158 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_20),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_39),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_49),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_46),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_89),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_85),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_49),
.B1(n_58),
.B2(n_56),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_74),
.B1(n_68),
.B2(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_61),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_58),
.B1(n_65),
.B2(n_53),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_52),
.B1(n_60),
.B2(n_63),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_66),
.B(n_51),
.C(n_5),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_98),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_87),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_97),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_68),
.B1(n_69),
.B2(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_100),
.B1(n_103),
.B2(n_2),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_47),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_59),
.B1(n_57),
.B2(n_55),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_48),
.B1(n_54),
.B2(n_5),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_54),
.C(n_22),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_54),
.C(n_23),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_29),
.B(n_45),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_110),
.Y(n_115)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_21),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_120),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_116),
.B1(n_117),
.B2(n_30),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_7),
.B(n_9),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_9),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_10),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_18),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_17),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_11),
.B(n_14),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_137),
.B1(n_138),
.B2(n_143),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_15),
.B(n_16),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_115),
.B(n_112),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_142),
.C(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_19),
.B(n_27),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_149),
.Y(n_152)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_119),
.B(n_133),
.Y(n_150)
);

OA21x2_ASAP7_75t_SL g153 ( 
.A1(n_150),
.A2(n_151),
.B(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_132),
.Y(n_154)
);

OAI31xp33_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_136),
.A3(n_152),
.B(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_148),
.B1(n_146),
.B2(n_144),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_135),
.B1(n_148),
.B2(n_127),
.Y(n_157)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_135),
.B1(n_124),
.B2(n_42),
.C(n_43),
.Y(n_158)
);


endmodule