module fake_jpeg_3865_n_39 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_39);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_16),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_4),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_2),
.A2(n_9),
.B(n_4),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_15),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_21),
.A3(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_31),
.B(n_27),
.Y(n_34)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_5),
.B1(n_10),
.B2(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_35),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_31),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_0),
.C2(n_17),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_39)
);


endmodule