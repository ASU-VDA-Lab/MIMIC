module fake_jpeg_629_n_84 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_84);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_84;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_0),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_31),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_28),
.Y(n_40)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_29),
.C(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_41),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_27),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_35),
.B1(n_40),
.B2(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_46),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_57),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_33),
.B(n_42),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_1),
.B(n_2),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_2),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_1),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_34),
.B1(n_24),
.B2(n_23),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_34),
.B1(n_11),
.B2(n_14),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_62),
.B1(n_15),
.B2(n_19),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_53),
.C(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_72),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_4),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_60),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_70),
.B(n_8),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_78),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_79),
.A2(n_75),
.B(n_73),
.Y(n_80)
);

AOI322xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_76),
.A3(n_17),
.B1(n_16),
.B2(n_18),
.C1(n_20),
.C2(n_10),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_6),
.B(n_9),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_10),
.Y(n_84)
);


endmodule