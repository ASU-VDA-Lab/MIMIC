module fake_jpeg_73_n_233 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_7),
.B(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_52),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_57),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_54),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_20),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_59),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_32),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_63),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_37),
.Y(n_67)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_67),
.B(n_76),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_81),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_37),
.B1(n_23),
.B2(n_33),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_82),
.B1(n_62),
.B2(n_58),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_20),
.B1(n_26),
.B2(n_29),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_73),
.A2(n_74),
.B1(n_77),
.B2(n_83),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_34),
.B1(n_36),
.B2(n_31),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_34),
.B1(n_31),
.B2(n_36),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_33),
.B1(n_25),
.B2(n_32),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_18),
.B1(n_24),
.B2(n_17),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_18),
.B1(n_30),
.B2(n_24),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_18),
.B1(n_27),
.B2(n_3),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_86),
.B1(n_99),
.B2(n_82),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_18),
.B1(n_27),
.B2(n_4),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_27),
.B1(n_1),
.B2(n_5),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_42),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_70),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_51),
.A2(n_27),
.B1(n_6),
.B2(n_8),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_27),
.B1(n_6),
.B2(n_8),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_109),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_63),
.B1(n_40),
.B2(n_45),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_110),
.B1(n_125),
.B2(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_1),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_116),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_45),
.C(n_9),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_81),
.C(n_96),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_1),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_112),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_11),
.B1(n_14),
.B2(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_68),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_78),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_80),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_90),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_129),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_66),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_130),
.A2(n_110),
.B(n_109),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_102),
.B1(n_101),
.B2(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_104),
.B1(n_103),
.B2(n_117),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_154),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_106),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_79),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_142),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_66),
.B(n_79),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_113),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_95),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_96),
.B(n_90),
.C(n_93),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_152),
.B(n_129),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_101),
.A2(n_95),
.B1(n_75),
.B2(n_93),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_118),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_93),
.B(n_75),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_93),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_136),
.C(n_142),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_111),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_162),
.Y(n_180)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_171),
.C(n_153),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_108),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_167),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_164),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_145),
.B(n_137),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_172),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_127),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_144),
.B(n_152),
.Y(n_181)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_119),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_133),
.B(n_143),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_126),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_75),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_148),
.B1(n_132),
.B2(n_154),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_178),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_161),
.A2(n_150),
.B1(n_145),
.B2(n_137),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_192),
.C(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_191),
.C(n_159),
.Y(n_194)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_139),
.C(n_138),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_171),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_194),
.C(n_197),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_161),
.A3(n_172),
.B1(n_173),
.B2(n_150),
.C1(n_165),
.C2(n_170),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_179),
.A3(n_180),
.B1(n_192),
.B2(n_187),
.C1(n_183),
.C2(n_191),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_165),
.C(n_170),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_174),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_169),
.C(n_155),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_176),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_188),
.C(n_185),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_181),
.B(n_180),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_210),
.A2(n_196),
.B(n_205),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_180),
.B1(n_130),
.B2(n_150),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_214),
.B(n_194),
.CI(n_197),
.CON(n_215),
.SN(n_215)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_214),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_218),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_209),
.C(n_211),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_210),
.B(n_206),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_221),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_223),
.C(n_185),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_206),
.C(n_213),
.Y(n_223)
);

AOI21x1_ASAP7_75t_SL g226 ( 
.A1(n_224),
.A2(n_216),
.B(n_218),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_220),
.B(n_225),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_162),
.B(n_143),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_230),
.B(n_231),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_156),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_228),
.Y(n_233)
);


endmodule