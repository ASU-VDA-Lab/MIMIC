module fake_netlist_1_316_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_6), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
NOR2xp33_ASAP7_75t_R g20 ( .A(n_16), .B(n_3), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_15), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_15), .Y(n_23) );
BUFx2_ASAP7_75t_L g24 ( .A(n_12), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
AND2x4_ASAP7_75t_L g26 ( .A(n_21), .B(n_11), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_14), .B1(n_17), .B2(n_13), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_19), .Y(n_28) );
NOR4xp25_ASAP7_75t_SL g29 ( .A(n_25), .B(n_23), .C(n_20), .D(n_0), .Y(n_29) );
BUFx2_ASAP7_75t_L g30 ( .A(n_26), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx1_ASAP7_75t_SL g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AOI221x1_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_27), .B1(n_13), .B2(n_22), .C(n_26), .Y(n_34) );
NOR3xp33_ASAP7_75t_SL g35 ( .A(n_32), .B(n_29), .C(n_30), .Y(n_35) );
NAND4xp25_ASAP7_75t_L g36 ( .A(n_34), .B(n_2), .C(n_13), .D(n_20), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
NOR2xp33_ASAP7_75t_L g38 ( .A(n_34), .B(n_13), .Y(n_38) );
INVx1_ASAP7_75t_SL g39 ( .A(n_37), .Y(n_39) );
NOR3xp33_ASAP7_75t_L g40 ( .A(n_36), .B(n_5), .C(n_7), .Y(n_40) );
INVx3_ASAP7_75t_L g41 ( .A(n_39), .Y(n_41) );
AOI22xp5_ASAP7_75t_L g42 ( .A1(n_41), .A2(n_40), .B1(n_38), .B2(n_9), .Y(n_42) );
endmodule