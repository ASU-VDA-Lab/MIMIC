module fake_jpeg_2869_n_421 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_421);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx3_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_55),
.B(n_57),
.Y(n_136)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g115 ( 
.A(n_56),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_15),
.A2(n_28),
.B(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_61),
.B(n_77),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_88),
.Y(n_130)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_20),
.B(n_14),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_92),
.Y(n_118)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_90),
.B(n_91),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_44),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_0),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_31),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_95),
.Y(n_121)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_22),
.B1(n_37),
.B2(n_28),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_98),
.Y(n_140)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_50),
.A2(n_38),
.B1(n_46),
.B2(n_22),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_101),
.A2(n_103),
.B1(n_111),
.B2(n_129),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_46),
.B1(n_38),
.B2(n_24),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_110),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_37),
.B1(n_22),
.B2(n_26),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_24),
.B1(n_25),
.B2(n_21),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_59),
.A2(n_21),
.B1(n_25),
.B2(n_39),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_85),
.A2(n_90),
.B1(n_37),
.B2(n_63),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_137),
.B1(n_138),
.B2(n_76),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_74),
.A2(n_16),
.B1(n_41),
.B2(n_39),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_58),
.A2(n_47),
.B1(n_41),
.B2(n_33),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_73),
.A2(n_47),
.B1(n_33),
.B2(n_30),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_72),
.B1(n_68),
.B2(n_56),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_75),
.B(n_30),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_51),
.B(n_16),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_147),
.B(n_69),
.Y(n_163)
);

HAxp5_ASAP7_75t_SL g153 ( 
.A(n_69),
.B(n_4),
.CON(n_153),
.SN(n_153)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_93),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_158),
.Y(n_209)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_86),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_78),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_165),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_78),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_115),
.Y(n_166)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_178),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_122),
.A2(n_97),
.B1(n_62),
.B2(n_64),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_137),
.B1(n_110),
.B2(n_138),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_176),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_96),
.B1(n_76),
.B2(n_60),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_175),
.B1(n_126),
.B2(n_106),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_84),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_126),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_79),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_125),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_104),
.B(n_66),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_183),
.B(n_186),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_193),
.B1(n_102),
.B2(n_150),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_130),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_4),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_65),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_195),
.Y(n_215)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_123),
.B(n_5),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_123),
.B(n_5),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_5),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_101),
.A2(n_82),
.B1(n_80),
.B2(n_65),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_152),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_102),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_221),
.B1(n_195),
.B2(n_183),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_143),
.A3(n_132),
.B1(n_153),
.B2(n_111),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_199),
.A2(n_220),
.B(n_167),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_201),
.A2(n_109),
.B1(n_194),
.B2(n_180),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_108),
.B(n_117),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_166),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_214),
.B(n_217),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_162),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_124),
.B(n_113),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_174),
.A2(n_119),
.B1(n_131),
.B2(n_152),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_162),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_174),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_133),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_230),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_164),
.B1(n_189),
.B2(n_192),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_236),
.B1(n_242),
.B2(n_251),
.Y(n_261)
);

BUFx8_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_238),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_216),
.A2(n_178),
.B1(n_185),
.B2(n_184),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_170),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_237),
.B(n_256),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_158),
.C(n_161),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_229),
.Y(n_262)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_186),
.B1(n_159),
.B2(n_154),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_250),
.B1(n_255),
.B2(n_196),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_131),
.B1(n_119),
.B2(n_150),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_201),
.A2(n_181),
.B1(n_195),
.B2(n_168),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_217),
.B1(n_222),
.B2(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_99),
.B1(n_116),
.B2(n_179),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_221),
.A2(n_116),
.B1(n_99),
.B2(n_156),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_157),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_200),
.Y(n_280)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_197),
.B(n_188),
.C(n_169),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_215),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_229),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_234),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_264),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_218),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_197),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_274),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_218),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_268),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_SL g274 ( 
.A(n_233),
.B(n_215),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_211),
.B1(n_206),
.B2(n_212),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_278),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_235),
.A2(n_220),
.B(n_199),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_286),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_208),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_198),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_283),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_234),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_234),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_248),
.Y(n_293)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_288),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_241),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_289),
.B(n_303),
.Y(n_316)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_300),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_293),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_198),
.Y(n_322)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_296),
.Y(n_321)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_297),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_254),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_308),
.Y(n_323)
);

AO21x2_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_243),
.B(n_238),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_255),
.Y(n_331)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_231),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_306),
.B(n_310),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_248),
.B1(n_236),
.B2(n_246),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_273),
.B1(n_276),
.B2(n_268),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_274),
.B(n_260),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_287),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_260),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_279),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_312),
.A2(n_326),
.B1(n_333),
.B2(n_331),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_278),
.C(n_267),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_317),
.C(n_325),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_273),
.C(n_272),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_309),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_319),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_301),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_272),
.C(n_270),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_305),
.A2(n_284),
.B1(n_270),
.B2(n_266),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_298),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_327),
.A2(n_334),
.B1(n_228),
.B2(n_224),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_295),
.C(n_311),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_308),
.C(n_307),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_261),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_330),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_R g349 ( 
.A(n_331),
.B(n_258),
.C(n_252),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_279),
.Y(n_332)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_332),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_292),
.A2(n_242),
.B1(n_282),
.B2(n_257),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_300),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_340),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_297),
.C(n_282),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_343),
.C(n_350),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_313),
.A2(n_304),
.B(n_301),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_339),
.A2(n_321),
.B(n_320),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_292),
.B1(n_304),
.B2(n_305),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_341),
.A2(n_344),
.B1(n_352),
.B2(n_353),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_301),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_347),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_231),
.C(n_225),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_324),
.A2(n_290),
.B1(n_230),
.B2(n_244),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_345),
.A2(n_202),
.B1(n_219),
.B2(n_203),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_240),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_318),
.A2(n_333),
.B1(n_312),
.B2(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_348),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_322),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_225),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_315),
.A2(n_251),
.B1(n_228),
.B2(n_200),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_205),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_205),
.C(n_190),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_340),
.A2(n_315),
.B(n_329),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_357),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_342),
.A2(n_332),
.B(n_330),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_359),
.Y(n_382)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_346),
.B(n_203),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_366),
.Y(n_371)
);

OAI321xp33_ASAP7_75t_L g362 ( 
.A1(n_351),
.A2(n_200),
.A3(n_249),
.B1(n_202),
.B2(n_219),
.C(n_10),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_362),
.A2(n_369),
.B(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_365),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_249),
.C(n_42),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_335),
.C(n_336),
.Y(n_372)
);

XNOR2x1_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_249),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_349),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_6),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_368),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_338),
.C(n_364),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_373),
.B(n_377),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_374),
.A2(n_367),
.B1(n_366),
.B2(n_365),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_354),
.C(n_337),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_379),
.A2(n_12),
.B1(n_13),
.B2(n_36),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_357),
.A2(n_347),
.B(n_337),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_380),
.A2(n_36),
.B(n_42),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_6),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_381),
.B(n_8),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_360),
.A2(n_352),
.B(n_9),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_383),
.A2(n_8),
.B(n_12),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_382),
.A2(n_356),
.B1(n_355),
.B2(n_368),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_386),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_372),
.C(n_376),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_382),
.A2(n_364),
.B1(n_370),
.B2(n_359),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_388),
.Y(n_401)
);

FAx1_ASAP7_75t_SL g389 ( 
.A(n_375),
.B(n_369),
.CI(n_9),
.CON(n_389),
.SN(n_389)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_390),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_378),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_376),
.A2(n_12),
.B(n_13),
.Y(n_392)
);

AOI21xp33_ASAP7_75t_SL g395 ( 
.A1(n_392),
.A2(n_393),
.B(n_371),
.Y(n_395)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_395),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_394),
.B(n_373),
.C(n_377),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_400),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_399),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_383),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_13),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_390),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_386),
.Y(n_407)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_407),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_396),
.A2(n_392),
.B(n_389),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_408),
.A2(n_402),
.B(n_407),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_409),
.B(n_410),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_389),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_405),
.B(n_399),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_412),
.B(n_42),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_413),
.A2(n_406),
.B(n_404),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g418 ( 
.A(n_415),
.Y(n_418)
);

O2A1O1Ixp33_ASAP7_75t_SL g416 ( 
.A1(n_414),
.A2(n_13),
.B(n_42),
.C(n_411),
.Y(n_416)
);

BUFx24_ASAP7_75t_SL g419 ( 
.A(n_418),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_419),
.Y(n_420)
);

AO21x1_ASAP7_75t_L g421 ( 
.A1(n_420),
.A2(n_417),
.B(n_416),
.Y(n_421)
);


endmodule