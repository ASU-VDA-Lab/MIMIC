module fake_jpeg_85_n_194 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_194);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_7),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_1),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_69),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_78),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_83),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_57),
.B1(n_51),
.B2(n_65),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_82),
.B1(n_90),
.B2(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_57),
.B1(n_61),
.B2(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_62),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_61),
.B1(n_55),
.B2(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_59),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_84),
.B(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_107),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_99),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_73),
.B1(n_81),
.B2(n_87),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_75),
.B1(n_71),
.B2(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_77),
.B1(n_56),
.B2(n_52),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_58),
.A3(n_67),
.B1(n_53),
.B2(n_60),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_58),
.Y(n_112)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_91),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_106),
.C(n_101),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_70),
.B1(n_55),
.B2(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_6),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_43),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_128),
.C(n_7),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_75),
.B1(n_71),
.B2(n_60),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_66),
.B1(n_54),
.B2(n_77),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_56),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_127),
.C(n_44),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_23),
.B(n_46),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_1),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_48),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_4),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_4),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_140),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_5),
.B(n_6),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_147),
.B(n_9),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_5),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_8),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_8),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_41),
.C(n_25),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_9),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_29),
.B1(n_13),
.B2(n_14),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_15),
.C(n_16),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_34),
.C(n_33),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_163),
.C(n_15),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_148),
.B1(n_143),
.B2(n_139),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_166),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_31),
.C(n_30),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_147),
.B1(n_13),
.B2(n_14),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_171),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_10),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_173),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_16),
.B(n_17),
.C(n_161),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_155),
.B(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_152),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_176),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_167),
.B(n_165),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_181),
.B1(n_180),
.B2(n_182),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_164),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_185),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_169),
.B1(n_162),
.B2(n_154),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_187),
.B(n_151),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_153),
.C(n_158),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_189),
.A2(n_179),
.B(n_173),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_188),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

AOI31xp33_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_187),
.A3(n_174),
.B(n_163),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_159),
.Y(n_194)
);


endmodule