module real_aes_8372_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_693;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_0), .A2(n_205), .B1(n_344), .B2(n_510), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_1), .A2(n_214), .B1(n_331), .B2(n_458), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_2), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_3), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_4), .B(n_329), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_5), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_6), .A2(n_16), .B1(n_557), .B2(n_698), .Y(n_697) );
AOI22xp5_ASAP7_75t_SL g623 ( .A1(n_7), .A2(n_50), .B1(n_288), .B2(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_8), .A2(n_19), .B1(n_262), .B2(n_431), .Y(n_603) );
INVx1_ASAP7_75t_L g675 ( .A(n_9), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_9), .A2(n_675), .B1(n_679), .B2(n_706), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_10), .B(n_329), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_11), .A2(n_64), .B1(n_555), .B2(n_557), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_12), .A2(n_108), .B1(n_293), .B2(n_296), .Y(n_292) );
XOR2x2_ASAP7_75t_L g469 ( .A(n_13), .B(n_470), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_14), .A2(n_155), .B1(n_435), .B2(n_461), .Y(n_472) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_15), .A2(n_123), .B1(n_495), .B2(n_497), .Y(n_494) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_17), .A2(n_93), .B1(n_113), .B2(n_417), .C1(n_465), .C2(n_466), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_18), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_20), .A2(n_29), .B1(n_305), .B2(n_317), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_21), .A2(n_215), .B1(n_305), .B2(n_498), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_22), .A2(n_546), .B1(n_583), .B2(n_584), .Y(n_545) );
INVx1_ASAP7_75t_L g584 ( .A(n_22), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_23), .A2(n_151), .B1(n_273), .B2(n_278), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_24), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_25), .Y(n_378) );
AO22x2_ASAP7_75t_L g246 ( .A1(n_26), .A2(n_74), .B1(n_247), .B2(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g641 ( .A(n_26), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_27), .Y(n_436) );
AOI22xp5_ASAP7_75t_SL g622 ( .A1(n_28), .A2(n_219), .B1(n_341), .B2(n_344), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_30), .A2(n_54), .B1(n_517), .B2(n_518), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_31), .B(n_327), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_32), .A2(n_138), .B1(n_274), .B2(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_33), .A2(n_70), .B1(n_268), .B2(n_512), .Y(n_562) );
AOI22xp5_ASAP7_75t_SL g618 ( .A1(n_34), .A2(n_121), .B1(n_343), .B2(n_389), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_35), .A2(n_46), .B1(n_416), .B2(n_417), .Y(n_415) );
AOI222xp33_ASAP7_75t_L g604 ( .A1(n_36), .A2(n_111), .B1(n_169), .B2(n_416), .C1(n_417), .C2(n_465), .Y(n_604) );
AO22x2_ASAP7_75t_L g251 ( .A1(n_37), .A2(n_76), .B1(n_247), .B2(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g642 ( .A(n_37), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_38), .A2(n_57), .B1(n_300), .B2(n_305), .Y(n_299) );
AOI222xp33_ASAP7_75t_L g309 ( .A1(n_39), .A2(n_137), .B1(n_179), .B2(n_310), .C1(n_312), .C2(n_316), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_40), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_41), .A2(n_139), .B1(n_431), .B2(n_452), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_42), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_43), .A2(n_71), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_44), .A2(n_116), .B1(n_704), .B2(n_705), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_45), .Y(n_420) );
XOR2xp5_ASAP7_75t_L g448 ( .A(n_47), .B(n_449), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_48), .A2(n_196), .B1(n_389), .B2(n_602), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_49), .A2(n_488), .B1(n_489), .B2(n_520), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_49), .Y(n_488) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_51), .A2(n_117), .B1(n_302), .B2(n_305), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_52), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_53), .A2(n_197), .B1(n_396), .B2(n_477), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_55), .A2(n_98), .B1(n_452), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_56), .A2(n_112), .B1(n_387), .B2(n_389), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_58), .A2(n_163), .B1(n_274), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g390 ( .A1(n_59), .A2(n_99), .B1(n_350), .B2(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_60), .A2(n_129), .B1(n_331), .B2(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g483 ( .A(n_61), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_62), .B(n_293), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_63), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_65), .A2(n_79), .B1(n_283), .B2(n_288), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_66), .A2(n_207), .B1(n_458), .B2(n_616), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_67), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_68), .A2(n_209), .B1(n_318), .B2(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_69), .A2(n_75), .B1(n_455), .B2(n_456), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_72), .A2(n_177), .B1(n_306), .B2(n_458), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_73), .A2(n_109), .B1(n_349), .B2(n_394), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_77), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_78), .B(n_503), .Y(n_614) );
INVx1_ASAP7_75t_L g229 ( .A(n_80), .Y(n_229) );
AOI22xp33_ASAP7_75t_SL g340 ( .A1(n_81), .A2(n_135), .B1(n_283), .B2(n_341), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_82), .A2(n_94), .B1(n_257), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_83), .A2(n_120), .B1(n_317), .B2(n_375), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_84), .A2(n_162), .B1(n_242), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_85), .A2(n_97), .B1(n_257), .B2(n_427), .Y(n_590) );
INVx1_ASAP7_75t_L g226 ( .A(n_86), .Y(n_226) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_87), .A2(n_95), .B1(n_349), .B2(n_350), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_88), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_89), .B(n_498), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_90), .A2(n_124), .B1(n_262), .B2(n_268), .Y(n_261) );
OA22x2_ASAP7_75t_L g360 ( .A1(n_91), .A2(n_361), .B1(n_362), .B2(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_91), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_92), .A2(n_96), .B1(n_512), .B2(n_514), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_100), .A2(n_181), .B1(n_387), .B2(n_427), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_101), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_102), .A2(n_107), .B1(n_240), .B2(n_257), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_103), .A2(n_148), .B1(n_317), .B2(n_495), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_104), .A2(n_141), .B1(n_592), .B2(n_593), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_105), .Y(n_661) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_106), .A2(n_182), .B1(n_290), .B2(n_430), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_110), .Y(n_657) );
XNOR2x2_ASAP7_75t_L g236 ( .A(n_114), .B(n_237), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_115), .A2(n_136), .B1(n_288), .B2(n_347), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_118), .Y(n_610) );
INVx2_ASAP7_75t_L g230 ( .A(n_119), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_122), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_125), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_126), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_127), .A2(n_186), .B1(n_349), .B2(n_649), .Y(n_648) );
OA22x2_ASAP7_75t_L g321 ( .A1(n_128), .A2(n_322), .B1(n_323), .B2(n_352), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_128), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_130), .B(n_310), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_131), .B(n_298), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_132), .A2(n_218), .B1(n_429), .B2(n_431), .Y(n_428) );
AND2x6_ASAP7_75t_L g225 ( .A(n_133), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_133), .Y(n_635) );
AO22x2_ASAP7_75t_L g256 ( .A1(n_134), .A2(n_191), .B1(n_247), .B2(n_252), .Y(n_256) );
AOI22xp5_ASAP7_75t_SL g619 ( .A1(n_140), .A2(n_190), .B1(n_350), .B2(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_142), .A2(n_195), .B1(n_341), .B2(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_143), .A2(n_206), .B1(n_300), .B2(n_616), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_144), .B(n_665), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_145), .A2(n_223), .B(n_231), .C(n_643), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_146), .B(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_147), .A2(n_178), .B1(n_302), .B2(n_313), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_149), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_150), .A2(n_202), .B1(n_351), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_152), .A2(n_158), .B1(n_396), .B2(n_398), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_153), .A2(n_221), .B1(n_455), .B2(n_456), .Y(n_480) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_154), .A2(n_198), .B1(n_247), .B2(n_248), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_156), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_157), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_159), .A2(n_175), .B1(n_316), .B2(n_375), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_160), .A2(n_208), .B1(n_350), .B2(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_161), .B(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_164), .A2(n_180), .B1(n_343), .B2(n_344), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_165), .A2(n_183), .B1(n_283), .B2(n_288), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_166), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_167), .Y(n_577) );
INVx1_ASAP7_75t_L g625 ( .A(n_168), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_170), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_171), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_172), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_173), .A2(n_174), .B1(n_288), .B2(n_396), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_176), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_184), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_185), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_187), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_188), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_189), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_191), .B(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_192), .A2(n_220), .B1(n_280), .B2(n_285), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_193), .Y(n_568) );
XOR2xp5_ASAP7_75t_L g644 ( .A(n_194), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g638 ( .A(n_198), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_199), .Y(n_533) );
OA22x2_ASAP7_75t_L g400 ( .A1(n_200), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_400) );
CKINVDCx16_ASAP7_75t_R g401 ( .A(n_200), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_201), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_203), .B(n_503), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_204), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_210), .Y(n_682) );
INVx1_ASAP7_75t_L g247 ( .A(n_211), .Y(n_247) );
INVx1_ASAP7_75t_L g249 ( .A(n_211), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_212), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_213), .A2(n_216), .B1(n_262), .B2(n_398), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_217), .B(n_327), .Y(n_613) );
INVx2_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_226), .Y(n_634) );
OA21x2_ASAP7_75t_L g673 ( .A1(n_227), .A2(n_633), .B(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_523), .B1(n_628), .B2(n_629), .C(n_630), .Y(n_231) );
INVx1_ASAP7_75t_L g628 ( .A(n_232), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B1(n_354), .B2(n_522), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_235), .A2(n_236), .B1(n_320), .B2(n_353), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND4xp75_ASAP7_75t_L g237 ( .A(n_238), .B(n_271), .C(n_291), .D(n_309), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_261), .Y(n_238) );
INVx4_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g510 ( .A(n_241), .Y(n_510) );
INVx4_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx3_ASAP7_75t_L g349 ( .A(n_243), .Y(n_349) );
BUFx3_ASAP7_75t_L g389 ( .A(n_243), .Y(n_389) );
BUFx3_ASAP7_75t_L g452 ( .A(n_243), .Y(n_452) );
INVx2_ASAP7_75t_L g559 ( .A(n_243), .Y(n_559) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_253), .Y(n_243) );
AND2x4_ASAP7_75t_L g258 ( .A(n_244), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g275 ( .A(n_244), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g281 ( .A(n_244), .B(n_265), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_244), .B(n_265), .Y(n_439) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
AND2x2_ASAP7_75t_L g267 ( .A(n_245), .B(n_251), .Y(n_267) );
OR2x2_ASAP7_75t_L g287 ( .A(n_245), .B(n_251), .Y(n_287) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g304 ( .A(n_246), .B(n_256), .Y(n_304) );
AND2x2_ASAP7_75t_L g308 ( .A(n_246), .B(n_251), .Y(n_308) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g252 ( .A(n_249), .Y(n_252) );
AND2x2_ASAP7_75t_L g314 ( .A(n_250), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g380 ( .A(n_250), .Y(n_380) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g270 ( .A(n_251), .Y(n_270) );
AND2x4_ASAP7_75t_L g295 ( .A(n_253), .B(n_286), .Y(n_295) );
AND2x6_ASAP7_75t_L g298 ( .A(n_253), .B(n_267), .Y(n_298) );
INVx1_ASAP7_75t_L g369 ( .A(n_253), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g372 ( .A(n_253), .B(n_267), .Y(n_372) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_254), .B(n_256), .Y(n_260) );
INVx1_ASAP7_75t_L g266 ( .A(n_254), .Y(n_266) );
INVx1_ASAP7_75t_L g277 ( .A(n_254), .Y(n_277) );
INVx1_ASAP7_75t_L g315 ( .A(n_254), .Y(n_315) );
AND2x2_ASAP7_75t_L g276 ( .A(n_255), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g265 ( .A(n_256), .B(n_266), .Y(n_265) );
BUFx2_ASAP7_75t_L g698 ( .A(n_257), .Y(n_698) );
BUFx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g344 ( .A(n_258), .Y(n_344) );
BUFx3_ASAP7_75t_L g394 ( .A(n_258), .Y(n_394) );
INVx1_ASAP7_75t_L g444 ( .A(n_258), .Y(n_444) );
BUFx3_ASAP7_75t_L g542 ( .A(n_258), .Y(n_542) );
BUFx2_ASAP7_75t_SL g649 ( .A(n_258), .Y(n_649) );
AND2x2_ASAP7_75t_L g530 ( .A(n_259), .B(n_380), .Y(n_530) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x6_ASAP7_75t_L g269 ( .A(n_260), .B(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g347 ( .A(n_263), .Y(n_347) );
INVx5_ASAP7_75t_L g391 ( .A(n_263), .Y(n_391) );
INVx4_ASAP7_75t_L g430 ( .A(n_263), .Y(n_430) );
INVx2_ASAP7_75t_L g474 ( .A(n_263), .Y(n_474) );
BUFx3_ASAP7_75t_L g513 ( .A(n_263), .Y(n_513) );
INVx8_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g307 ( .A(n_266), .Y(n_307) );
AND2x4_ASAP7_75t_L g290 ( .A(n_267), .B(n_276), .Y(n_290) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx6_ASAP7_75t_SL g351 ( .A(n_269), .Y(n_351) );
INVx1_ASAP7_75t_SL g514 ( .A(n_269), .Y(n_514) );
INVx1_ASAP7_75t_L g303 ( .A(n_270), .Y(n_303) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_282), .Y(n_271) );
BUFx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_274), .Y(n_517) );
INVx3_ASAP7_75t_L g556 ( .A(n_274), .Y(n_556) );
BUFx3_ASAP7_75t_L g702 ( .A(n_274), .Y(n_702) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_SL g343 ( .A(n_275), .Y(n_343) );
INVx2_ASAP7_75t_L g388 ( .A(n_275), .Y(n_388) );
BUFx2_ASAP7_75t_SL g477 ( .A(n_275), .Y(n_477) );
AND2x6_ASAP7_75t_L g285 ( .A(n_276), .B(n_286), .Y(n_285) );
AND2x6_ASAP7_75t_L g311 ( .A(n_276), .B(n_308), .Y(n_311) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx4f_ASAP7_75t_SL g518 ( .A(n_280), .Y(n_518) );
BUFx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx3_ASAP7_75t_L g341 ( .A(n_281), .Y(n_341) );
BUFx3_ASAP7_75t_L g461 ( .A(n_281), .Y(n_461) );
BUFx3_ASAP7_75t_L g593 ( .A(n_281), .Y(n_593) );
INVx4_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g427 ( .A(n_284), .Y(n_427) );
INVx5_ASAP7_75t_SL g463 ( .A(n_284), .Y(n_463) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_284), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_284), .A2(n_289), .B1(n_654), .B2(n_655), .Y(n_653) );
INVx11_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx11_ASAP7_75t_L g397 ( .A(n_285), .Y(n_397) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g368 ( .A(n_287), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g435 ( .A(n_289), .Y(n_435) );
INVx3_ASAP7_75t_L g602 ( .A(n_289), .Y(n_602) );
INVx6_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx3_ASAP7_75t_L g398 ( .A(n_290), .Y(n_398) );
BUFx3_ASAP7_75t_L g552 ( .A(n_290), .Y(n_552) );
AND2x2_ASAP7_75t_SL g291 ( .A(n_292), .B(n_299), .Y(n_291) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_293), .Y(n_503) );
INVx5_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g329 ( .A(n_294), .Y(n_329) );
INVx2_ASAP7_75t_L g455 ( .A(n_294), .Y(n_455) );
INVx4_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g327 ( .A(n_297), .Y(n_327) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
BUFx4f_ASAP7_75t_L g456 ( .A(n_298), .Y(n_456) );
BUFx2_ASAP7_75t_L g501 ( .A(n_298), .Y(n_501) );
BUFx2_ASAP7_75t_L g665 ( .A(n_298), .Y(n_665) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g505 ( .A(n_301), .Y(n_505) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx2_ASAP7_75t_L g332 ( .A(n_302), .Y(n_332) );
BUFx3_ASAP7_75t_L g458 ( .A(n_302), .Y(n_458) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x4_ASAP7_75t_L g313 ( .A(n_304), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g318 ( .A(n_304), .B(n_319), .Y(n_318) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_304), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g507 ( .A(n_305), .Y(n_507) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g466 ( .A(n_306), .Y(n_466) );
BUFx2_ASAP7_75t_SL g616 ( .A(n_306), .Y(n_616) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g384 ( .A(n_307), .Y(n_384) );
INVx1_ASAP7_75t_L g383 ( .A(n_308), .Y(n_383) );
INVx3_ASAP7_75t_L g413 ( .A(n_310), .Y(n_413) );
BUFx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx4_ASAP7_75t_L g335 ( .A(n_311), .Y(n_335) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_311), .Y(n_465) );
INVx2_ASAP7_75t_L g573 ( .A(n_311), .Y(n_573) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_313), .Y(n_331) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_313), .Y(n_375) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_313), .Y(n_485) );
BUFx4f_ASAP7_75t_SL g571 ( .A(n_313), .Y(n_571) );
INVx1_ASAP7_75t_L g319 ( .A(n_315), .Y(n_319) );
INVx1_ASAP7_75t_L g580 ( .A(n_316), .Y(n_580) );
BUFx4f_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g418 ( .A(n_317), .Y(n_418) );
BUFx12f_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_318), .Y(n_498) );
INVx1_ASAP7_75t_L g353 ( .A(n_320), .Y(n_353) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g352 ( .A(n_323), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_324), .B(n_338), .Y(n_323) );
NOR2xp67_ASAP7_75t_SL g324 ( .A(n_325), .B(n_333), .Y(n_324) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .C(n_330), .Y(n_325) );
OAI21xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_336), .B(n_337), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_335), .A2(n_533), .B(n_534), .Y(n_532) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_335), .A2(n_610), .B(n_611), .Y(n_609) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_335), .A2(n_661), .B(n_662), .Y(n_660) );
NOR2x1_ASAP7_75t_L g338 ( .A(n_339), .B(n_345), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g431 ( .A(n_351), .Y(n_431) );
BUFx2_ASAP7_75t_L g705 ( .A(n_351), .Y(n_705) );
INVx1_ASAP7_75t_L g522 ( .A(n_354), .Y(n_522) );
XOR2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_445), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_399), .B2(n_400), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND3x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_385), .C(n_392), .Y(n_363) );
NOR3xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_373), .C(n_377), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_370), .B2(n_371), .Y(n_365) );
BUFx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_368), .Y(n_408) );
INVx2_ASAP7_75t_L g567 ( .A(n_368), .Y(n_567) );
BUFx3_ASAP7_75t_L g410 ( .A(n_371), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_371), .A2(n_565), .B1(n_566), .B2(n_568), .Y(n_564) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g597 ( .A(n_372), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
BUFx2_ASAP7_75t_L g416 ( .A(n_375), .Y(n_416) );
INVx4_ASAP7_75t_L g496 ( .A(n_375), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B1(n_381), .B2(n_382), .Y(n_377) );
OAI22xp33_ASAP7_75t_SL g419 ( .A1(n_379), .A2(n_420), .B1(n_421), .B2(n_423), .Y(n_419) );
INVx4_ASAP7_75t_L g576 ( .A(n_379), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_379), .A2(n_582), .B1(n_693), .B2(n_694), .Y(n_692) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_382), .Y(n_422) );
BUFx2_ASAP7_75t_L g582 ( .A(n_382), .Y(n_582) );
OR2x6_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx3_ASAP7_75t_L g592 ( .A(n_388), .Y(n_592) );
INVx1_ASAP7_75t_L g442 ( .A(n_389), .Y(n_442) );
BUFx2_ASAP7_75t_L g704 ( .A(n_391), .Y(n_704) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx4_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g624 ( .A(n_397), .Y(n_624) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_424), .Y(n_403) );
NOR3xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_412), .C(n_419), .Y(n_404) );
OAI22xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_409), .B1(n_410), .B2(n_411), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_408), .A2(n_682), .B1(n_683), .B2(n_684), .Y(n_681) );
OAI21xp33_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B(n_415), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g482 ( .A1(n_413), .A2(n_483), .B(n_484), .Y(n_482) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_432), .C(n_440), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g620 ( .A(n_430), .Y(n_620) );
INVx2_ASAP7_75t_L g652 ( .A(n_430), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_436), .B2(n_437), .Y(n_432) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_437), .A2(n_556), .B1(n_657), .B2(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_440) );
OAI221xp5_ASAP7_75t_SL g558 ( .A1(n_444), .A2(n_559), .B1(n_560), .B2(n_561), .C(n_562), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B1(n_467), .B2(n_468), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND5xp2_ASAP7_75t_SL g449 ( .A(n_450), .B(n_451), .C(n_453), .D(n_459), .E(n_464), .Y(n_449) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_454), .B(n_457), .Y(n_453) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
BUFx3_ASAP7_75t_L g557 ( .A(n_461), .Y(n_557) );
INVx2_ASAP7_75t_L g492 ( .A(n_465), .Y(n_492) );
INVx2_ASAP7_75t_SL g686 ( .A(n_465), .Y(n_686) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AO22x1_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_486), .B1(n_487), .B2(n_521), .Y(n_468) );
INVx1_ASAP7_75t_SL g521 ( .A(n_469), .Y(n_521) );
NOR4xp75_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .C(n_479), .D(n_482), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_472), .B(n_473), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_476), .B(n_478), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_480), .B(n_481), .Y(n_479) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_485), .Y(n_689) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g520 ( .A(n_489), .Y(n_520) );
NAND3x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_508), .C(n_515), .Y(n_489) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_491), .B(n_499), .Y(n_490) );
OAI21xp5_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_493), .B(n_494), .Y(n_491) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx4f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .C(n_504), .Y(n_499) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
INVx1_ASAP7_75t_L g629 ( .A(n_523), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_544), .B2(n_627), .Y(n_523) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
XOR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_543), .Y(n_525) );
NAND3x1_ASAP7_75t_SL g526 ( .A(n_527), .B(n_531), .C(n_539), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_532), .B(n_535), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .C(n_538), .Y(n_535) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_SL g627 ( .A(n_544), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_585), .B1(n_586), .B2(n_626), .Y(n_544) );
INVx2_ASAP7_75t_L g626 ( .A(n_545), .Y(n_626) );
INVx1_ASAP7_75t_L g583 ( .A(n_546), .Y(n_583) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_547), .B(n_563), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_558), .Y(n_547) );
OAI221xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_550), .B1(n_551), .B2(n_553), .C(n_554), .Y(n_548) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NOR3xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_569), .C(n_578), .Y(n_563) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
OAI222xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_572), .B1(n_573), .B2(n_574), .C1(n_575), .C2(n_577), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B1(n_581), .B2(n_582), .Y(n_578) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
XNOR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_606), .Y(n_586) );
XOR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_605), .Y(n_587) );
NAND4xp75_ASAP7_75t_L g588 ( .A(n_589), .B(n_594), .C(n_600), .D(n_604), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OA211x2_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_598), .C(n_599), .Y(n_594) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_SL g684 ( .A(n_597), .Y(n_684) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
XOR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_625), .Y(n_606) );
NAND3x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_617), .C(n_621), .Y(n_607) );
NOR2x1_ASAP7_75t_L g608 ( .A(n_609), .B(n_612), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .C(n_615), .Y(n_612) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
NOR2x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .Y(n_631) );
OR2x2_ASAP7_75t_SL g709 ( .A(n_632), .B(n_637), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_634), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_634), .B(n_672), .Y(n_674) );
CKINVDCx16_ASAP7_75t_R g672 ( .A(n_635), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
OAI322xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_668), .A3(n_669), .B1(n_673), .B2(n_675), .C1(n_676), .C2(n_707), .Y(n_643) );
AND2x2_ASAP7_75t_SL g645 ( .A(n_646), .B(n_659), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_653), .C(n_656), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .C(n_667), .Y(n_663) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g706 ( .A(n_679), .Y(n_706) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_695), .Y(n_679) );
NOR3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_685), .C(n_692), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_688), .B2(n_690), .C(n_691), .Y(n_685) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_700), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_708), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_709), .Y(n_708) );
endmodule