module real_aes_9117_n_367 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_367);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_367;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_1067;
wire n_518;
wire n_792;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_1040;
wire n_415;
wire n_572;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_370;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_1098;
wire n_824;
wire n_875;
wire n_467;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_976;
wire n_1049;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_369;
wire n_1070;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_996;
wire n_523;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_973;
wire n_1081;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_1006;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_1079;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1028;
wire n_727;
wire n_1014;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_691;
wire n_765;
wire n_481;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_717;
wire n_456;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_823;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_1045;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_968;
wire n_743;
wire n_710;
wire n_393;
wire n_652;
wire n_1097;
wire n_703;
wire n_500;
wire n_601;
wire n_1101;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g773 ( .A1(n_0), .A2(n_161), .B1(n_651), .B2(n_774), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_1), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_2), .B(n_475), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_3), .B(n_470), .Y(n_1011) );
XOR2x2_ASAP7_75t_L g728 ( .A(n_4), .B(n_729), .Y(n_728) );
OA22x2_ASAP7_75t_L g382 ( .A1(n_5), .A2(n_383), .B1(n_384), .B2(n_476), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_5), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_6), .A2(n_557), .B1(n_591), .B2(n_592), .Y(n_556) );
INVx1_ASAP7_75t_L g592 ( .A(n_6), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_7), .A2(n_271), .B1(n_526), .B2(n_612), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_8), .A2(n_334), .B1(n_724), .B2(n_856), .Y(n_1035) );
AOI22xp5_ASAP7_75t_SL g649 ( .A1(n_9), .A2(n_364), .B1(n_650), .B2(n_651), .Y(n_649) );
AO22x2_ASAP7_75t_L g401 ( .A1(n_10), .A2(n_205), .B1(n_393), .B2(n_398), .Y(n_401) );
INVx1_ASAP7_75t_L g1060 ( .A(n_10), .Y(n_1060) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_11), .Y(n_885) );
AOI22xp33_ASAP7_75t_SL g959 ( .A1(n_12), .A2(n_192), .B1(n_722), .B2(n_734), .Y(n_959) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_13), .A2(n_283), .B1(n_466), .B2(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_SL g643 ( .A1(n_14), .A2(n_230), .B1(n_616), .B2(n_644), .Y(n_643) );
AO22x1_ASAP7_75t_L g695 ( .A1(n_15), .A2(n_696), .B1(n_726), .B2(n_727), .Y(n_695) );
INVx1_ASAP7_75t_L g726 ( .A(n_15), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_16), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_17), .A2(n_24), .B1(n_612), .B2(n_934), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_18), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_19), .A2(n_366), .B1(n_665), .B2(n_789), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_20), .A2(n_358), .B1(n_426), .B2(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g911 ( .A(n_21), .Y(n_911) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_22), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_23), .A2(n_355), .B1(n_549), .B2(n_737), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_25), .A2(n_250), .B1(n_427), .B2(n_499), .Y(n_910) );
AOI22xp33_ASAP7_75t_SL g1012 ( .A1(n_26), .A2(n_319), .B1(n_678), .B2(n_864), .Y(n_1012) );
INVx1_ASAP7_75t_L g748 ( .A(n_27), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g639 ( .A1(n_28), .A2(n_163), .B1(n_640), .B2(n_641), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_29), .A2(n_324), .B1(n_431), .B2(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_30), .A2(n_86), .B1(n_458), .B2(n_494), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_31), .A2(n_101), .B1(n_544), .B2(n_572), .Y(n_571) );
AO22x2_ASAP7_75t_L g403 ( .A1(n_32), .A2(n_107), .B1(n_393), .B2(n_394), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g1014 ( .A(n_33), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_34), .A2(n_186), .B1(n_426), .B2(n_429), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g986 ( .A1(n_35), .A2(n_93), .B1(n_682), .B2(n_987), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_36), .A2(n_261), .B1(n_566), .B2(n_956), .Y(n_955) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_37), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g775 ( .A1(n_38), .A2(n_308), .B1(n_544), .B2(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_39), .A2(n_210), .B1(n_599), .B2(n_600), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_40), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g927 ( .A(n_41), .Y(n_927) );
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_42), .A2(n_256), .B1(n_422), .B2(n_437), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_43), .A2(n_212), .B1(n_600), .B2(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_44), .B(n_525), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_45), .A2(n_253), .B1(n_524), .B2(n_525), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_46), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_47), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_48), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_49), .A2(n_180), .B1(n_525), .B2(n_633), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_50), .A2(n_347), .B1(n_739), .B2(n_917), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_51), .B(n_747), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g1018 ( .A1(n_52), .A2(n_304), .B1(n_650), .B2(n_956), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_53), .A2(n_199), .B1(n_664), .B2(n_665), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_54), .A2(n_173), .B1(n_426), .B2(n_565), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g1074 ( .A(n_55), .Y(n_1074) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_56), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_57), .A2(n_350), .B1(n_412), .B2(n_427), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_58), .A2(n_279), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g654 ( .A(n_59), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_60), .A2(n_102), .B1(n_668), .B2(n_719), .Y(n_718) );
AOI222xp33_ASAP7_75t_L g621 ( .A1(n_61), .A2(n_190), .B1(n_222), .B2(n_446), .C1(n_622), .C2(n_623), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_62), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_63), .A2(n_254), .B1(n_420), .B2(n_549), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_64), .A2(n_264), .B1(n_615), .B2(n_653), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_65), .A2(n_92), .B1(n_410), .B2(n_420), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_66), .A2(n_239), .B1(n_452), .B2(n_464), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_67), .A2(n_215), .B1(n_599), .B2(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_68), .A2(n_147), .B1(n_644), .B2(n_651), .Y(n_1019) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_69), .Y(n_561) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_70), .A2(n_368), .B(n_376), .C(n_1062), .Y(n_367) );
AOI22xp5_ASAP7_75t_SL g645 ( .A1(n_71), .A2(n_236), .B1(n_646), .B2(n_647), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_72), .A2(n_232), .B1(n_549), .B2(n_551), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_73), .Y(n_849) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_74), .A2(n_263), .B1(n_404), .B2(n_498), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_75), .A2(n_287), .B1(n_602), .B2(n_665), .Y(n_957) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_76), .A2(n_201), .B1(n_440), .B2(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_77), .A2(n_113), .B1(n_615), .B2(n_616), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g902 ( .A(n_78), .Y(n_902) );
AO22x2_ASAP7_75t_L g397 ( .A1(n_79), .A2(n_243), .B1(n_393), .B2(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g1057 ( .A(n_79), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_80), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_81), .A2(n_241), .B1(n_435), .B2(n_620), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g1067 ( .A(n_82), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_83), .A2(n_88), .B1(n_429), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_84), .A2(n_170), .B1(n_612), .B2(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_SL g994 ( .A1(n_85), .A2(n_301), .B1(n_404), .B2(n_854), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_87), .A2(n_362), .B1(n_618), .B2(n_787), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_89), .Y(n_563) );
AOI22xp5_ASAP7_75t_SL g652 ( .A1(n_90), .A2(n_196), .B1(n_420), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_91), .A2(n_280), .B1(n_618), .B2(n_619), .Y(n_617) );
AOI211xp5_ASAP7_75t_L g995 ( .A1(n_94), .A2(n_644), .B(n_996), .C(n_1001), .Y(n_995) );
AOI22xp33_ASAP7_75t_SL g989 ( .A1(n_95), .A2(n_269), .B1(n_463), .B2(n_466), .Y(n_989) );
AOI222xp33_ASAP7_75t_L g796 ( .A1(n_96), .A2(n_214), .B1(n_226), .B2(n_446), .C1(n_466), .C2(n_623), .Y(n_796) );
INVx1_ASAP7_75t_L g935 ( .A(n_97), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_98), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_99), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_100), .A2(n_181), .B1(n_488), .B2(n_612), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_103), .A2(n_187), .B1(n_470), .B2(n_473), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_104), .A2(n_657), .B1(n_687), .B2(n_688), .Y(n_656) );
INVx1_ASAP7_75t_L g687 ( .A(n_104), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_105), .A2(n_112), .B1(n_622), .B2(n_623), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_106), .A2(n_166), .B1(n_451), .B2(n_464), .Y(n_973) );
INVx1_ASAP7_75t_L g1061 ( .A(n_107), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_108), .A2(n_235), .B1(n_619), .B2(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_109), .B(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_110), .Y(n_859) );
XOR2xp5_ASAP7_75t_L g784 ( .A(n_111), .B(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_114), .A2(n_315), .B1(n_464), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_115), .A2(n_184), .B1(n_388), .B2(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_116), .A2(n_341), .B1(n_787), .B2(n_856), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_117), .B(n_610), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_118), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_119), .A2(n_174), .B1(n_541), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_120), .A2(n_298), .B1(n_742), .B2(n_743), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g767 ( .A1(n_121), .A2(n_194), .B1(n_768), .B2(n_770), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_122), .A2(n_224), .B1(n_653), .B2(n_1079), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_123), .A2(n_134), .B1(n_488), .B2(n_524), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_124), .A2(n_310), .B1(n_647), .B2(n_739), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_125), .A2(n_317), .B1(n_572), .B2(n_618), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_126), .A2(n_225), .B1(n_464), .B2(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_127), .A2(n_231), .B1(n_463), .B2(n_466), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_128), .A2(n_351), .B1(n_993), .B2(n_1086), .Y(n_1085) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_129), .A2(n_330), .B1(n_488), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_130), .A2(n_191), .B1(n_435), .B2(n_440), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_131), .A2(n_175), .B1(n_473), .B2(n_610), .Y(n_1038) );
XNOR2x2_ASAP7_75t_L g1029 ( .A(n_132), .B(n_1030), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_133), .A2(n_143), .B1(n_599), .B2(n_854), .Y(n_853) );
OA22x2_ASAP7_75t_L g1005 ( .A1(n_135), .A2(n_1006), .B1(n_1007), .B2(n_1024), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_135), .Y(n_1006) );
INVx1_ASAP7_75t_L g508 ( .A(n_136), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_137), .B(n_475), .Y(n_906) );
AND2x6_ASAP7_75t_L g370 ( .A(n_138), .B(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_138), .Y(n_1054) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_139), .A2(n_354), .B1(n_650), .B2(n_665), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_140), .B(n_931), .Y(n_930) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_141), .B(n_609), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_142), .Y(n_706) );
AOI22xp33_ASAP7_75t_SL g892 ( .A1(n_144), .A2(n_335), .B1(n_549), .B2(n_787), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_145), .A2(n_177), .B1(n_566), .B2(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g764 ( .A(n_146), .B(n_765), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_148), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g975 ( .A1(n_149), .A2(n_167), .B1(n_503), .B2(n_976), .Y(n_975) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_150), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_151), .Y(n_952) );
AOI222xp33_ASAP7_75t_L g1040 ( .A1(n_152), .A2(n_193), .B1(n_325), .B2(n_588), .C1(n_704), .C2(n_747), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_153), .A2(n_285), .B1(n_599), .B2(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g990 ( .A1(n_154), .A2(n_217), .B1(n_610), .B2(n_765), .Y(n_990) );
AO22x2_ASAP7_75t_L g392 ( .A1(n_155), .A2(n_233), .B1(n_393), .B2(n_394), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g1058 ( .A(n_155), .B(n_1059), .Y(n_1058) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_156), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g1002 ( .A(n_157), .Y(n_1002) );
AOI22xp33_ASAP7_75t_SL g909 ( .A1(n_158), .A2(n_274), .B1(n_389), .B2(n_414), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_159), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g992 ( .A1(n_160), .A2(n_252), .B1(n_787), .B2(n_993), .Y(n_992) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_162), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_164), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_165), .A2(n_169), .B1(n_640), .B2(n_678), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_168), .A2(n_244), .B1(n_427), .B2(n_618), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_171), .A2(n_300), .B1(n_426), .B2(n_1084), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_172), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_176), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_178), .Y(n_948) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_179), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_182), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_183), .A2(n_284), .B1(n_619), .B2(n_739), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_185), .B(n_637), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_188), .A2(n_234), .B1(n_412), .B2(n_427), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_189), .A2(n_282), .B1(n_572), .B2(n_667), .Y(n_1081) );
XNOR2xp5_ASAP7_75t_L g981 ( .A(n_195), .B(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_197), .A2(n_223), .B1(n_616), .B2(n_826), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g889 ( .A1(n_198), .A2(n_216), .B1(n_504), .B2(n_647), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_200), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_202), .A2(n_320), .B1(n_776), .B2(n_851), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_203), .A2(n_327), .B1(n_667), .B2(n_668), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_204), .A2(n_221), .B1(n_665), .B2(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_206), .B(n_609), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_207), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_208), .A2(n_309), .B1(n_566), .B2(n_600), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_209), .A2(n_249), .B1(n_431), .B2(n_506), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_211), .B(n_776), .Y(n_1000) );
OA22x2_ASAP7_75t_L g873 ( .A1(n_213), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_213), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_218), .A2(n_237), .B1(n_498), .B2(n_602), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_219), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_220), .A2(n_311), .B1(n_429), .B2(n_600), .Y(n_1032) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_227), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_228), .A2(n_278), .B1(n_498), .B2(n_506), .Y(n_964) );
INVx2_ASAP7_75t_L g375 ( .A(n_229), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_238), .A2(n_267), .B1(n_641), .B2(n_934), .Y(n_933) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_240), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g1071 ( .A(n_242), .Y(n_1071) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_245), .A2(n_842), .B1(n_870), .B2(n_871), .Y(n_841) );
INVx1_ASAP7_75t_L g870 ( .A(n_245), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g945 ( .A(n_246), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_247), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_248), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_251), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_255), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_257), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_258), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_259), .Y(n_815) );
INVx1_ASAP7_75t_L g1098 ( .A(n_260), .Y(n_1098) );
AOI22x1_ASAP7_75t_L g1099 ( .A1(n_260), .A2(n_1064), .B1(n_1089), .B2(n_1098), .Y(n_1099) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_262), .Y(n_968) );
OA22x2_ASAP7_75t_L g806 ( .A1(n_265), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_806) );
CKINVDCx16_ASAP7_75t_R g807 ( .A(n_265), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_266), .B(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_268), .A2(n_337), .B1(n_647), .B2(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g393 ( .A(n_270), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_270), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_272), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_273), .A2(n_321), .B1(n_619), .B2(n_719), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_275), .B(n_470), .Y(n_932) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_276), .A2(n_312), .B1(n_503), .B2(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_277), .A2(n_352), .B1(n_388), .B2(n_404), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_281), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_286), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_288), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_289), .A2(n_1064), .B1(n_1088), .B2(n_1089), .Y(n_1063) );
CKINVDCx20_ASAP7_75t_R g1088 ( .A(n_289), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_290), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_291), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_292), .A2(n_756), .B1(n_757), .B2(n_781), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_292), .Y(n_756) );
XNOR2x1_ASAP7_75t_L g941 ( .A(n_293), .B(n_942), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_294), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_295), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_296), .A2(n_345), .B1(n_467), .B2(n_640), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_297), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_299), .Y(n_978) );
AND2x2_ASAP7_75t_L g374 ( .A(n_302), .B(n_375), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_303), .Y(n_1075) );
INVx1_ASAP7_75t_L g371 ( .A(n_305), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_306), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_307), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_313), .A2(n_360), .B1(n_458), .B2(n_466), .Y(n_949) );
AOI22xp33_ASAP7_75t_SL g1021 ( .A1(n_314), .A2(n_323), .B1(n_420), .B2(n_1022), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_316), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_318), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_322), .B(n_742), .Y(n_971) );
CKINVDCx20_ASAP7_75t_R g1072 ( .A(n_326), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_328), .A2(n_357), .B1(n_526), .B2(n_612), .Y(n_969) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_329), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_331), .B(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_332), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_333), .A2(n_365), .B1(n_742), .B2(n_743), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g928 ( .A1(n_336), .A2(n_343), .B1(n_524), .B2(n_588), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_338), .A2(n_348), .B1(n_420), .B2(n_956), .Y(n_1036) );
XNOR2x1_ASAP7_75t_L g509 ( .A(n_339), .B(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_340), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g997 ( .A(n_342), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_344), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_346), .B(n_475), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_349), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_353), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_356), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_359), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_361), .B(n_637), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_363), .Y(n_711) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_371), .Y(n_1053) );
OAI21xp5_ASAP7_75t_L g1096 ( .A1(n_372), .A2(n_1052), .B(n_1097), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_799), .B1(n_1047), .B2(n_1048), .C(n_1049), .Y(n_376) );
INVx1_ASAP7_75t_L g1047 ( .A(n_377), .Y(n_1047) );
AOI22xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_690), .B1(n_691), .B2(n_798), .Y(n_377) );
INVx1_ASAP7_75t_L g798 ( .A(n_378), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_552), .B2(n_553), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B1(n_477), .B2(n_478), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g476 ( .A(n_384), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_443), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_424), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_409), .Y(n_386) );
BUFx4f_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g725 ( .A(n_389), .Y(n_725) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g498 ( .A(n_390), .Y(n_498) );
BUFx3_ASAP7_75t_L g566 ( .A(n_390), .Y(n_566) );
BUFx3_ASAP7_75t_L g650 ( .A(n_390), .Y(n_650) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_399), .Y(n_390) );
AND2x2_ASAP7_75t_L g439 ( .A(n_391), .B(n_423), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_391), .B(n_399), .Y(n_834) );
NAND2xp5_ASAP7_75t_SL g999 ( .A(n_391), .B(n_423), .Y(n_999) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_392), .B(n_397), .Y(n_408) );
INVx2_ASAP7_75t_L g418 ( .A(n_392), .Y(n_418) );
AND2x2_ASAP7_75t_L g455 ( .A(n_392), .B(n_401), .Y(n_455) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_395), .Y(n_398) );
INVx1_ASAP7_75t_L g468 ( .A(n_396), .Y(n_468) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g419 ( .A(n_397), .Y(n_419) );
AND2x2_ASAP7_75t_L g433 ( .A(n_397), .B(n_418), .Y(n_433) );
INVx1_ASAP7_75t_L g454 ( .A(n_397), .Y(n_454) );
AND2x4_ASAP7_75t_L g406 ( .A(n_399), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g428 ( .A(n_399), .B(n_417), .Y(n_428) );
AND2x4_ASAP7_75t_L g432 ( .A(n_399), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
OR2x2_ASAP7_75t_L g416 ( .A(n_400), .B(n_403), .Y(n_416) );
AND2x2_ASAP7_75t_L g423 ( .A(n_400), .B(n_403), .Y(n_423) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g448 ( .A(n_401), .B(n_403), .Y(n_448) );
AND2x2_ASAP7_75t_L g453 ( .A(n_402), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g507 ( .A(n_402), .Y(n_507) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g442 ( .A(n_403), .Y(n_442) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI221xp5_ASAP7_75t_SL g567 ( .A1(n_405), .A2(n_568), .B1(n_569), .B2(n_570), .C(n_571), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_405), .A2(n_836), .B1(n_837), .B2(n_838), .Y(n_835) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g499 ( .A(n_406), .Y(n_499) );
BUFx3_ASAP7_75t_L g600 ( .A(n_406), .Y(n_600) );
BUFx2_ASAP7_75t_L g651 ( .A(n_406), .Y(n_651) );
BUFx3_ASAP7_75t_L g665 ( .A(n_406), .Y(n_665) );
BUFx2_ASAP7_75t_SL g848 ( .A(n_406), .Y(n_848) );
BUFx2_ASAP7_75t_SL g917 ( .A(n_406), .Y(n_917) );
AND2x2_ASAP7_75t_L g506 ( .A(n_407), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x6_ASAP7_75t_L g441 ( .A(n_408), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx5_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_413), .Y(n_560) );
INVx2_ASAP7_75t_L g599 ( .A(n_413), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_413), .A2(n_421), .B1(n_920), .B2(n_921), .Y(n_919) );
INVx4_ASAP7_75t_L g956 ( .A(n_413), .Y(n_956) );
INVx2_ASAP7_75t_SL g976 ( .A(n_413), .Y(n_976) );
INVx11_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx11_ASAP7_75t_L g550 ( .A(n_414), .Y(n_550) );
AND2x6_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
AND2x4_ASAP7_75t_L g472 ( .A(n_415), .B(n_433), .Y(n_472) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g515 ( .A(n_416), .B(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_L g422 ( .A(n_417), .B(n_423), .Y(n_422) );
AND2x6_ASAP7_75t_L g447 ( .A(n_417), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g615 ( .A(n_421), .Y(n_615) );
INVx2_ASAP7_75t_L g722 ( .A(n_421), .Y(n_722) );
INVx2_ASAP7_75t_L g732 ( .A(n_421), .Y(n_732) );
INVx6_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g503 ( .A(n_422), .Y(n_503) );
BUFx3_ASAP7_75t_L g551 ( .A(n_422), .Y(n_551) );
BUFx3_ASAP7_75t_L g787 ( .A(n_422), .Y(n_787) );
AND2x6_ASAP7_75t_L g475 ( .A(n_423), .B(n_433), .Y(n_475) );
NAND2x1p5_ASAP7_75t_L g520 ( .A(n_423), .B(n_433), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_434), .Y(n_424) );
BUFx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g542 ( .A(n_427), .Y(n_542) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_427), .Y(n_779) );
BUFx3_ASAP7_75t_L g856 ( .A(n_427), .Y(n_856) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g603 ( .A(n_428), .Y(n_603) );
BUFx2_ASAP7_75t_SL g644 ( .A(n_428), .Y(n_644) );
BUFx2_ASAP7_75t_SL g737 ( .A(n_428), .Y(n_737) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g774 ( .A(n_430), .Y(n_774) );
INVx4_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g568 ( .A(n_432), .Y(n_568) );
BUFx3_ASAP7_75t_L g616 ( .A(n_432), .Y(n_616) );
BUFx3_ASAP7_75t_L g739 ( .A(n_432), .Y(n_739) );
BUFx3_ASAP7_75t_L g789 ( .A(n_432), .Y(n_789) );
INVx1_ASAP7_75t_L g516 ( .A(n_433), .Y(n_516) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g646 ( .A(n_437), .Y(n_646) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_437), .Y(n_719) );
INVx4_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx5_ASAP7_75t_L g504 ( .A(n_438), .Y(n_504) );
BUFx3_ASAP7_75t_L g545 ( .A(n_438), .Y(n_545) );
INVx3_ASAP7_75t_L g618 ( .A(n_438), .Y(n_618) );
INVx2_ASAP7_75t_L g734 ( .A(n_438), .Y(n_734) );
INVx1_ASAP7_75t_L g1022 ( .A(n_438), .Y(n_1022) );
INVx8_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g572 ( .A(n_441), .Y(n_572) );
INVx6_ASAP7_75t_SL g620 ( .A(n_441), .Y(n_620) );
INVx1_ASAP7_75t_SL g776 ( .A(n_441), .Y(n_776) );
INVx1_ASAP7_75t_L g465 ( .A(n_442), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_461), .Y(n_443) );
OAI222xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_449), .B1(n_450), .B2(n_456), .C1(n_457), .C2(n_460), .Y(n_444) );
OAI222xp33_ASAP7_75t_L g702 ( .A1(n_445), .A2(n_703), .B1(n_705), .B2(n_706), .C1(n_707), .C2(n_709), .Y(n_702) );
OAI222xp33_ASAP7_75t_L g865 ( .A1(n_445), .A2(n_677), .B1(n_866), .B2(n_867), .C1(n_868), .C2(n_869), .Y(n_865) );
INVx2_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g760 ( .A(n_446), .Y(n_760) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g486 ( .A(n_447), .Y(n_486) );
INVx4_ASAP7_75t_L g630 ( .A(n_447), .Y(n_630) );
BUFx3_ASAP7_75t_L g747 ( .A(n_447), .Y(n_747) );
AND2x4_ASAP7_75t_L g467 ( .A(n_448), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g536 ( .A(n_448), .Y(n_536) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g580 ( .A(n_451), .Y(n_580) );
BUFx4f_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_452), .Y(n_494) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_452), .Y(n_524) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_452), .Y(n_678) );
BUFx2_ASAP7_75t_L g704 ( .A(n_452), .Y(n_704) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
INVx1_ASAP7_75t_L g459 ( .A(n_454), .Y(n_459) );
AND2x4_ASAP7_75t_L g458 ( .A(n_455), .B(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g464 ( .A(n_455), .B(n_465), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g531 ( .A(n_455), .B(n_507), .Y(n_531) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx12f_ASAP7_75t_L g488 ( .A(n_458), .Y(n_488) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_458), .Y(n_526) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_458), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_469), .Y(n_461) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g640 ( .A(n_464), .Y(n_640) );
INVx1_ASAP7_75t_L g769 ( .A(n_464), .Y(n_769) );
BUFx2_ASAP7_75t_L g864 ( .A(n_464), .Y(n_864) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_467), .Y(n_612) );
BUFx2_ASAP7_75t_SL g641 ( .A(n_467), .Y(n_641) );
INVx1_ASAP7_75t_L g537 ( .A(n_468), .Y(n_537) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g491 ( .A(n_471), .Y(n_491) );
INVx5_ASAP7_75t_L g610 ( .A(n_471), .Y(n_610) );
INVx2_ASAP7_75t_L g742 ( .A(n_471), .Y(n_742) );
INVx4_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g637 ( .A(n_474), .Y(n_637) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
BUFx4f_ASAP7_75t_L g743 ( .A(n_475), .Y(n_743) );
BUFx2_ASAP7_75t_L g765 ( .A(n_475), .Y(n_765) );
BUFx2_ASAP7_75t_L g931 ( .A(n_475), .Y(n_931) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
XNOR2x1_ASAP7_75t_SL g478 ( .A(n_479), .B(n_509), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AO22x2_ASAP7_75t_L g783 ( .A1(n_480), .A2(n_481), .B1(n_784), .B2(n_797), .Y(n_783) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
XOR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_508), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_483), .B(n_495), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_489), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_487), .Y(n_484) );
OAI21xp33_ASAP7_75t_SL g521 ( .A1(n_486), .A2(n_522), .B(n_523), .Y(n_521) );
OAI222xp33_ASAP7_75t_L g579 ( .A1(n_486), .A2(n_580), .B1(n_581), .B2(n_582), .C1(n_583), .C2(n_584), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g1066 ( .A1(n_486), .A2(n_677), .B1(n_1067), .B2(n_1068), .C(n_1069), .Y(n_1066) );
BUFx4f_ASAP7_75t_SL g588 ( .A(n_488), .Y(n_588) );
INVx2_ASAP7_75t_L g624 ( .A(n_488), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .C(n_493), .Y(n_489) );
BUFx6f_ASAP7_75t_L g987 ( .A(n_494), .Y(n_987) );
NOR2x1_ASAP7_75t_L g495 ( .A(n_496), .B(n_501), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_500), .Y(n_496) );
INVx2_ASAP7_75t_L g1080 ( .A(n_499), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .Y(n_501) );
INVx3_ASAP7_75t_L g562 ( .A(n_503), .Y(n_562) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_504), .Y(n_667) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_538), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .C(n_527), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_517), .B2(n_518), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_514), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_514), .A2(n_519), .B1(n_879), .B2(n_880), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_514), .A2(n_673), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
BUFx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g577 ( .A(n_515), .Y(n_577) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_515), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_515), .A2(n_673), .B1(n_945), .B2(n_946), .Y(n_944) );
OAI22xp5_ASAP7_75t_SL g811 ( .A1(n_518), .A2(n_812), .B1(n_815), .B2(n_816), .Y(n_811) );
BUFx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_519), .A2(n_575), .B1(n_576), .B2(n_578), .Y(n_574) );
INVx2_ASAP7_75t_L g861 ( .A(n_519), .Y(n_861) );
BUFx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g607 ( .A(n_520), .Y(n_607) );
BUFx2_ASAP7_75t_L g622 ( .A(n_524), .Y(n_622) );
INVx4_ASAP7_75t_L g634 ( .A(n_524), .Y(n_634) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B1(n_532), .B2(n_533), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_529), .A2(n_684), .B1(n_685), .B2(n_686), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_529), .A2(n_533), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
INVx3_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g583 ( .A(n_530), .Y(n_583) );
INVx4_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx3_ASAP7_75t_L g712 ( .A(n_531), .Y(n_712) );
OAI22xp33_ASAP7_75t_SL g820 ( .A1(n_531), .A2(n_686), .B1(n_821), .B2(n_822), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_531), .A2(n_535), .B1(n_885), .B2(n_886), .Y(n_884) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g686 ( .A(n_534), .Y(n_686) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g590 ( .A(n_535), .Y(n_590) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_546), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_542), .A2(n_832), .B1(n_923), .B2(n_924), .Y(n_922) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx4_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_SL g653 ( .A(n_550), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g1001 ( .A(n_550), .B(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1087 ( .A(n_551), .Y(n_1087) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_SL g553 ( .A1(n_554), .A2(n_555), .B1(n_656), .B2(n_689), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_593), .B1(n_594), .B2(n_655), .Y(n_555) );
INVx2_ASAP7_75t_L g655 ( .A(n_556), .Y(n_655) );
INVx1_ASAP7_75t_L g591 ( .A(n_557), .Y(n_591) );
AND2x2_ASAP7_75t_SL g557 ( .A(n_558), .B(n_573), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_567), .Y(n_558) );
OAI221xp5_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_561), .B1(n_562), .B2(n_563), .C(n_564), .Y(n_559) );
BUFx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g664 ( .A(n_568), .Y(n_664) );
INVx1_ASAP7_75t_L g717 ( .A(n_568), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_579), .C(n_585), .Y(n_573) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g700 ( .A(n_577), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g950 ( .A1(n_583), .A2(n_703), .B1(n_951), .B2(n_952), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_589), .B2(n_590), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
XNOR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_626), .Y(n_594) );
XOR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_625), .Y(n_595) );
NAND4xp75_ASAP7_75t_L g596 ( .A(n_597), .B(n_604), .C(n_613), .D(n_621), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
INVx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx3_ASAP7_75t_L g826 ( .A(n_603), .Y(n_826) );
OA211x2_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B(n_608), .C(n_611), .Y(n_604) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g673 ( .A(n_607), .Y(n_673) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g771 ( .A(n_612), .Y(n_771) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
INVx1_ASAP7_75t_L g837 ( .A(n_616), .Y(n_837) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx2_ASAP7_75t_L g647 ( .A(n_620), .Y(n_647) );
BUFx4f_ASAP7_75t_SL g668 ( .A(n_620), .Y(n_668) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
XOR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_654), .Y(n_626) );
NAND3x1_ASAP7_75t_L g627 ( .A(n_628), .B(n_642), .C(n_648), .Y(n_627) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_629), .B(n_635), .Y(n_628) );
OAI21xp5_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_631), .B(n_632), .Y(n_629) );
BUFx2_ASAP7_75t_L g675 ( .A(n_630), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g901 ( .A1(n_630), .A2(n_902), .B(n_903), .Y(n_901) );
OAI21xp5_ASAP7_75t_SL g926 ( .A1(n_630), .A2(n_927), .B(n_928), .Y(n_926) );
OAI21xp5_ASAP7_75t_L g967 ( .A1(n_630), .A2(n_968), .B(n_969), .Y(n_967) );
INVx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .C(n_639), .Y(n_635) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .Y(n_648) );
BUFx2_ASAP7_75t_L g993 ( .A(n_650), .Y(n_993) );
INVx1_ASAP7_75t_L g689 ( .A(n_656), .Y(n_689) );
INVx1_ASAP7_75t_SL g688 ( .A(n_657), .Y(n_688) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_658), .B(n_669), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_674), .C(n_683), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_673), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_677), .B2(n_679), .C(n_680), .Y(n_674) );
OAI21xp5_ASAP7_75t_SL g1013 ( .A1(n_675), .A2(n_1014), .B(n_1015), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
INVxp67_ASAP7_75t_L g868 ( .A(n_681), .Y(n_868) );
BUFx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx3_ASAP7_75t_L g708 ( .A(n_682), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_686), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
XOR2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_751), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_728), .B2(n_750), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g727 ( .A(n_696), .Y(n_727) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_714), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_702), .C(n_710), .Y(n_697) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_720), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_721), .B(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g750 ( .A(n_728), .Y(n_750) );
NOR4xp75_ASAP7_75t_L g729 ( .A(n_730), .B(n_735), .C(n_740), .D(n_745), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_731), .B(n_733), .Y(n_730) );
INVx2_ASAP7_75t_L g830 ( .A(n_732), .Y(n_830) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_734), .Y(n_851) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_736), .B(n_738), .Y(n_735) );
BUFx2_ASAP7_75t_L g854 ( .A(n_739), .Y(n_854) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_741), .B(n_744), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g745 ( .A1(n_746), .A2(n_748), .B(n_749), .Y(n_745) );
OAI21xp33_ASAP7_75t_SL g817 ( .A1(n_746), .A2(n_818), .B(n_819), .Y(n_817) );
OAI21xp33_ASAP7_75t_L g947 ( .A1(n_746), .A2(n_948), .B(n_949), .Y(n_947) );
INVx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_782), .B2(n_783), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
BUFx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g781 ( .A(n_757), .Y(n_781) );
NAND3x1_ASAP7_75t_L g757 ( .A(n_758), .B(n_772), .C(n_777), .Y(n_757) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_759), .B(n_763), .Y(n_758) );
OAI21xp5_ASAP7_75t_SL g759 ( .A1(n_760), .A2(n_761), .B(n_762), .Y(n_759) );
OAI21xp5_ASAP7_75t_SL g984 ( .A1(n_760), .A2(n_985), .B(n_986), .Y(n_984) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .C(n_767), .Y(n_763) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g934 ( .A(n_769), .Y(n_934) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g772 ( .A(n_773), .B(n_775), .Y(n_772) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_780), .Y(n_777) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g797 ( .A(n_784), .Y(n_797) );
NAND5xp2_ASAP7_75t_SL g785 ( .A(n_786), .B(n_788), .C(n_790), .D(n_793), .E(n_796), .Y(n_785) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_789), .Y(n_1084) );
AND2x2_ASAP7_75t_SL g790 ( .A(n_791), .B(n_792), .Y(n_790) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g1048 ( .A(n_799), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_802), .B1(n_939), .B2(n_1046), .Y(n_799) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
XNOR2xp5_ASAP7_75t_SL g802 ( .A(n_803), .B(n_872), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_805), .B1(n_839), .B2(n_840), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_823), .Y(n_809) );
NOR3xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_817), .C(n_820), .Y(n_810) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OAI221xp5_ASAP7_75t_SL g858 ( .A1(n_814), .A2(n_859), .B1(n_860), .B2(n_862), .C(n_863), .Y(n_858) );
NOR3xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_828), .C(n_835), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_827), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_828) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g845 ( .A(n_833), .Y(n_845) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g871 ( .A(n_842), .Y(n_871) );
AND2x2_ASAP7_75t_SL g842 ( .A(n_843), .B(n_857), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_844), .B(n_852), .Y(n_843) );
OAI221xp5_ASAP7_75t_SL g844 ( .A1(n_845), .A2(n_846), .B1(n_847), .B2(n_849), .C(n_850), .Y(n_844) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_855), .Y(n_852) );
NOR2xp33_ASAP7_75t_SL g857 ( .A(n_858), .B(n_865), .Y(n_857) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_893), .B1(n_937), .B2(n_938), .Y(n_872) );
INVx2_ASAP7_75t_SL g937 ( .A(n_873), .Y(n_937) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AND3x1_ASAP7_75t_L g876 ( .A(n_877), .B(n_887), .C(n_890), .Y(n_876) );
NOR3xp33_ASAP7_75t_L g877 ( .A(n_878), .B(n_881), .C(n_884), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
AND2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
AND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g938 ( .A(n_893), .Y(n_938) );
OA22x2_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_895), .B1(n_912), .B2(n_936), .Y(n_893) );
INVx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
XOR2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_911), .Y(n_895) );
NAND3x1_ASAP7_75t_SL g896 ( .A(n_897), .B(n_900), .C(n_908), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
NOR2x1_ASAP7_75t_L g900 ( .A(n_901), .B(n_904), .Y(n_900) );
NAND3xp33_ASAP7_75t_L g904 ( .A(n_905), .B(n_906), .C(n_907), .Y(n_904) );
AND2x2_ASAP7_75t_L g908 ( .A(n_909), .B(n_910), .Y(n_908) );
INVx1_ASAP7_75t_L g936 ( .A(n_912), .Y(n_936) );
XOR2x2_ASAP7_75t_L g912 ( .A(n_913), .B(n_935), .Y(n_912) );
AND2x2_ASAP7_75t_SL g913 ( .A(n_914), .B(n_925), .Y(n_913) );
NOR3xp33_ASAP7_75t_L g914 ( .A(n_915), .B(n_919), .C(n_922), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_916), .B(n_918), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_926), .B(n_929), .Y(n_925) );
NAND3xp33_ASAP7_75t_L g929 ( .A(n_930), .B(n_932), .C(n_933), .Y(n_929) );
INVx1_ASAP7_75t_L g1046 ( .A(n_939), .Y(n_1046) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_979), .B1(n_1044), .B2(n_1045), .Y(n_939) );
INVx2_ASAP7_75t_L g1044 ( .A(n_940), .Y(n_1044) );
XOR2x2_ASAP7_75t_L g940 ( .A(n_941), .B(n_961), .Y(n_940) );
AND2x2_ASAP7_75t_L g942 ( .A(n_943), .B(n_953), .Y(n_942) );
NOR3xp33_ASAP7_75t_L g943 ( .A(n_944), .B(n_947), .C(n_950), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_958), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_957), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .Y(n_958) );
INVx2_ASAP7_75t_L g1028 ( .A(n_961), .Y(n_1028) );
XOR2x2_ASAP7_75t_L g961 ( .A(n_962), .B(n_978), .Y(n_961) );
NAND3x1_ASAP7_75t_L g962 ( .A(n_963), .B(n_966), .C(n_974), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_964), .B(n_965), .Y(n_963) );
NOR2x1_ASAP7_75t_L g966 ( .A(n_967), .B(n_970), .Y(n_966) );
NAND3xp33_ASAP7_75t_L g970 ( .A(n_971), .B(n_972), .C(n_973), .Y(n_970) );
AND2x2_ASAP7_75t_L g974 ( .A(n_975), .B(n_977), .Y(n_974) );
INVx1_ASAP7_75t_L g1045 ( .A(n_979), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_1026), .B1(n_1042), .B2(n_1043), .Y(n_979) );
INVx1_ASAP7_75t_L g1042 ( .A(n_980), .Y(n_1042) );
AOI22xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_1003), .B1(n_1004), .B2(n_1025), .Y(n_980) );
INVx1_ASAP7_75t_L g1025 ( .A(n_981), .Y(n_1025) );
NAND3x1_ASAP7_75t_L g982 ( .A(n_983), .B(n_991), .C(n_995), .Y(n_982) );
NOR2xp33_ASAP7_75t_L g983 ( .A(n_984), .B(n_988), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_989), .B(n_990), .Y(n_988) );
AND2x2_ASAP7_75t_L g991 ( .A(n_992), .B(n_994), .Y(n_991) );
OAI21xp33_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_998), .B(n_1000), .Y(n_996) );
BUFx2_ASAP7_75t_R g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1024 ( .A(n_1007), .Y(n_1024) );
NAND2x1p5_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1016), .Y(n_1007) );
NOR2xp67_ASAP7_75t_SL g1008 ( .A(n_1009), .B(n_1013), .Y(n_1008) );
NAND3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .C(n_1012), .Y(n_1009) );
NOR2x1_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1020), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1023), .Y(n_1020) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1026), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g1026 ( .A1(n_1027), .A2(n_1028), .B1(n_1029), .B2(n_1041), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1029), .Y(n_1041) );
NAND4xp75_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1034), .C(n_1037), .D(n_1040), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
AND2x2_ASAP7_75t_SL g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
INVx1_ASAP7_75t_SL g1049 ( .A(n_1050), .Y(n_1049) );
NOR2x1_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1055), .Y(n_1050) );
OR2x2_ASAP7_75t_SL g1102 ( .A(n_1051), .B(n_1056), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1054), .Y(n_1051) );
CKINVDCx20_ASAP7_75t_R g1091 ( .A(n_1052), .Y(n_1091) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_1053), .B(n_1094), .Y(n_1097) );
CKINVDCx16_ASAP7_75t_R g1094 ( .A(n_1054), .Y(n_1094) );
CKINVDCx20_ASAP7_75t_R g1055 ( .A(n_1056), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1058), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1061), .Y(n_1059) );
OAI322xp33_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1090), .A3(n_1092), .B1(n_1095), .B2(n_1098), .C1(n_1099), .C2(n_1100), .Y(n_1062) );
INVx2_ASAP7_75t_SL g1089 ( .A(n_1064), .Y(n_1089) );
AND2x4_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1076), .Y(n_1064) );
NOR3xp33_ASAP7_75t_SL g1065 ( .A(n_1066), .B(n_1070), .C(n_1073), .Y(n_1065) );
NOR2x1_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1082), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1081), .Y(n_1077) );
INVx2_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1085), .Y(n_1082) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
CKINVDCx16_ASAP7_75t_R g1095 ( .A(n_1096), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_1101), .Y(n_1100) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_1102), .Y(n_1101) );
endmodule