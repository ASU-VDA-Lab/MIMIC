module fake_jpeg_24459_n_348 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_20),
.B1(n_16),
.B2(n_23),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_21),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_58),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_68),
.B1(n_29),
.B2(n_24),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_20),
.B1(n_16),
.B2(n_23),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_67),
.B1(n_70),
.B2(n_76),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_50),
.B1(n_46),
.B2(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_64),
.B1(n_72),
.B2(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_69),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_16),
.B1(n_23),
.B2(n_32),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_17),
.B1(n_19),
.B2(n_32),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_13),
.B(n_14),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_25),
.B1(n_19),
.B2(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_73),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_17),
.B1(n_27),
.B2(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_35),
.B1(n_33),
.B2(n_31),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_37),
.A2(n_35),
.B1(n_33),
.B2(n_31),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_47),
.B1(n_45),
.B2(n_31),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_87),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_85),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_86),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_91),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_90),
.A2(n_121),
.B1(n_57),
.B2(n_66),
.Y(n_145)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_92),
.B(n_111),
.Y(n_130)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_33),
.B1(n_29),
.B2(n_24),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_110),
.B1(n_59),
.B2(n_77),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_115),
.B(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_103),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_29),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_63),
.Y(n_109)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_24),
.B1(n_18),
.B2(n_14),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_74),
.B(n_14),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_13),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_116),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_65),
.A2(n_12),
.B1(n_11),
.B2(n_18),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_12),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_63),
.B(n_81),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_61),
.B(n_73),
.Y(n_128)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_0),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_54),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_127),
.B1(n_133),
.B2(n_103),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_63),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_137),
.B(n_151),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_79),
.B1(n_66),
.B2(n_57),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_132),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_75),
.C(n_64),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_140),
.C(n_152),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_93),
.B1(n_102),
.B2(n_90),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_72),
.B(n_75),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_78),
.C(n_66),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_147),
.B1(n_97),
.B2(n_91),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_95),
.A2(n_57),
.B1(n_56),
.B2(n_3),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_93),
.A2(n_1),
.B(n_2),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_1),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_153),
.B(n_157),
.Y(n_219)
);

AO21x2_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_93),
.B(n_121),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_154),
.A2(n_164),
.B(n_148),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_104),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_159),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_158),
.B1(n_168),
.B2(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_83),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_120),
.B1(n_104),
.B2(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_117),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_150),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_107),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_96),
.B(n_87),
.C(n_118),
.Y(n_164)
);

BUFx24_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

XOR2x2_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_89),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_166),
.B(n_6),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_169),
.B1(n_175),
.B2(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_114),
.B1(n_84),
.B2(n_109),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_108),
.B1(n_86),
.B2(n_85),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_176),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_11),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_180),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_3),
.B(n_4),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_151),
.B(n_128),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_113),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_122),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_177),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_123),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_178),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_130),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_181),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_4),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_132),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_135),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_148),
.B(n_131),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_5),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_129),
.B(n_105),
.C(n_7),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_149),
.C(n_129),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_188),
.B(n_203),
.C(n_216),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_193),
.A2(n_214),
.B1(n_217),
.B2(n_218),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_151),
.B(n_124),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_207),
.B(n_221),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_199),
.A2(n_175),
.B(n_165),
.Y(n_241)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_154),
.A2(n_166),
.B1(n_174),
.B2(n_172),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_205),
.B(n_170),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_124),
.B1(n_126),
.B2(n_139),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_204),
.B1(n_201),
.B2(n_195),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_126),
.C(n_139),
.Y(n_203)
);

OAI22x1_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_146),
.B1(n_134),
.B2(n_136),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_164),
.B1(n_165),
.B2(n_169),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_136),
.B(n_130),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_170),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_131),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_203),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_156),
.A2(n_138),
.B1(n_8),
.B2(n_9),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_183),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_138),
.C(n_9),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_154),
.A2(n_8),
.B1(n_10),
.B2(n_158),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_10),
.B1(n_168),
.B2(n_176),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_159),
.A2(n_10),
.A3(n_155),
.B1(n_178),
.B2(n_167),
.C1(n_185),
.C2(n_177),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_220),
.B(n_188),
.CI(n_216),
.CON(n_249),
.SN(n_249)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_174),
.A2(n_10),
.B(n_153),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_193),
.B1(n_205),
.B2(n_199),
.Y(n_251)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_213),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_232),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_206),
.B(n_161),
.Y(n_225)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_206),
.B(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_226),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_162),
.Y(n_227)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_227),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_200),
.C(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_230),
.Y(n_255)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_190),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_238),
.B1(n_243),
.B2(n_246),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_248),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_240),
.B(n_241),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_187),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_165),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_197),
.Y(n_253)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_200),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_194),
.C(n_196),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_254),
.C(n_259),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_251),
.A2(n_261),
.B1(n_247),
.B2(n_239),
.Y(n_288)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_212),
.C(n_215),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_247),
.A2(n_205),
.B1(n_195),
.B2(n_192),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_257),
.A2(n_230),
.B1(n_246),
.B2(n_236),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_198),
.C(n_209),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_267),
.C(n_272),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_235),
.B1(n_222),
.B2(n_244),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_248),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_237),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_194),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_249),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_196),
.C(n_231),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_273),
.A2(n_282),
.B(n_286),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_254),
.C(n_260),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_224),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_278),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_241),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_229),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_280),
.B(n_281),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_255),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_234),
.Y(n_283)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_287),
.B1(n_291),
.B2(n_252),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_258),
.B1(n_257),
.B2(n_242),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_269),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_290),
.B(n_249),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_239),
.B(n_238),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_251),
.B1(n_223),
.B2(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_296),
.A2(n_297),
.B1(n_303),
.B2(n_304),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_272),
.B1(n_242),
.B2(n_259),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_305),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_301),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_264),
.B1(n_267),
.B2(n_262),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_285),
.C(n_275),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_279),
.C(n_285),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_320),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_302),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_311),
.B(n_318),
.Y(n_329)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_296),
.A2(n_291),
.B(n_289),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_304),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_297),
.C(n_299),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_300),
.B1(n_298),
.B2(n_294),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_289),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_317),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_312),
.B(n_313),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_303),
.B1(n_294),
.B2(n_301),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_324),
.B(n_325),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_262),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_278),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_305),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_318),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_331),
.B(n_335),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_336),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_310),
.C(n_316),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_313),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_SL g340 ( 
.A(n_331),
.B(n_322),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_332),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_335),
.C(n_326),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_342),
.B(n_343),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_339),
.C(n_330),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_334),
.B(n_338),
.Y(n_346)
);

AOI32xp33_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_321),
.A3(n_319),
.B1(n_333),
.B2(n_315),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_347),
.B(n_315),
.Y(n_348)
);


endmodule