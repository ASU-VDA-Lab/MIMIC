module real_jpeg_27983_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_0),
.A2(n_42),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_1),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_2),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_73)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_5),
.A2(n_18),
.B1(n_19),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_5),
.A2(n_31),
.B1(n_42),
.B2(n_45),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_69)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_6),
.A2(n_18),
.B(n_20),
.C(n_21),
.D(n_29),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_18),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_6),
.B(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_25),
.Y(n_81)
);

A2O1A1O1Ixp25_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_25),
.B(n_37),
.C(n_81),
.D(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_6),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_6),
.A2(n_58),
.B(n_74),
.Y(n_103)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_10),
.A2(n_36),
.B1(n_42),
.B2(n_45),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_77),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_76),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_64),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_15),
.B(n_64),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_48),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_33),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_19),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI32xp33_ASAP7_75t_L g61 ( 
.A1(n_19),
.A2(n_20),
.A3(n_25),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_24),
.B(n_28),
.Y(n_63)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_24),
.A2(n_39),
.A3(n_45),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_38),
.B(n_40),
.C(n_41),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_38),
.Y(n_40)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_41),
.B2(n_46),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_66),
.B(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_38),
.B(n_42),
.Y(n_82)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_59),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_45),
.B(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_61),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_57),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_53),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_92),
.B(n_101),
.Y(n_100)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_75),
.Y(n_74)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_99),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_70),
.C(n_72),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_88),
.B(n_108),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_79),
.B(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_83),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_96),
.B(n_107),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_95),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_102),
.B(n_106),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);


endmodule