module fake_jpeg_5138_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_23),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_17),
.B1(n_16),
.B2(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_53),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_16),
.B1(n_31),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_55),
.B1(n_26),
.B2(n_23),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_61),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_32),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_36),
.B1(n_39),
.B2(n_28),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_34),
.B1(n_42),
.B2(n_40),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_73),
.B1(n_63),
.B2(n_24),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_42),
.B1(n_34),
.B2(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_80),
.B1(n_59),
.B2(n_49),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_35),
.C(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_26),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_42),
.B1(n_32),
.B2(n_36),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_102),
.B1(n_103),
.B2(n_20),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_90),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_97),
.B1(n_67),
.B2(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_56),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_69),
.B(n_54),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_51),
.B1(n_59),
.B2(n_52),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_76),
.B1(n_73),
.B2(n_66),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_114),
.B1(n_116),
.B2(n_120),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_90),
.B1(n_98),
.B2(n_92),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_74),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.C(n_117),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_68),
.C(n_74),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_70),
.B(n_78),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_33),
.B(n_30),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_36),
.B1(n_72),
.B2(n_78),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_53),
.B1(n_44),
.B2(n_72),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_102),
.C(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_52),
.B1(n_20),
.B2(n_29),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_0),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_47),
.B1(n_15),
.B2(n_52),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_47),
.B1(n_33),
.B2(n_19),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_47),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_136),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_130),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_95),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_132),
.C(n_144),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_123),
.B1(n_110),
.B2(n_109),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_30),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_93),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_135),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_1),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_139),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_27),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_138),
.A2(n_143),
.B(n_124),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_91),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_27),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_145),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_113),
.B(n_111),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_27),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_27),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_143),
.A2(n_112),
.B(n_116),
.C(n_114),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_141),
.B1(n_144),
.B2(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_159),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_111),
.A3(n_120),
.B1(n_109),
.B2(n_122),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_132),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_110),
.C(n_108),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_1),
.C(n_2),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_162),
.B1(n_1),
.B2(n_2),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_134),
.B(n_128),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_28),
.B1(n_27),
.B2(n_6),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_130),
.B(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_171),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_152),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_172),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_150),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_168),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_138),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_174),
.C(n_179),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_146),
.B1(n_148),
.B2(n_159),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_14),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_185),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_178),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_162),
.B1(n_154),
.B2(n_146),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_149),
.C(n_163),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_188),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_163),
.C(n_151),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_146),
.C(n_156),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_182),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_174),
.B(n_176),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_170),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_194),
.B(n_195),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_171),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_200),
.B(n_198),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_165),
.B1(n_179),
.B2(n_10),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_180),
.B1(n_9),
.B2(n_11),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_8),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_205),
.B(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_186),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_187),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_194),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_180),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_209),
.C(n_210),
.Y(n_216)
);

NOR4xp25_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_184),
.C(n_9),
.D(n_11),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_184),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_201),
.C(n_202),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_214),
.B(n_215),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_8),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_9),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_11),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_220),
.Y(n_222)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_14),
.B(n_12),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_12),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_218),
.A2(n_211),
.B(n_13),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_223),
.C(n_12),
.Y(n_225)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_225),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_224),
.Y(n_227)
);


endmodule