module fake_jpeg_15571_n_81 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_81);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_81;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx6_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_7),
.B(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_29),
.Y(n_33)
);

NOR2xp67_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_27),
.B(n_8),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_2),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_20),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_39),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_39),
.B(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_12),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_20),
.B1(n_17),
.B2(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_30),
.B1(n_23),
.B2(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_23),
.A2(n_17),
.B1(n_22),
.B2(n_18),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_24),
.A2(n_29),
.B1(n_25),
.B2(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_47),
.B1(n_3),
.B2(n_6),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_18),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_3),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_24),
.A2(n_18),
.B1(n_5),
.B2(n_6),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_10),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_25),
.B(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_58),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_38),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_9),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_3),
.B1(n_7),
.B2(n_10),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_37),
.B1(n_45),
.B2(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_61),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_46),
.C(n_41),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_53),
.C(n_55),
.Y(n_72)
);

XOR2x2_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_44),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_51),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_70),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_73),
.B(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_55),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_40),
.B1(n_35),
.B2(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_65),
.B1(n_64),
.B2(n_66),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

AOI321xp33_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_76),
.A3(n_74),
.B1(n_78),
.B2(n_57),
.C(n_42),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_57),
.B(n_61),
.Y(n_81)
);


endmodule