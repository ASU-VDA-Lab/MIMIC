module fake_ariane_2870_n_857 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_857);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_857;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_818;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_721;
wire n_600;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_260;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_809;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_755;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_767;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_106),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_33),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_124),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_116),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_120),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_18),
.B(n_100),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_25),
.Y(n_205)
);

BUFx2_ASAP7_75t_SL g206 ( 
.A(n_189),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_64),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_11),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_81),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_69),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_39),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_86),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_101),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_99),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_102),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_53),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_59),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_142),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_32),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_123),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_78),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_4),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_117),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_149),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_96),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_132),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_55),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_5),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_4),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_85),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_6),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_89),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_80),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_35),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_178),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_68),
.Y(n_240)
);

CKINVDCx11_ASAP7_75t_R g241 ( 
.A(n_60),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_6),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_166),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_40),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_146),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_159),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_76),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_136),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_122),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_87),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_168),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_51),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_155),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_148),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_88),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_143),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_108),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_115),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_46),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_62),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_154),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_54),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_3),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_147),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_204),
.B(n_0),
.Y(n_266)
);

OAI22x1_ASAP7_75t_R g267 ( 
.A1(n_235),
.A2(n_242),
.B1(n_201),
.B2(n_225),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_215),
.B(n_1),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_17),
.Y(n_272)
);

OA21x2_ASAP7_75t_L g273 ( 
.A1(n_209),
.A2(n_1),
.B(n_2),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_210),
.A2(n_224),
.B(n_211),
.Y(n_276)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_222),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_229),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_241),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

NOR2x1_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_19),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_220),
.A2(n_95),
.B(n_191),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_198),
.Y(n_294)
);

NOR2x1_ASAP7_75t_L g295 ( 
.A(n_238),
.B(n_20),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_193),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_246),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_7),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_200),
.B(n_7),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_245),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_205),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_212),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_195),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_306)
);

BUFx12f_ASAP7_75t_L g307 ( 
.A(n_207),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_251),
.B(n_8),
.Y(n_309)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_257),
.A2(n_9),
.B(n_10),
.Y(n_313)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_206),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_297),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_282),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_275),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_282),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_314),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_278),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_278),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_R g324 ( 
.A(n_286),
.B(n_194),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_308),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_309),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_307),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_271),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_267),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_271),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_314),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_311),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_300),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_314),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_300),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_270),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_311),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_299),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_291),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_280),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_291),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_303),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_292),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_303),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_285),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_303),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_289),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_296),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_255),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_292),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_292),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_292),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_296),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_287),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_294),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_312),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_294),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_277),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

NOR3xp33_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_306),
.C(n_281),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_347),
.B(n_266),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_302),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_318),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_294),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_324),
.B(n_315),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

NOR3xp33_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_295),
.C(n_265),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_321),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_294),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_332),
.B(n_315),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_319),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_322),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_366),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_327),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_340),
.B(n_304),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_336),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_334),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_339),
.B(n_315),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_276),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_352),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_343),
.B(n_304),
.Y(n_396)
);

BUFx6f_ASAP7_75t_SL g397 ( 
.A(n_339),
.Y(n_397)
);

NAND3xp33_ASAP7_75t_L g398 ( 
.A(n_334),
.B(n_276),
.C(n_273),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_304),
.Y(n_399)
);

AND2x6_ASAP7_75t_L g400 ( 
.A(n_351),
.B(n_272),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_341),
.B(n_361),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_341),
.B(n_255),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_320),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_362),
.B(n_196),
.Y(n_405)
);

XOR2x2_ASAP7_75t_L g406 ( 
.A(n_335),
.B(n_288),
.Y(n_406)
);

A2O1A1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_345),
.A2(n_290),
.B(n_284),
.C(n_293),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_355),
.A2(n_276),
.B(n_283),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_313),
.C(n_273),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_358),
.B(n_269),
.Y(n_410)
);

NOR3xp33_ASAP7_75t_L g411 ( 
.A(n_348),
.B(n_269),
.C(n_203),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_350),
.B(n_304),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_365),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_326),
.B(n_197),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_346),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_364),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_354),
.B(n_305),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g418 ( 
.A1(n_328),
.A2(n_313),
.B1(n_273),
.B2(n_305),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_327),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_323),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_356),
.B(n_310),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_331),
.B(n_199),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_357),
.B(n_310),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_327),
.B(n_305),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_342),
.B(n_202),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_333),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_333),
.B(n_305),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_333),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_333),
.B(n_283),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_345),
.B(n_310),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_345),
.B(n_277),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_347),
.B(n_277),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_345),
.B(n_277),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_373),
.A2(n_313),
.B1(n_301),
.B2(n_298),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_213),
.Y(n_437)
);

NOR2x1p5_ASAP7_75t_L g438 ( 
.A(n_375),
.B(n_214),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_386),
.B(n_284),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_391),
.B(n_216),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_385),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_293),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_374),
.B(n_217),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_404),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_219),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_386),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_379),
.A2(n_243),
.B1(n_221),
.B2(n_223),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_394),
.B(n_203),
.Y(n_449)
);

AND2x4_ASAP7_75t_SL g450 ( 
.A(n_415),
.B(n_301),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_430),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_392),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_398),
.A2(n_298),
.B1(n_287),
.B2(n_262),
.Y(n_454)
);

NOR3xp33_ASAP7_75t_SL g455 ( 
.A(n_414),
.B(n_426),
.C(n_423),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_372),
.A2(n_249),
.B1(n_260),
.B2(n_259),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_226),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_397),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_369),
.B(n_228),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_410),
.B(n_11),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_380),
.B(n_230),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_SL g464 ( 
.A(n_371),
.B(n_256),
.C(n_237),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_397),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_388),
.B(n_411),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_402),
.B(n_287),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_389),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_384),
.Y(n_470)
);

NAND3xp33_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_254),
.C(n_252),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_370),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_406),
.A2(n_239),
.B1(n_236),
.B2(n_14),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_401),
.B(n_12),
.Y(n_474)
);

NAND2x1p5_ASAP7_75t_L g475 ( 
.A(n_413),
.B(n_287),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_435),
.B(n_12),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_393),
.B(n_13),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_398),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_377),
.B(n_15),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_432),
.B(n_16),
.Y(n_481)
);

INVx5_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_416),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_434),
.B(n_16),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_425),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_419),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_403),
.B(n_21),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_399),
.B(n_22),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_407),
.A2(n_23),
.B(n_24),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_408),
.A2(n_26),
.B(n_27),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_376),
.B(n_192),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_428),
.Y(n_493)
);

NOR2xp67_ASAP7_75t_L g494 ( 
.A(n_412),
.B(n_28),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_405),
.B(n_190),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_418),
.A2(n_409),
.B1(n_394),
.B2(n_400),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_382),
.B(n_29),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_429),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_417),
.B(n_30),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_409),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_422),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_381),
.B(n_37),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_419),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_400),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_453),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_441),
.Y(n_507)
);

AOI222xp33_ASAP7_75t_L g508 ( 
.A1(n_473),
.A2(n_396),
.B1(n_390),
.B2(n_427),
.C1(n_43),
.C2(n_44),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_449),
.A2(n_427),
.B(n_41),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_447),
.B(n_439),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_444),
.A2(n_427),
.B(n_42),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_SL g513 ( 
.A(n_455),
.B(n_38),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_457),
.B(n_45),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_47),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_469),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_48),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_487),
.B(n_49),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_446),
.A2(n_50),
.B(n_52),
.Y(n_519)
);

A2O1A1Ixp33_ASAP7_75t_SL g520 ( 
.A1(n_489),
.A2(n_188),
.B(n_57),
.C(n_58),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_474),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_491),
.A2(n_56),
.B(n_61),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_437),
.A2(n_485),
.B(n_488),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_442),
.B(n_63),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_462),
.A2(n_65),
.B(n_66),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_482),
.B(n_67),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_490),
.A2(n_70),
.B(n_71),
.Y(n_528)
);

OAI21xp33_ASAP7_75t_L g529 ( 
.A1(n_476),
.A2(n_72),
.B(n_73),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_460),
.B(n_74),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_450),
.Y(n_531)
);

NOR2x1_ASAP7_75t_R g532 ( 
.A(n_458),
.B(n_75),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_482),
.B(n_77),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_465),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_474),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_497),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

OAI21xp33_ASAP7_75t_L g538 ( 
.A1(n_478),
.A2(n_84),
.B(n_90),
.Y(n_538)
);

O2A1O1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_461),
.A2(n_91),
.B(n_92),
.C(n_93),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_482),
.B(n_94),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_466),
.B(n_97),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_493),
.A2(n_98),
.B(n_103),
.Y(n_542)
);

O2A1O1Ixp33_ASAP7_75t_L g543 ( 
.A1(n_477),
.A2(n_104),
.B(n_105),
.C(n_107),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_472),
.B(n_464),
.Y(n_544)
);

O2A1O1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_440),
.A2(n_109),
.B(n_110),
.C(n_111),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_438),
.B(n_112),
.Y(n_547)
);

BUFx6f_ASAP7_75t_SL g548 ( 
.A(n_505),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_469),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_492),
.B(n_113),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_448),
.B(n_185),
.Y(n_551)
);

OA22x2_ASAP7_75t_L g552 ( 
.A1(n_452),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_449),
.B(n_125),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_484),
.B(n_126),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_454),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_499),
.A2(n_131),
.B(n_133),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_470),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_436),
.A2(n_134),
.B(n_135),
.Y(n_558)
);

AO21x1_ASAP7_75t_L g559 ( 
.A1(n_495),
.A2(n_137),
.B(n_138),
.Y(n_559)
);

AOI21xp33_ASAP7_75t_L g560 ( 
.A1(n_479),
.A2(n_139),
.B(n_140),
.Y(n_560)
);

O2A1O1Ixp33_ASAP7_75t_L g561 ( 
.A1(n_480),
.A2(n_141),
.B(n_144),
.C(n_150),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_481),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_503),
.B(n_151),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_501),
.A2(n_152),
.B(n_153),
.Y(n_564)
);

BUFx4_ASAP7_75t_R g565 ( 
.A(n_534),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g566 ( 
.A1(n_528),
.A2(n_500),
.B(n_498),
.Y(n_566)
);

AO21x2_ASAP7_75t_L g567 ( 
.A1(n_524),
.A2(n_494),
.B(n_503),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_558),
.A2(n_502),
.B(n_504),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_546),
.Y(n_569)
);

AOI22x1_ASAP7_75t_L g570 ( 
.A1(n_511),
.A2(n_475),
.B1(n_467),
.B2(n_486),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_514),
.A2(n_449),
.B(n_562),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_507),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_537),
.Y(n_573)
);

BUFx8_ASAP7_75t_L g574 ( 
.A(n_548),
.Y(n_574)
);

BUFx4f_ASAP7_75t_SL g575 ( 
.A(n_506),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_523),
.A2(n_459),
.B(n_471),
.Y(n_576)
);

OAI21x1_ASAP7_75t_L g577 ( 
.A1(n_509),
.A2(n_449),
.B(n_456),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_557),
.Y(n_578)
);

AOI22x1_ASAP7_75t_L g579 ( 
.A1(n_519),
.A2(n_496),
.B1(n_486),
.B2(n_468),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_522),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_521),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_512),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_510),
.Y(n_583)
);

BUFx12f_ASAP7_75t_L g584 ( 
.A(n_535),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_515),
.Y(n_585)
);

AO21x2_ASAP7_75t_L g586 ( 
.A1(n_530),
.A2(n_496),
.B(n_486),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_546),
.Y(n_587)
);

BUFx8_ASAP7_75t_SL g588 ( 
.A(n_548),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_516),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_531),
.Y(n_590)
);

OA21x2_ASAP7_75t_L g591 ( 
.A1(n_538),
.A2(n_496),
.B(n_468),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_544),
.B(n_468),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_553),
.A2(n_463),
.B(n_157),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_552),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_541),
.A2(n_538),
.B(n_518),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_516),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_549),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_508),
.B(n_463),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_549),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_525),
.A2(n_156),
.B(n_160),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_542),
.A2(n_526),
.B(n_550),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_547),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_554),
.Y(n_603)
);

AOI22x1_ASAP7_75t_L g604 ( 
.A1(n_556),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_513),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_517),
.B(n_165),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_564),
.A2(n_167),
.B(n_170),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_564),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_536),
.Y(n_609)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_555),
.A2(n_172),
.B(n_173),
.Y(n_610)
);

NOR2x1_ASAP7_75t_R g611 ( 
.A(n_532),
.B(n_174),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_563),
.Y(n_612)
);

INVx6_ASAP7_75t_L g613 ( 
.A(n_532),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_578),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_582),
.B(n_551),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_572),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_594),
.B(n_527),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_573),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_578),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_580),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_612),
.B(n_540),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_575),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_565),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_612),
.A2(n_559),
.B1(n_529),
.B2(n_539),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_568),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_569),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_595),
.A2(n_533),
.B(n_520),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_591),
.A2(n_560),
.B(n_545),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_589),
.Y(n_629)
);

BUFx4f_ASAP7_75t_SL g630 ( 
.A(n_574),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_598),
.B(n_561),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_591),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_591),
.Y(n_634)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_574),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_581),
.B(n_543),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_575),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_609),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_607),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_609),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_581),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_574),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_583),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_592),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_602),
.A2(n_183),
.B1(n_184),
.B2(n_585),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_592),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_592),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_569),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_607),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_613),
.B(n_565),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_613),
.B(n_602),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_569),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_586),
.Y(n_653)
);

AOI21x1_ASAP7_75t_L g654 ( 
.A1(n_571),
.A2(n_601),
.B(n_576),
.Y(n_654)
);

INVx6_ASAP7_75t_L g655 ( 
.A(n_569),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_584),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_584),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_616),
.Y(n_658)
);

CKINVDCx12_ASAP7_75t_R g659 ( 
.A(n_630),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_623),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_618),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_623),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_629),
.B(n_586),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_635),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_657),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_623),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_619),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_R g668 ( 
.A(n_650),
.B(n_605),
.Y(n_668)
);

NOR3xp33_ASAP7_75t_SL g669 ( 
.A(n_615),
.B(n_605),
.C(n_613),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_R g670 ( 
.A(n_635),
.B(n_587),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_620),
.Y(n_671)
);

NAND2x1p5_ASAP7_75t_L g672 ( 
.A(n_648),
.B(n_596),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_641),
.Y(n_673)
);

NOR3xp33_ASAP7_75t_SL g674 ( 
.A(n_651),
.B(n_611),
.C(n_588),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_622),
.B(n_588),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_643),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_629),
.B(n_577),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_632),
.A2(n_606),
.B1(n_603),
.B2(n_590),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_614),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_626),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_614),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_648),
.B(n_596),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_626),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_631),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_648),
.B(n_599),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_631),
.B(n_577),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_632),
.B(n_608),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_644),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_656),
.B(n_617),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_646),
.B(n_603),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_626),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_642),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_657),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_617),
.B(n_597),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_647),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_626),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_624),
.A2(n_606),
.B1(n_597),
.B2(n_599),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_652),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_652),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_621),
.B(n_608),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_621),
.B(n_606),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_636),
.A2(n_603),
.B1(n_590),
.B2(n_567),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_642),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_676),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_687),
.B(n_634),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_658),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_687),
.B(n_634),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_673),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_661),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_698),
.B(n_603),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_701),
.B(n_633),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_677),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_665),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_701),
.B(n_652),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_665),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_681),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_671),
.B(n_637),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_700),
.B(n_652),
.Y(n_719)
);

NAND2x1p5_ASAP7_75t_L g720 ( 
.A(n_682),
.B(n_652),
.Y(n_720)
);

OR2x2_ASAP7_75t_SL g721 ( 
.A(n_693),
.B(n_655),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_702),
.B(n_653),
.Y(n_722)
);

AOI221xp5_ASAP7_75t_L g723 ( 
.A1(n_689),
.A2(n_678),
.B1(n_695),
.B2(n_702),
.C(n_638),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_677),
.B(n_654),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_686),
.B(n_654),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_679),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_688),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_680),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_696),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_686),
.B(n_625),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_683),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_684),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_667),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_682),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_692),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_694),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_713),
.B(n_663),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_705),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_709),
.B(n_694),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_707),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_717),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_711),
.A2(n_669),
.B1(n_645),
.B2(n_640),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_712),
.B(n_690),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_710),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_727),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_706),
.B(n_699),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_729),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_714),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_706),
.B(n_697),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_711),
.A2(n_567),
.B1(n_703),
.B2(n_668),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_718),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_708),
.B(n_712),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_714),
.B(n_691),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_715),
.B(n_704),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_726),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_708),
.B(n_700),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_717),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_732),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_715),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_730),
.B(n_700),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_716),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_755),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_742),
.A2(n_723),
.B1(n_722),
.B2(n_668),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_759),
.B(n_731),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_759),
.B(n_731),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_752),
.B(n_735),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_751),
.B(n_738),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_759),
.B(n_735),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_741),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_749),
.B(n_728),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_756),
.B(n_724),
.Y(n_771)
);

INVx3_ASAP7_75t_SL g772 ( 
.A(n_748),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_748),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_756),
.B(n_715),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_740),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_749),
.B(n_730),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_761),
.B(n_734),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_760),
.B(n_716),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_744),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_762),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_772),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_762),
.B(n_745),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_775),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_779),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_772),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_767),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_766),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_770),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_788),
.B(n_776),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_786),
.A2(n_763),
.B1(n_721),
.B2(n_773),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_781),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_782),
.A2(n_763),
.B(n_777),
.Y(n_792)
);

OAI21xp33_ASAP7_75t_L g793 ( 
.A1(n_780),
.A2(n_777),
.B(n_765),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_791),
.Y(n_794)
);

AOI21xp33_ASAP7_75t_SL g795 ( 
.A1(n_792),
.A2(n_785),
.B(n_664),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_SL g796 ( 
.A1(n_790),
.A2(n_737),
.B1(n_736),
.B2(n_743),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_793),
.B(n_664),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_789),
.A2(n_750),
.B1(n_784),
.B2(n_783),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_789),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_799),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_794),
.Y(n_801)
);

NOR4xp75_ASAP7_75t_L g802 ( 
.A(n_795),
.B(n_782),
.C(n_659),
.D(n_754),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_798),
.B(n_787),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_803),
.A2(n_797),
.B(n_796),
.Y(n_804)
);

NOR2x1_ASAP7_75t_L g805 ( 
.A(n_800),
.B(n_675),
.Y(n_805)
);

AOI211xp5_ASAP7_75t_L g806 ( 
.A1(n_804),
.A2(n_801),
.B(n_802),
.C(n_704),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_805),
.Y(n_807)
);

OAI211xp5_ASAP7_75t_SL g808 ( 
.A1(n_805),
.A2(n_739),
.B(n_674),
.C(n_753),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_807),
.A2(n_806),
.B1(n_808),
.B2(n_764),
.Y(n_809)
);

AND3x4_ASAP7_75t_L g810 ( 
.A(n_806),
.B(n_764),
.C(n_736),
.Y(n_810)
);

NOR2x1_ASAP7_75t_L g811 ( 
.A(n_807),
.B(n_660),
.Y(n_811)
);

AO22x2_ASAP7_75t_SL g812 ( 
.A1(n_807),
.A2(n_670),
.B1(n_778),
.B2(n_768),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_807),
.A2(n_750),
.B1(n_747),
.B2(n_758),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_807),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_814),
.B(n_771),
.Y(n_815)
);

INVx3_ASAP7_75t_SL g816 ( 
.A(n_812),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_813),
.A2(n_809),
.B1(n_810),
.B2(n_811),
.Y(n_817)
);

AND2x2_ASAP7_75t_SL g818 ( 
.A(n_812),
.B(n_670),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_SL g819 ( 
.A1(n_809),
.A2(n_662),
.B(n_666),
.Y(n_819)
);

AND3x2_ASAP7_75t_L g820 ( 
.A(n_814),
.B(n_764),
.C(n_771),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_814),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_821),
.Y(n_822)
);

NOR2x1_ASAP7_75t_L g823 ( 
.A(n_819),
.B(n_587),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_816),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_815),
.B(n_774),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_817),
.A2(n_746),
.B1(n_685),
.B2(n_682),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_818),
.Y(n_827)
);

AOI32xp33_ASAP7_75t_L g828 ( 
.A1(n_820),
.A2(n_685),
.A3(n_746),
.B1(n_760),
.B2(n_566),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_824),
.A2(n_721),
.B1(n_720),
.B2(n_672),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_827),
.A2(n_685),
.B1(n_719),
.B2(n_655),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_822),
.Y(n_831)
);

XOR2xp5_ASAP7_75t_L g832 ( 
.A(n_826),
.B(n_743),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_825),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_823),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_828),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_824),
.A2(n_719),
.B1(n_655),
.B2(n_690),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_824),
.A2(n_720),
.B1(n_672),
.B2(n_734),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_835),
.A2(n_655),
.B1(n_719),
.B2(n_690),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_831),
.B(n_734),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_833),
.B(n_734),
.Y(n_840)
);

AOI31xp33_ASAP7_75t_L g841 ( 
.A1(n_834),
.A2(n_743),
.A3(n_737),
.B(n_725),
.Y(n_841)
);

AOI211xp5_ASAP7_75t_L g842 ( 
.A1(n_837),
.A2(n_610),
.B(n_576),
.C(n_600),
.Y(n_842)
);

OAI31xp33_ASAP7_75t_L g843 ( 
.A1(n_832),
.A2(n_769),
.A3(n_725),
.B(n_724),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_836),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_829),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_830),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_839),
.A2(n_690),
.B1(n_769),
.B2(n_627),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_845),
.Y(n_848)
);

OAI22x1_ASAP7_75t_SL g849 ( 
.A1(n_844),
.A2(n_604),
.B1(n_639),
.B2(n_649),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_840),
.A2(n_627),
.B1(n_570),
.B2(n_579),
.Y(n_850)
);

XOR2xp5_ASAP7_75t_L g851 ( 
.A(n_846),
.B(n_628),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_SL g852 ( 
.A1(n_848),
.A2(n_838),
.B(n_841),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_SL g853 ( 
.A1(n_851),
.A2(n_847),
.B1(n_849),
.B2(n_842),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_852),
.B(n_843),
.C(n_850),
.Y(n_854)
);

AO21x2_ASAP7_75t_L g855 ( 
.A1(n_854),
.A2(n_853),
.B(n_566),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_855),
.B(n_593),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_856),
.A2(n_757),
.B1(n_741),
.B2(n_733),
.Y(n_857)
);


endmodule