module fake_jpeg_31898_n_122 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_122);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_16),
.B(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_34),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_2),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_17),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_22),
.B1(n_11),
.B2(n_12),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_36),
.B1(n_39),
.B2(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_52),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_35),
.B1(n_24),
.B2(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_15),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_46),
.C(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_59),
.B1(n_66),
.B2(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_60),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_69),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_51),
.Y(n_69)
);

OA21x2_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_19),
.B(n_26),
.Y(n_71)
);

AO22x1_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_47),
.B1(n_53),
.B2(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_62),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_77),
.B1(n_85),
.B2(n_81),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_41),
.C(n_56),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_84),
.C(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_71),
.B1(n_72),
.B2(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_27),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_83),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_54),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_19),
.C(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_66),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_65),
.Y(n_98)
);

NOR4xp25_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_95),
.C(n_96),
.D(n_91),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_91),
.B1(n_57),
.B2(n_59),
.Y(n_103)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_71),
.B(n_57),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_64),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_100),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_78),
.C(n_65),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_88),
.B(n_92),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_110),
.B1(n_91),
.B2(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_114),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_98),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_105),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_111),
.C(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_120),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_118),
.C(n_117),
.Y(n_122)
);


endmodule