module real_aes_10574_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_402;
wire n_602;
wire n_552;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_598;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_0), .A2(n_64), .B1(n_128), .B2(n_130), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_1), .B(n_94), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_2), .B(n_59), .Y(n_617) );
AND2x2_ASAP7_75t_L g633 ( .A(n_2), .B(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_2), .Y(n_671) );
INVx1_ASAP7_75t_L g711 ( .A(n_2), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_3), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_4), .Y(n_195) );
INVx2_ASAP7_75t_L g514 ( .A(n_5), .Y(n_514) );
OR2x2_ASAP7_75t_L g546 ( .A(n_5), .B(n_529), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_6), .A2(n_70), .B1(n_598), .B2(n_600), .Y(n_597) );
OAI221xp5_ASAP7_75t_L g653 ( .A1(n_6), .A2(n_70), .B1(n_654), .B2(n_661), .C(n_665), .Y(n_653) );
BUFx2_ASAP7_75t_L g607 ( .A(n_7), .Y(n_607) );
OR2x2_ASAP7_75t_L g616 ( .A(n_7), .B(n_617), .Y(n_616) );
BUFx2_ASAP7_75t_L g620 ( .A(n_7), .Y(n_620) );
INVx1_ASAP7_75t_L g632 ( .A(n_7), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_8), .A2(n_32), .B1(n_108), .B2(n_114), .Y(n_226) );
INVx1_ASAP7_75t_L g497 ( .A(n_9), .Y(n_497) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_10), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_11), .A2(n_47), .B1(n_111), .B2(n_114), .Y(n_110) );
NAND3xp33_ASAP7_75t_L g167 ( .A(n_12), .B(n_114), .C(n_147), .Y(n_167) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_12), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_13), .A2(n_60), .B1(n_575), .B2(n_580), .Y(n_574) );
INVx1_ASAP7_75t_L g676 ( .A(n_13), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_14), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_15), .B(n_161), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_16), .B(n_129), .Y(n_178) );
NAND3xp33_ASAP7_75t_L g162 ( .A(n_17), .B(n_104), .C(n_106), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_18), .A2(n_23), .B1(n_106), .B2(n_108), .Y(n_126) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_19), .A2(n_22), .B1(n_567), .B2(n_569), .C(n_572), .Y(n_566) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_19), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_20), .B(n_161), .Y(n_212) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_21), .Y(n_104) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_22), .Y(n_689) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_24), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_25), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g513 ( .A(n_26), .Y(n_513) );
INVx1_ASAP7_75t_L g529 ( .A(n_26), .Y(n_529) );
INVx1_ASAP7_75t_L g552 ( .A(n_27), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_28), .A2(n_40), .B1(n_111), .B2(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_29), .B(n_104), .Y(n_159) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_29), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_30), .A2(n_537), .B1(n_538), .B2(n_713), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_30), .Y(n_713) );
OAI21x1_ASAP7_75t_L g95 ( .A1(n_31), .A2(n_51), .B(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g118 ( .A(n_33), .B(n_119), .Y(n_118) );
AND2x6_ASAP7_75t_L g99 ( .A(n_34), .B(n_100), .Y(n_99) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_34), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_34), .B(n_506), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_35), .A2(n_67), .B1(n_594), .B2(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g646 ( .A(n_35), .Y(n_646) );
NAND2x1p5_ASAP7_75t_L g168 ( .A(n_36), .B(n_119), .Y(n_168) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_37), .A2(n_63), .B1(n_569), .B2(n_589), .C(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g641 ( .A(n_37), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_38), .B(n_129), .Y(n_214) );
INVx1_ASAP7_75t_L g100 ( .A(n_39), .Y(n_100) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_39), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_41), .B(n_119), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_42), .B(n_106), .Y(n_184) );
INVx1_ASAP7_75t_L g565 ( .A(n_43), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_44), .B(n_106), .Y(n_149) );
NAND2x1_ASAP7_75t_L g219 ( .A(n_45), .B(n_119), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_46), .B(n_147), .Y(n_190) );
INVx2_ASAP7_75t_L g615 ( .A(n_48), .Y(n_615) );
INVx1_ASAP7_75t_L g608 ( .A(n_49), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_50), .B(n_142), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_52), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_53), .B(n_147), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_54), .A2(n_57), .B1(n_106), .B2(n_108), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_55), .Y(n_199) );
BUFx10_ASAP7_75t_L g523 ( .A(n_56), .Y(n_523) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_57), .Y(n_489) );
INVx1_ASAP7_75t_SL g136 ( .A(n_58), .Y(n_136) );
INVx2_ASAP7_75t_L g634 ( .A(n_59), .Y(n_634) );
INVx1_ASAP7_75t_L g692 ( .A(n_60), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_61), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_62), .Y(n_217) );
INVx1_ASAP7_75t_L g635 ( .A(n_63), .Y(n_635) );
INVx2_ASAP7_75t_L g96 ( .A(n_65), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_66), .B(n_147), .Y(n_164) );
INVx1_ASAP7_75t_L g625 ( .A(n_67), .Y(n_625) );
INVx1_ASAP7_75t_L g587 ( .A(n_68), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_69), .B(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_71), .Y(n_501) );
INVx2_ASAP7_75t_L g614 ( .A(n_72), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_73), .B(n_109), .Y(n_146) );
INVx1_ASAP7_75t_L g549 ( .A(n_74), .Y(n_549) );
BUFx3_ASAP7_75t_L g563 ( .A(n_74), .Y(n_563) );
BUFx3_ASAP7_75t_L g521 ( .A(n_75), .Y(n_521) );
INVx1_ASAP7_75t_L g551 ( .A(n_75), .Y(n_551) );
INVx1_ASAP7_75t_L g543 ( .A(n_76), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_477), .B(n_484), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
OR2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_391), .Y(n_82) );
NAND4xp25_ASAP7_75t_L g83 ( .A(n_84), .B(n_302), .C(n_346), .D(n_380), .Y(n_83) );
NOR2xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_258), .Y(n_84) );
OAI221xp5_ASAP7_75t_L g85 ( .A1(n_86), .A2(n_169), .B1(n_202), .B2(n_231), .C(n_239), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_122), .Y(n_87) );
OR2x2_ASAP7_75t_L g371 ( .A(n_88), .B(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_88), .B(n_263), .Y(n_422) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g275 ( .A(n_89), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g234 ( .A(n_90), .Y(n_234) );
INVx1_ASAP7_75t_L g269 ( .A(n_90), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_90), .B(n_124), .Y(n_324) );
INVxp67_ASAP7_75t_SL g356 ( .A(n_90), .Y(n_356) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_90), .Y(n_362) );
OAI21x1_ASAP7_75t_L g90 ( .A1(n_91), .A2(n_101), .B(n_117), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g91 ( .A(n_92), .B(n_97), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
BUFx5_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g135 ( .A(n_94), .Y(n_135) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_94), .Y(n_201) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_L g121 ( .A(n_95), .Y(n_121) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_97), .Y(n_478) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx8_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_98), .A2(n_191), .B(n_201), .Y(n_200) );
INVx8_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g153 ( .A(n_99), .Y(n_153) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_99), .A2(n_158), .B(n_163), .Y(n_157) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_99), .A2(n_177), .B(n_180), .Y(n_176) );
BUFx2_ASAP7_75t_L g218 ( .A(n_99), .Y(n_218) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_101), .A2(n_254), .B(n_255), .Y(n_253) );
OA22x2_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_105), .B1(n_110), .B2(n_115), .Y(n_101) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_102), .A2(n_115), .B1(n_126), .B2(n_127), .Y(n_125) );
INVx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_103), .A2(n_149), .B(n_150), .Y(n_148) );
AOI21x1_ASAP7_75t_L g213 ( .A1(n_103), .A2(n_214), .B(n_215), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_103), .Y(n_225) );
BUFx12f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx5_ASAP7_75t_L g116 ( .A(n_104), .Y(n_116) );
INVx5_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_104), .A2(n_181), .B1(n_182), .B2(n_184), .Y(n_180) );
OAI321xp33_ASAP7_75t_L g188 ( .A1(n_104), .A2(n_106), .A3(n_128), .B1(n_189), .B2(n_190), .C(n_191), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_106), .A2(n_145), .B(n_146), .C(n_147), .Y(n_144) );
INVx2_ASAP7_75t_SL g166 ( .A(n_106), .Y(n_166) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_107), .Y(n_109) );
INVx1_ASAP7_75t_L g113 ( .A(n_107), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_107), .Y(n_114) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_107), .Y(n_129) );
INVx2_ASAP7_75t_L g211 ( .A(n_107), .Y(n_211) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g151 ( .A(n_109), .Y(n_151) );
INVx2_ASAP7_75t_L g161 ( .A(n_109), .Y(n_161) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g130 ( .A(n_113), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_115), .A2(n_225), .B1(n_226), .B2(n_227), .Y(n_224) );
CKINVDCx6p67_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
AOI21x1_ASAP7_75t_L g177 ( .A1(n_116), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_116), .A2(n_193), .B(n_198), .Y(n_192) );
AOI21x1_ASAP7_75t_L g208 ( .A1(n_116), .A2(n_209), .B(n_212), .Y(n_208) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVxp67_ASAP7_75t_L g255 ( .A(n_118), .Y(n_255) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_121), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_121), .B(n_153), .Y(n_152) );
NOR2x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_137), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_123), .B(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_123), .Y(n_339) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g265 ( .A(n_124), .Y(n_265) );
INVx1_ASAP7_75t_L g289 ( .A(n_124), .Y(n_289) );
AND2x2_ASAP7_75t_L g365 ( .A(n_124), .B(n_253), .Y(n_365) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_124), .Y(n_377) );
AO31x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_131), .A3(n_133), .B(n_134), .Y(n_124) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g183 ( .A(n_129), .Y(n_183) );
INVx2_ASAP7_75t_L g197 ( .A(n_129), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_129), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g483 ( .A(n_129), .Y(n_483) );
INVx3_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx3_ASAP7_75t_L g156 ( .A(n_132), .Y(n_156) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_132), .Y(n_254) );
AND2x2_ASAP7_75t_L g223 ( .A(n_133), .B(n_156), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
INVx1_ASAP7_75t_L g142 ( .A(n_135), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_135), .B(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g395 ( .A(n_138), .Y(n_395) );
AND2x2_ASAP7_75t_L g455 ( .A(n_138), .B(n_234), .Y(n_455) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_154), .Y(n_138) );
INVx2_ASAP7_75t_L g236 ( .A(n_139), .Y(n_236) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g278 ( .A(n_140), .Y(n_278) );
AND2x2_ASAP7_75t_L g354 ( .A(n_140), .B(n_154), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_148), .B(n_152), .Y(n_143) );
NAND2xp33_ASAP7_75t_L g480 ( .A(n_147), .B(n_481), .Y(n_480) );
BUFx3_ASAP7_75t_L g257 ( .A(n_154), .Y(n_257) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_168), .Y(n_154) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_155), .A2(n_157), .B(n_168), .Y(n_238) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_162), .Y(n_158) );
INVxp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_167), .Y(n_163) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_170), .B(n_387), .Y(n_386) );
AOI32xp33_ASAP7_75t_L g432 ( .A1(n_170), .A2(n_411), .A3(n_433), .B1(n_435), .B2(n_438), .Y(n_432) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_171), .B(n_280), .Y(n_425) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g443 ( .A(n_172), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_186), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g248 ( .A(n_174), .Y(n_248) );
AND2x2_ASAP7_75t_L g272 ( .A(n_174), .B(n_186), .Y(n_272) );
OAI21x1_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_185), .Y(n_174) );
OAI21x1_ASAP7_75t_L g206 ( .A1(n_175), .A2(n_207), .B(n_219), .Y(n_206) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_175), .A2(n_207), .B(n_219), .Y(n_243) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_175), .A2(n_176), .B(n_185), .Y(n_287) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_183), .B(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g284 ( .A(n_186), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g298 ( .A(n_186), .B(n_249), .Y(n_298) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g220 ( .A(n_187), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g244 ( .A(n_187), .Y(n_244) );
OAI21x1_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_192), .B(n_200), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_196), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_220), .Y(n_203) );
AND2x2_ASAP7_75t_L g396 ( .A(n_204), .B(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_205), .B(n_244), .Y(n_421) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_205), .Y(n_428) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g281 ( .A(n_206), .Y(n_281) );
OAI21x1_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_213), .B(n_218), .Y(n_207) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g228 ( .A(n_211), .Y(n_228) );
INVx4_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g299 ( .A(n_220), .B(n_248), .Y(n_299) );
AND2x2_ASAP7_75t_L g397 ( .A(n_220), .B(n_315), .Y(n_397) );
BUFx3_ASAP7_75t_L g429 ( .A(n_220), .Y(n_429) );
INVx1_ASAP7_75t_L g449 ( .A(n_220), .Y(n_449) );
OR2x2_ASAP7_75t_L g280 ( .A(n_221), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g320 ( .A(n_221), .Y(n_320) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_221), .Y(n_473) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
AOI21x1_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_229), .Y(n_222) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_231), .A2(n_424), .B1(n_426), .B2(n_427), .Y(n_423) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g338 ( .A(n_232), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
INVx2_ASAP7_75t_L g306 ( .A(n_233), .Y(n_306) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g330 ( .A(n_234), .B(n_309), .Y(n_330) );
INVx1_ASAP7_75t_L g372 ( .A(n_235), .Y(n_372) );
AND2x2_ASAP7_75t_L g383 ( .A(n_235), .B(n_344), .Y(n_383) );
AND2x2_ASAP7_75t_L g406 ( .A(n_235), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
AND2x2_ASAP7_75t_L g252 ( .A(n_236), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g268 ( .A(n_236), .Y(n_268) );
AND2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g361 ( .A(n_237), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_237), .B(n_278), .Y(n_470) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g301 ( .A(n_238), .B(n_253), .Y(n_301) );
OAI21xp33_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_245), .B(n_250), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g335 ( .A(n_243), .Y(n_335) );
AND2x2_ASAP7_75t_L g261 ( .A(n_244), .B(n_249), .Y(n_261) );
INVx2_ASAP7_75t_L g316 ( .A(n_244), .Y(n_316) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_246), .A2(n_312), .B(n_403), .C(n_405), .Y(n_402) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_249), .Y(n_444) );
NOR2x1p5_ASAP7_75t_SL g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g273 ( .A(n_252), .B(n_264), .Y(n_273) );
INVx2_ASAP7_75t_L g308 ( .A(n_257), .Y(n_308) );
AND2x2_ASAP7_75t_L g453 ( .A(n_257), .B(n_365), .Y(n_453) );
NOR2xp67_ASAP7_75t_L g460 ( .A(n_257), .B(n_461), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_274), .C(n_290), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B1(n_270), .B2(n_273), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g367 ( .A(n_261), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g379 ( .A(n_261), .B(n_296), .Y(n_379) );
INVx2_ASAP7_75t_L g414 ( .A(n_261), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_261), .B(n_417), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_262), .A2(n_291), .B1(n_299), .B2(n_300), .Y(n_290) );
NOR2x1p5_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g277 ( .A(n_265), .Y(n_277) );
AND2x4_ASAP7_75t_L g309 ( .A(n_265), .B(n_278), .Y(n_309) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NOR2xp67_ASAP7_75t_L g288 ( .A(n_268), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g326 ( .A(n_268), .Y(n_326) );
OR2x6_ASAP7_75t_L g446 ( .A(n_269), .B(n_363), .Y(n_446) );
AND2x2_ASAP7_75t_L g458 ( .A(n_269), .B(n_354), .Y(n_458) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_SL g279 ( .A(n_272), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g331 ( .A(n_272), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_272), .B(n_312), .Y(n_389) );
AND2x2_ASAP7_75t_L g475 ( .A(n_272), .B(n_333), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B1(n_282), .B2(n_288), .Y(n_274) );
AND2x4_ASAP7_75t_L g300 ( .A(n_276), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVxp67_ASAP7_75t_L g461 ( .A(n_277), .Y(n_461) );
OR2x2_ASAP7_75t_L g283 ( .A(n_280), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g348 ( .A(n_280), .Y(n_348) );
INVx2_ASAP7_75t_L g293 ( .A(n_281), .Y(n_293) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_281), .Y(n_388) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g439 ( .A(n_285), .B(n_293), .Y(n_439) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_SL g342 ( .A(n_286), .Y(n_342) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g297 ( .A(n_287), .Y(n_297) );
AND2x2_ASAP7_75t_L g471 ( .A(n_288), .B(n_301), .Y(n_471) );
INVx1_ASAP7_75t_L g351 ( .A(n_289), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
OR2x2_ASAP7_75t_L g318 ( .A(n_292), .B(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g312 ( .A(n_293), .Y(n_312) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_295), .Y(n_382) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_297), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g373 ( .A(n_298), .B(n_344), .Y(n_373) );
OR2x2_ASAP7_75t_L g456 ( .A(n_298), .B(n_312), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g464 ( .A(n_298), .B(n_315), .Y(n_464) );
INVx1_ASAP7_75t_L g400 ( .A(n_299), .Y(n_400) );
INVx2_ASAP7_75t_L g415 ( .A(n_300), .Y(n_415) );
AOI211x1_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_310), .B(n_317), .C(n_336), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_306), .A2(n_393), .B(n_396), .C(n_398), .Y(n_392) );
INVx1_ASAP7_75t_L g390 ( .A(n_307), .Y(n_390) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_308), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_308), .B(n_323), .Y(n_426) );
INVx2_ASAP7_75t_L g363 ( .A(n_309), .Y(n_363) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx4_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
BUFx2_ASAP7_75t_L g404 ( .A(n_316), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_327), .Y(n_317) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_319), .Y(n_358) );
AND2x2_ASAP7_75t_L g334 ( .A(n_320), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g345 ( .A(n_320), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_321), .A2(n_337), .B(n_340), .Y(n_336) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_323), .B(n_326), .Y(n_329) );
AND2x2_ASAP7_75t_L g410 ( .A(n_323), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVxp67_ASAP7_75t_L g407 ( .A(n_324), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_324), .B(n_470), .Y(n_476) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B(n_331), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AO22x1_ASAP7_75t_L g442 ( .A1(n_330), .A2(n_443), .B1(n_445), .B2(n_447), .Y(n_442) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g344 ( .A(n_335), .Y(n_344) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AND2x2_ASAP7_75t_L g347 ( .A(n_342), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g417 ( .A(n_342), .B(n_369), .Y(n_417) );
INVx1_ASAP7_75t_L g434 ( .A(n_343), .Y(n_434) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx2_ASAP7_75t_L g369 ( .A(n_344), .Y(n_369) );
AOI211xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_349), .B(n_357), .C(n_370), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_351), .B1(n_381), .B2(n_384), .C(n_385), .Y(n_380) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
AND2x2_ASAP7_75t_L g375 ( .A(n_354), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g412 ( .A(n_354), .Y(n_412) );
INVx1_ASAP7_75t_L g437 ( .A(n_355), .Y(n_437) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_364), .B2(n_366), .Y(n_357) );
INVx1_ASAP7_75t_L g441 ( .A(n_359), .Y(n_441) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI22xp33_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_373), .B1(n_374), .B2(n_378), .Y(n_370) );
INVx1_ASAP7_75t_L g384 ( .A(n_373), .Y(n_384) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx2_ASAP7_75t_L g399 ( .A(n_383), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B(n_390), .Y(n_385) );
OR2x2_ASAP7_75t_L g413 ( .A(n_387), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND3xp33_ASAP7_75t_SL g391 ( .A(n_392), .B(n_401), .C(n_430), .Y(n_391) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g436 ( .A(n_395), .B(n_437), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_408), .C(n_423), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_413), .B1(n_415), .B2(n_416), .C(n_418), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_421), .B(n_473), .Y(n_472) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_429), .B(n_441), .Y(n_440) );
NOR4xp25_ASAP7_75t_L g430 ( .A(n_431), .B(n_442), .C(n_450), .D(n_465), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_432), .B(n_440), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_437), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g448 ( .A(n_439), .B(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_451), .B(n_457), .Y(n_450) );
AO21x1_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_454), .B(n_456), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_462), .Y(n_457) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_466), .B(n_474), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_471), .B(n_472), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
AO21x1_ASAP7_75t_L g723 ( .A1(n_480), .A2(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_537), .B1(n_712), .B2(n_714), .C(n_717), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_503), .B1(n_532), .B2(n_533), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_486), .A2(n_532), .B1(n_719), .B2(n_720), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_492), .B1(n_493), .B2(n_502), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_487), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g491 ( .A(n_490), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_500), .B2(n_501), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_496), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_497), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_504), .Y(n_719) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_508), .Y(n_504) );
OR2x4_ASAP7_75t_L g536 ( .A(n_505), .B(n_509), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_506), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g724 ( .A(n_506), .Y(n_724) );
INVx1_ASAP7_75t_L g716 ( .A(n_507), .Y(n_716) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI31xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_515), .A3(n_522), .B(n_524), .Y(n_509) );
BUFx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
BUFx3_ASAP7_75t_L g573 ( .A(n_512), .Y(n_573) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
AND2x4_ASAP7_75t_L g592 ( .A(n_513), .B(n_530), .Y(n_592) );
INVx2_ASAP7_75t_L g530 ( .A(n_514), .Y(n_530) );
INVxp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g531 ( .A(n_518), .Y(n_531) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x4_ASAP7_75t_L g578 ( .A(n_520), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g556 ( .A(n_521), .B(n_549), .Y(n_556) );
AND2x2_ASAP7_75t_L g562 ( .A(n_521), .B(n_563), .Y(n_562) );
INVx6_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVxp67_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
BUFx2_ASAP7_75t_L g583 ( .A(n_527), .Y(n_583) );
AND2x4_ASAP7_75t_L g599 ( .A(n_527), .B(n_531), .Y(n_599) );
AND2x4_ASAP7_75t_L g601 ( .A(n_527), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g621 ( .A(n_527), .B(n_578), .Y(n_621) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx8_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g720 ( .A(n_535), .Y(n_720) );
INVx8_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_537), .A2(n_718), .B1(n_721), .B2(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_622), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_604), .B1(n_608), .B2(n_609), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_557), .C(n_584), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_552), .B2(n_553), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_543), .A2(n_565), .B1(n_701), .B2(n_702), .Y(n_700) );
INVx6_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
OR2x2_ASAP7_75t_L g554 ( .A(n_546), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g564 ( .A(n_546), .Y(n_564) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_L g568 ( .A(n_551), .B(n_563), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_552), .A2(n_587), .B1(n_694), .B2(n_697), .Y(n_693) );
INVx4_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_556), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_565), .B1(n_566), .B2(n_574), .C(n_582), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
AND2x4_ASAP7_75t_L g582 ( .A(n_561), .B(n_583), .Y(n_582) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_562), .Y(n_571) );
INVx2_ASAP7_75t_L g579 ( .A(n_563), .Y(n_579) );
AND2x2_ASAP7_75t_L g585 ( .A(n_564), .B(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_568), .Y(n_586) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_568), .Y(n_594) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx6_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g590 ( .A(n_578), .Y(n_590) );
INVx1_ASAP7_75t_L g603 ( .A(n_579), .Y(n_603) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g596 ( .A(n_581), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .B1(n_588), .B2(n_593), .C(n_597), .Y(n_584) );
INVx2_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
BUFx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
CKINVDCx8_ASAP7_75t_R g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x6_ASAP7_75t_L g669 ( .A(n_607), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_611), .B(n_618), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_616), .Y(n_611) );
INVx2_ASAP7_75t_SL g675 ( .A(n_612), .Y(n_675) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_612), .Y(n_701) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x4_ASAP7_75t_L g629 ( .A(n_614), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g639 ( .A(n_614), .Y(n_639) );
AND2x2_ASAP7_75t_L g645 ( .A(n_614), .B(n_615), .Y(n_645) );
INVx2_ASAP7_75t_L g650 ( .A(n_614), .Y(n_650) );
INVx1_ASAP7_75t_L g682 ( .A(n_614), .Y(n_682) );
INVx2_ASAP7_75t_L g630 ( .A(n_615), .Y(n_630) );
INVx1_ASAP7_75t_L g652 ( .A(n_615), .Y(n_652) );
INVx1_ASAP7_75t_L g659 ( .A(n_615), .Y(n_659) );
INVx1_ASAP7_75t_L g681 ( .A(n_615), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_615), .B(n_650), .Y(n_688) );
INVx3_ASAP7_75t_L g660 ( .A(n_616), .Y(n_660) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_653), .C(n_668), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_624), .B(n_640), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_635), .B2(n_636), .Y(n_624) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_631), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_L g691 ( .A(n_628), .Y(n_691) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g699 ( .A(n_629), .Y(n_699) );
AND2x4_ASAP7_75t_L g638 ( .A(n_630), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g636 ( .A(n_631), .B(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_L g642 ( .A(n_631), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_631), .B(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g708 ( .A(n_632), .Y(n_708) );
INVx1_ASAP7_75t_L g672 ( .A(n_634), .Y(n_672) );
INVx1_ASAP7_75t_L g710 ( .A(n_634), .Y(n_710) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx3_ASAP7_75t_L g667 ( .A(n_638), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_646), .B2(n_647), .Y(n_640) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g664 ( .A(n_650), .Y(n_664) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2x1_ASAP7_75t_SL g656 ( .A(n_657), .B(n_660), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_660), .B(n_663), .Y(n_662) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_660), .B(n_667), .Y(n_666) );
BUFx4f_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI33xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_673), .A3(n_684), .B1(n_693), .B2(n_700), .B3(n_705), .Y(n_668) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B1(n_677), .B2(n_683), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_681), .B(n_682), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g696 ( .A(n_688), .Y(n_696) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx3_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx6_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x6_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
BUFx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx2_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
endmodule