module fake_jpeg_3406_n_686 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_686);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_686;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_332;
wire n_92;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_19),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_7),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_62),
.B(n_72),
.Y(n_179)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_0),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_74),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_41),
.B(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_77),
.Y(n_187)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_79),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_80),
.B(n_81),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_0),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_82),
.B(n_88),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_86),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_87),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_40),
.Y(n_88)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_89),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_40),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_90),
.B(n_94),
.Y(n_166)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_91),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_47),
.B(n_1),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_92),
.B(n_5),
.Y(n_211)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_93),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_40),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g186 ( 
.A(n_95),
.Y(n_186)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_97),
.Y(n_225)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_98),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_38),
.B(n_3),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_99),
.B(n_107),
.Y(n_204)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

CKINVDCx9p33_ASAP7_75t_R g229 ( 
.A(n_102),
.Y(n_229)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_54),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_106),
.B(n_120),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_41),
.B(n_17),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx5_ASAP7_75t_SL g185 ( 
.A(n_110),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_21),
.B(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_112),
.B(n_113),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_17),
.Y(n_113)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_114),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_44),
.B(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_115),
.B(n_118),
.Y(n_212)
);

BUFx8_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_44),
.B(n_3),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_119),
.B(n_123),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_34),
.B(n_18),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_22),
.B(n_4),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_22),
.B(n_4),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_128),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_34),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_34),
.Y(n_130)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_59),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_53),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_46),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_30),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_133),
.B(n_151),
.Y(n_264)
);

INVx6_ASAP7_75t_SL g138 ( 
.A(n_102),
.Y(n_138)
);

CKINVDCx9p33_ASAP7_75t_R g270 ( 
.A(n_138),
.Y(n_270)
);

CKINVDCx12_ASAP7_75t_R g139 ( 
.A(n_102),
.Y(n_139)
);

CKINVDCx12_ASAP7_75t_R g233 ( 
.A(n_139),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_72),
.B(n_80),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_141),
.B(n_162),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g151 ( 
.A(n_125),
.B(n_30),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_119),
.A2(n_43),
.B1(n_58),
.B2(n_57),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_160),
.A2(n_196),
.B1(n_205),
.B2(n_131),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_99),
.B(n_43),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_116),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_164),
.B(n_168),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_81),
.B(n_32),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_116),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_169),
.B(n_181),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_100),
.B(n_28),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_182),
.B(n_190),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_122),
.A2(n_59),
.B1(n_51),
.B2(n_45),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_183),
.A2(n_59),
.B1(n_51),
.B2(n_23),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_115),
.B(n_28),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_118),
.B(n_24),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_201),
.Y(n_231)
);

HAxp5_ASAP7_75t_SL g193 ( 
.A(n_92),
.B(n_46),
.CON(n_193),
.SN(n_193)
);

INVx2_ASAP7_75t_R g300 ( 
.A(n_193),
.Y(n_300)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_71),
.Y(n_195)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_60),
.A2(n_27),
.B1(n_58),
.B2(n_57),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_93),
.Y(n_197)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_63),
.B(n_24),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_121),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_202),
.B(n_217),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_92),
.B(n_45),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_219),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_70),
.A2(n_27),
.B1(n_49),
.B2(n_48),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_76),
.B(n_23),
.C(n_45),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_206),
.B(n_86),
.C(n_67),
.Y(n_268)
);

BUFx12_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_23),
.Y(n_245)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_213),
.Y(n_275)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_96),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_77),
.Y(n_218)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_98),
.B(n_33),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_109),
.B(n_49),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_223),
.Y(n_252)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_103),
.Y(n_222)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_78),
.B(n_48),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_61),
.B(n_36),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_226),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_105),
.B(n_36),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_65),
.B(n_33),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_228),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_126),
.B(n_129),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_124),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_230),
.B(n_117),
.Y(n_283)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_51),
.C(n_30),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_232),
.B(n_277),
.Y(n_341)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_157),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_234),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_136),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_235),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_157),
.Y(n_236)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_236),
.Y(n_354)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_237),
.Y(n_316)
);

INVx13_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_238),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_156),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_242),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_243),
.A2(n_249),
.B1(n_287),
.B2(n_297),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_146),
.A2(n_89),
.B1(n_84),
.B2(n_114),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_244),
.A2(n_247),
.B1(n_249),
.B2(n_287),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_245),
.B(n_246),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_146),
.A2(n_85),
.B1(n_91),
.B2(n_104),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_144),
.A2(n_83),
.B1(n_68),
.B2(n_101),
.Y(n_249)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_138),
.Y(n_251)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

INVx11_ASAP7_75t_L g326 ( 
.A(n_253),
.Y(n_326)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_154),
.Y(n_255)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_255),
.Y(n_335)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_136),
.Y(n_261)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_261),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_221),
.B(n_66),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_263),
.B(n_266),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_156),
.Y(n_265)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_265),
.Y(n_320)
);

CKINVDCx12_ASAP7_75t_R g266 ( 
.A(n_185),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_143),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_267),
.B(n_271),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_268),
.B(n_214),
.Y(n_355)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_154),
.Y(n_269)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_269),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_204),
.B(n_180),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_212),
.B(n_79),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_273),
.B(n_276),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_147),
.Y(n_274)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_274),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_163),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_209),
.B(n_87),
.Y(n_277)
);

AOI21xp33_ASAP7_75t_L g278 ( 
.A1(n_148),
.A2(n_86),
.B(n_53),
.Y(n_278)
);

AOI32xp33_ASAP7_75t_L g339 ( 
.A1(n_278),
.A2(n_300),
.A3(n_270),
.B1(n_231),
.B2(n_257),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_279),
.Y(n_349)
);

INVx5_ASAP7_75t_SL g280 ( 
.A(n_208),
.Y(n_280)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_155),
.Y(n_281)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_159),
.Y(n_282)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_283),
.Y(n_350)
);

CKINVDCx12_ASAP7_75t_R g284 ( 
.A(n_134),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_284),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_147),
.Y(n_285)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_159),
.Y(n_286)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_144),
.A2(n_111),
.B1(n_97),
.B2(n_69),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_166),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_289),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_175),
.B(n_86),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_203),
.A2(n_53),
.B1(n_7),
.B2(n_8),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_290),
.A2(n_310),
.B1(n_293),
.B2(n_260),
.Y(n_331)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_218),
.Y(n_291)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_195),
.Y(n_292)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_6),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_296),
.Y(n_327)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_222),
.Y(n_294)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_177),
.B(n_7),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_295),
.B(n_299),
.Y(n_364)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_152),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_144),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_297),
.A2(n_309),
.B(n_310),
.Y(n_334)
);

CKINVDCx12_ASAP7_75t_R g298 ( 
.A(n_170),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_298),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_191),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_304),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_L g302 ( 
.A1(n_183),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_193),
.B1(n_206),
.B2(n_186),
.Y(n_322)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_191),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_152),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_305),
.B(n_306),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_173),
.B(n_10),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_176),
.B(n_15),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_308),
.Y(n_343)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_140),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_178),
.B(n_133),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_211),
.B(n_15),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_199),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_311),
.B(n_312),
.Y(n_373)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_194),
.Y(n_312)
);

CKINVDCx12_ASAP7_75t_R g313 ( 
.A(n_186),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g340 ( 
.A(n_313),
.B(n_314),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g314 ( 
.A(n_140),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_322),
.A2(n_323),
.B1(n_359),
.B2(n_368),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_264),
.A2(n_194),
.B1(n_158),
.B2(n_187),
.Y(n_323)
);

OAI22x1_ASAP7_75t_SL g329 ( 
.A1(n_264),
.A2(n_155),
.B1(n_151),
.B2(n_214),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_329),
.A2(n_336),
.B1(n_346),
.B2(n_357),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_268),
.A2(n_207),
.B(n_216),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_330),
.A2(n_244),
.B(n_270),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_331),
.B(n_258),
.Y(n_384)
);

OA22x2_ASAP7_75t_SL g332 ( 
.A1(n_300),
.A2(n_199),
.B1(n_167),
.B2(n_137),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g386 ( 
.A(n_332),
.B(n_282),
.C(n_255),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_248),
.A2(n_187),
.B1(n_158),
.B2(n_210),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g408 ( 
.A(n_339),
.B(n_251),
.C(n_305),
.Y(n_408)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_289),
.A2(n_184),
.B1(n_225),
.B2(n_171),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_252),
.A2(n_225),
.B1(n_188),
.B2(n_171),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_348),
.A2(n_351),
.B1(n_361),
.B2(n_365),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_240),
.A2(n_165),
.B1(n_188),
.B2(n_172),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_355),
.B(n_308),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_243),
.A2(n_210),
.B1(n_142),
.B2(n_167),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_302),
.A2(n_142),
.B1(n_137),
.B2(n_189),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_245),
.A2(n_150),
.B1(n_198),
.B2(n_165),
.Y(n_361)
);

AO22x1_ASAP7_75t_SL g366 ( 
.A1(n_312),
.A2(n_189),
.B1(n_200),
.B2(n_150),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_376),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_259),
.A2(n_172),
.B1(n_198),
.B2(n_174),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_239),
.A2(n_153),
.B1(n_145),
.B2(n_216),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_371),
.A2(n_145),
.B1(n_238),
.B2(n_256),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g375 ( 
.A(n_254),
.B(n_161),
.CI(n_153),
.CON(n_375),
.SN(n_375)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_375),
.B(n_303),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_247),
.A2(n_200),
.B1(n_174),
.B2(n_149),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_377),
.Y(n_426)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_378),
.Y(n_436)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_379),
.Y(n_460)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_373),
.Y(n_380)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_382),
.B(n_384),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_385),
.A2(n_418),
.B(n_424),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_386),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_275),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_387),
.B(n_389),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_388),
.A2(n_407),
.B1(n_420),
.B2(n_421),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_374),
.B(n_304),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_317),
.A2(n_135),
.B1(n_149),
.B2(n_261),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_391),
.A2(n_400),
.B1(n_416),
.B2(n_423),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_301),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_392),
.B(n_393),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_280),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_394),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_345),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_396),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_343),
.B(n_241),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_397),
.B(n_415),
.Y(n_451)
);

INVx8_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_317),
.A2(n_135),
.B1(n_294),
.B2(n_291),
.Y(n_400)
);

A2O1A1Ixp33_ASAP7_75t_L g401 ( 
.A1(n_330),
.A2(n_262),
.B(n_272),
.C(n_233),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_401),
.A2(n_409),
.B(n_413),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_343),
.B(n_292),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_402),
.B(n_403),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_367),
.B(n_241),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_404),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_405),
.Y(n_433)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_360),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_SL g437 ( 
.A(n_408),
.B(n_411),
.C(n_425),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_269),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_347),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_410),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_356),
.B(n_286),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_358),
.B(n_314),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_355),
.B(n_296),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_317),
.A2(n_285),
.B1(n_274),
.B2(n_235),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_349),
.B(n_314),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_417),
.A2(n_419),
.B(n_422),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_340),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_341),
.B(n_253),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_333),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_325),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_319),
.B(n_253),
.Y(n_422)
);

INVx8_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_327),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_327),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_398),
.A2(n_322),
.B1(n_353),
.B2(n_359),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_427),
.B(n_431),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_329),
.C(n_327),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_429),
.B(n_439),
.C(n_443),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_398),
.A2(n_323),
.B1(n_368),
.B2(n_365),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_398),
.A2(n_332),
.B1(n_375),
.B2(n_334),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_438),
.B(n_441),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_340),
.C(n_320),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_383),
.A2(n_380),
.B1(n_378),
.B2(n_412),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_383),
.A2(n_332),
.B1(n_375),
.B2(n_334),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_448),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_340),
.C(n_336),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_403),
.B(n_325),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_447),
.B(n_452),
.C(n_453),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_412),
.A2(n_357),
.B1(n_376),
.B2(n_337),
.Y(n_448)
);

AO21x2_ASAP7_75t_SL g449 ( 
.A1(n_386),
.A2(n_401),
.B(n_385),
.Y(n_449)
);

AO22x2_ASAP7_75t_L g488 ( 
.A1(n_449),
.A2(n_438),
.B1(n_442),
.B2(n_441),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_418),
.B(n_384),
.C(n_396),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_389),
.B(n_328),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_402),
.A2(n_337),
.B1(n_342),
.B2(n_328),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_459),
.A2(n_414),
.B1(n_416),
.B2(n_391),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_414),
.A2(n_342),
.B1(n_370),
.B2(n_363),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_461),
.A2(n_379),
.B1(n_381),
.B2(n_394),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_411),
.B(n_338),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_462),
.B(n_390),
.Y(n_474)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_467),
.Y(n_524)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_465),
.Y(n_468)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_468),
.Y(n_527)
);

INVx13_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_469),
.Y(n_514)
);

INVx13_ASAP7_75t_L g470 ( 
.A(n_449),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_470),
.A2(n_475),
.B1(n_479),
.B2(n_485),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_471),
.A2(n_432),
.B1(n_461),
.B2(n_458),
.Y(n_520)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_465),
.Y(n_472)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_472),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_454),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_459),
.Y(n_476)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_476),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_436),
.A2(n_407),
.B1(n_392),
.B2(n_393),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_477),
.A2(n_484),
.B1(n_434),
.B2(n_443),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_450),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_460),
.Y(n_480)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_480),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_428),
.B(n_387),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_481),
.B(n_482),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_456),
.B(n_362),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_430),
.B(n_372),
.Y(n_483)
);

CKINVDCx14_ASAP7_75t_R g531 ( 
.A(n_483),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_436),
.A2(n_382),
.B1(n_408),
.B2(n_418),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_450),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_486),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_445),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_487),
.B(n_496),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_488),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_444),
.A2(n_422),
.B(n_413),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_489),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_430),
.B(n_417),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_490),
.B(n_491),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_433),
.B(n_419),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_433),
.B(n_352),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_495),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_444),
.A2(n_377),
.B(n_409),
.Y(n_493)
);

XNOR2x1_ASAP7_75t_SL g530 ( 
.A(n_493),
.B(n_429),
.Y(n_530)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

NAND3xp33_ASAP7_75t_L g495 ( 
.A(n_452),
.B(n_421),
.C(n_406),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_460),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_457),
.B(n_400),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_497),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_445),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_498),
.B(n_503),
.Y(n_523)
);

BUFx24_ASAP7_75t_L g500 ( 
.A(n_449),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_500),
.Y(n_518)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_466),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_505),
.Y(n_519)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_455),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_455),
.Y(n_505)
);

AND2x4_ASAP7_75t_SL g506 ( 
.A(n_493),
.B(n_434),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_506),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_510),
.B(n_533),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_473),
.A2(n_427),
.B1(n_431),
.B2(n_448),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_512),
.A2(n_516),
.B1(n_533),
.B2(n_537),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_473),
.A2(n_504),
.B1(n_499),
.B2(n_476),
.Y(n_516)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_484),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_517),
.B(n_426),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_520),
.A2(n_467),
.B1(n_469),
.B2(n_498),
.Y(n_572)
);

AO22x1_ASAP7_75t_SL g521 ( 
.A1(n_500),
.A2(n_464),
.B1(n_432),
.B2(n_453),
.Y(n_521)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_521),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_502),
.B(n_451),
.Y(n_525)
);

XNOR2x1_ASAP7_75t_L g549 ( 
.A(n_525),
.B(n_478),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_477),
.B(n_440),
.Y(n_526)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_526),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_530),
.A2(n_488),
.B(n_500),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_504),
.A2(n_464),
.B1(n_447),
.B2(n_463),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_502),
.B(n_435),
.Y(n_534)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_534),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_503),
.B(n_435),
.Y(n_536)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_536),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_499),
.A2(n_426),
.B1(n_457),
.B2(n_462),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_505),
.B(n_352),
.Y(n_540)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_540),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_486),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_541),
.B(n_487),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_478),
.B(n_451),
.C(n_439),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_489),
.C(n_437),
.Y(n_558)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_519),
.Y(n_546)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_546),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_547),
.A2(n_570),
.B1(n_572),
.B2(n_446),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_549),
.B(n_571),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_550),
.B(n_553),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_531),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_564),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_552),
.B(n_423),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_515),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_511),
.A2(n_514),
.B(n_518),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_554),
.A2(n_522),
.B(n_524),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_506),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_527),
.Y(n_559)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_559),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_479),
.C(n_485),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_560),
.B(n_561),
.C(n_565),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_525),
.B(n_437),
.C(n_468),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_512),
.A2(n_471),
.B1(n_488),
.B2(n_497),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_562),
.A2(n_528),
.B1(n_518),
.B2(n_514),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_523),
.B(n_472),
.Y(n_563)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_563),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_508),
.B(n_338),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_530),
.B(n_497),
.C(n_480),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_539),
.B(n_496),
.C(n_321),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_566),
.B(n_569),
.C(n_576),
.Y(n_602)
);

AO21x1_ASAP7_75t_L g586 ( 
.A1(n_567),
.A2(n_509),
.B(n_516),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_523),
.B(n_501),
.Y(n_568)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_568),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_510),
.B(n_321),
.C(n_363),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_528),
.A2(n_488),
.B1(n_500),
.B2(n_470),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_537),
.B(n_488),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_527),
.Y(n_573)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_573),
.Y(n_584)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_529),
.Y(n_575)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_575),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_508),
.B(n_335),
.C(n_354),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_580),
.B(n_597),
.Y(n_622)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_582),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_585),
.A2(n_587),
.B1(n_601),
.B2(n_575),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_586),
.A2(n_600),
.B(n_567),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_562),
.A2(n_535),
.B1(n_524),
.B2(n_506),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_588),
.A2(n_598),
.B1(n_545),
.B2(n_573),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_547),
.A2(n_535),
.B1(n_521),
.B2(n_532),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_590),
.B(n_591),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_544),
.A2(n_572),
.B1(n_554),
.B2(n_570),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_560),
.B(n_569),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_592),
.B(n_565),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_563),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_596),
.B(n_542),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_561),
.B(n_521),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_548),
.A2(n_522),
.B1(n_529),
.B2(n_541),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_568),
.Y(n_599)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_599),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_544),
.A2(n_538),
.B1(n_507),
.B2(n_513),
.Y(n_601)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_604),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_605),
.Y(n_634)
);

AOI21xp33_ASAP7_75t_L g606 ( 
.A1(n_581),
.A2(n_553),
.B(n_556),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_606),
.B(n_609),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_581),
.A2(n_557),
.B(n_558),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_608),
.B(n_616),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_592),
.B(n_549),
.C(n_571),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_610),
.B(n_612),
.Y(n_628)
);

BUFx12f_ASAP7_75t_SL g611 ( 
.A(n_594),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_611),
.A2(n_617),
.B(n_586),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_602),
.B(n_548),
.C(n_576),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_602),
.B(n_566),
.C(n_555),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_613),
.B(n_615),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_597),
.B(n_546),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_614),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_589),
.B(n_559),
.C(n_550),
.Y(n_615)
);

BUFx12f_ASAP7_75t_SL g617 ( 
.A(n_594),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_593),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_618),
.B(n_620),
.Y(n_639)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_578),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_589),
.B(n_538),
.C(n_574),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_621),
.B(n_622),
.C(n_615),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_590),
.B(n_542),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_623),
.B(n_598),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_624),
.A2(n_584),
.B1(n_595),
.B2(n_599),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_625),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_627),
.B(n_630),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_629),
.B(n_637),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_612),
.B(n_580),
.C(n_591),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_621),
.B(n_577),
.Y(n_631)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_631),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_635),
.A2(n_421),
.B1(n_423),
.B2(n_399),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_604),
.B(n_587),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_613),
.B(n_588),
.C(n_601),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_640),
.B(n_641),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_609),
.B(n_585),
.C(n_579),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_614),
.B(n_583),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g655 ( 
.A(n_642),
.B(n_421),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_627),
.B(n_607),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_643),
.B(n_646),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_630),
.B(n_610),
.C(n_603),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_639),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_647),
.B(n_650),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_626),
.B(n_618),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_632),
.A2(n_623),
.B(n_619),
.Y(n_651)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_651),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_638),
.A2(n_617),
.B(n_611),
.Y(n_652)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_652),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_636),
.A2(n_513),
.B1(n_494),
.B2(n_420),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_653),
.B(n_654),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_655),
.B(n_629),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_628),
.B(n_420),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_656),
.B(n_640),
.Y(n_667)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_658),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_648),
.B(n_633),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_662),
.A2(n_663),
.B1(n_667),
.B2(n_335),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_648),
.B(n_641),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_657),
.A2(n_638),
.B(n_634),
.Y(n_664)
);

AOI31xp67_ASAP7_75t_SL g675 ( 
.A1(n_664),
.A2(n_250),
.A3(n_366),
.B(n_388),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_644),
.B(n_634),
.C(n_642),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_668),
.B(n_657),
.C(n_646),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_669),
.A2(n_675),
.B(n_668),
.Y(n_676)
);

AOI322xp5_ASAP7_75t_L g670 ( 
.A1(n_664),
.A2(n_649),
.A3(n_637),
.B1(n_645),
.B2(n_653),
.C1(n_655),
.C2(n_420),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_SL g678 ( 
.A1(n_670),
.A2(n_671),
.B1(n_673),
.B2(n_316),
.Y(n_678)
);

AOI322xp5_ASAP7_75t_L g671 ( 
.A1(n_661),
.A2(n_399),
.A3(n_370),
.B1(n_326),
.B2(n_161),
.C1(n_250),
.C2(n_315),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_SL g677 ( 
.A1(n_672),
.A2(n_660),
.B(n_659),
.Y(n_677)
);

AOI322xp5_ASAP7_75t_L g673 ( 
.A1(n_666),
.A2(n_326),
.A3(n_250),
.B1(n_315),
.B2(n_318),
.C1(n_354),
.C2(n_366),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_676),
.B(n_677),
.Y(n_681)
);

AOI322xp5_ASAP7_75t_L g680 ( 
.A1(n_678),
.A2(n_679),
.A3(n_670),
.B1(n_236),
.B2(n_665),
.C1(n_237),
.C2(n_207),
.Y(n_680)
);

A2O1A1O1Ixp25_ASAP7_75t_L g679 ( 
.A1(n_674),
.A2(n_665),
.B(n_316),
.C(n_281),
.D(n_234),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_680),
.B(n_15),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_682),
.B(n_681),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_683),
.B(n_12),
.Y(n_684)
);

AO21x1_ASAP7_75t_L g685 ( 
.A1(n_684),
.A2(n_12),
.B(n_13),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_SL g686 ( 
.A(n_685),
.B(n_12),
.C(n_13),
.Y(n_686)
);


endmodule