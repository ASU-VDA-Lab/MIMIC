module fake_jpeg_9547_n_226 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_1),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_26),
.B1(n_22),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_48),
.A2(n_55),
.B1(n_57),
.B2(n_21),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_56),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_22),
.B1(n_25),
.B2(n_19),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_69),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_73),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_71),
.B(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_29),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_23),
.Y(n_80)
);

AO22x1_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_114)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_21),
.B(n_34),
.Y(n_86)
);

OAI22x1_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_97),
.B1(n_10),
.B2(n_12),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_3),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_17),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_24),
.B(n_29),
.C(n_32),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_28),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_99),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_3),
.Y(n_99)
);

NOR2xp67_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_111),
.Y(n_128)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_17),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_93),
.B(n_90),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_9),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_12),
.C(n_14),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_4),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_67),
.Y(n_132)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_76),
.B1(n_70),
.B2(n_68),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_82),
.B1(n_86),
.B2(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_125),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_101),
.B(n_114),
.Y(n_147)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_92),
.B(n_90),
.C(n_88),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_139),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_88),
.B1(n_83),
.B2(n_87),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_131),
.B1(n_74),
.B2(n_110),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_83),
.B1(n_87),
.B2(n_67),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_116),
.B(n_106),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_109),
.B(n_118),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_75),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_15),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_15),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_127),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_98),
.B(n_101),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_155),
.B(n_164),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_153),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_74),
.B(n_103),
.Y(n_155)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_145),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_16),
.B(n_126),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_176),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_125),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_128),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_181),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_135),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_164),
.B(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_134),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_152),
.C(n_165),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_187),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_158),
.C(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_158),
.C(n_154),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_166),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_182),
.C(n_191),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_161),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_196),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_173),
.B(n_147),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_156),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_188),
.B(n_160),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_203),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_208),
.B(n_201),
.Y(n_212)
);

OAI211xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_149),
.B(n_176),
.C(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_202),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_186),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_213),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);

AOI31xp67_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_200),
.A3(n_154),
.B(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_207),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_210),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_208),
.B(n_137),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_204),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_222),
.C(n_123),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_216),
.Y(n_226)
);


endmodule