module real_aes_17359_n_266 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_1523, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_266);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_1523;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_266;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_273;
wire n_1038;
wire n_1085;
wire n_276;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_0), .A2(n_71), .B1(n_314), .B2(n_333), .Y(n_332) );
INVxp33_ASAP7_75t_SL g438 ( .A(n_0), .Y(n_438) );
OAI22xp33_ASAP7_75t_L g1167 ( .A1(n_1), .A2(n_91), .B1(n_687), .B2(n_690), .Y(n_1167) );
INVxp67_ASAP7_75t_SL g1181 ( .A(n_1), .Y(n_1181) );
XOR2xp5_ASAP7_75t_L g1110 ( .A(n_2), .B(n_1111), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g1299 ( .A1(n_3), .A2(n_205), .B1(n_1260), .B2(n_1264), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_4), .A2(n_215), .B1(n_804), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_4), .A2(n_189), .B1(n_552), .B2(n_826), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g921 ( .A(n_5), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g1478 ( .A1(n_6), .A2(n_85), .B1(n_782), .B2(n_1479), .C(n_1480), .Y(n_1478) );
AOI22xp33_ASAP7_75t_SL g1502 ( .A1(n_6), .A2(n_142), .B1(n_321), .B2(n_497), .Y(n_1502) );
CKINVDCx5p33_ASAP7_75t_R g1489 ( .A(n_7), .Y(n_1489) );
CKINVDCx5p33_ASAP7_75t_R g1064 ( .A(n_8), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_9), .A2(n_46), .B1(n_804), .B2(n_808), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_9), .A2(n_212), .B1(n_412), .B2(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1153 ( .A(n_10), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_11), .A2(n_56), .B1(n_1260), .B2(n_1264), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1206 ( .A1(n_12), .A2(n_74), .B1(n_472), .B2(n_476), .Y(n_1206) );
OAI22xp33_ASAP7_75t_L g1240 ( .A1(n_12), .A2(n_41), .B1(n_687), .B2(n_690), .Y(n_1240) );
AOI221xp5_ASAP7_75t_L g965 ( .A1(n_13), .A2(n_243), .B1(n_823), .B2(n_966), .C(n_968), .Y(n_965) );
INVx1_ASAP7_75t_L g988 ( .A(n_13), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_14), .A2(n_196), .B1(n_608), .B2(n_693), .C(n_696), .Y(n_692) );
INVx1_ASAP7_75t_L g737 ( .A(n_14), .Y(n_737) );
INVx1_ASAP7_75t_L g281 ( .A(n_15), .Y(n_281) );
AND2x2_ASAP7_75t_L g394 ( .A(n_15), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g407 ( .A(n_15), .B(n_227), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_15), .B(n_291), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_16), .Y(n_1010) );
INVx1_ASAP7_75t_L g756 ( .A(n_17), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_17), .A2(n_40), .B1(n_649), .B2(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g1263 ( .A(n_18), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_18), .B(n_108), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_18), .B(n_1269), .Y(n_1271) );
INVx1_ASAP7_75t_L g800 ( .A(n_19), .Y(n_800) );
OAI221xp5_ASAP7_75t_L g830 ( .A1(n_19), .A2(n_165), .B1(n_831), .B2(n_834), .C(n_839), .Y(n_830) );
AOI21xp5_ASAP7_75t_L g1164 ( .A1(n_20), .A2(n_497), .B(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1194 ( .A(n_20), .Y(n_1194) );
AOI22xp5_ASAP7_75t_L g1281 ( .A1(n_21), .A2(n_37), .B1(n_1267), .B2(n_1270), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_22), .A2(n_157), .B1(n_695), .B2(n_911), .Y(n_1173) );
AOI32xp33_ASAP7_75t_L g1183 ( .A1(n_22), .A2(n_1135), .A3(n_1184), .B1(n_1186), .B2(n_1523), .Y(n_1183) );
OAI222xp33_ASAP7_75t_L g1466 ( .A1(n_23), .A2(n_158), .B1(n_835), .B2(n_1467), .C1(n_1468), .C2(n_1472), .Y(n_1466) );
INVx1_ASAP7_75t_L g1493 ( .A(n_23), .Y(n_1493) );
CKINVDCx5p33_ASAP7_75t_R g1018 ( .A(n_24), .Y(n_1018) );
OAI21xp5_ASAP7_75t_L g1141 ( .A1(n_25), .A2(n_659), .B(n_1142), .Y(n_1141) );
OAI22xp33_ASAP7_75t_L g1042 ( .A1(n_26), .A2(n_254), .B1(n_283), .B2(n_1043), .Y(n_1042) );
OAI22xp33_ASAP7_75t_L g1073 ( .A1(n_26), .A2(n_254), .B1(n_1074), .B2(n_1077), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_27), .B(n_610), .Y(n_1166) );
AOI221xp5_ASAP7_75t_L g1198 ( .A1(n_27), .A2(n_157), .B1(n_639), .B2(n_640), .C(n_942), .Y(n_1198) );
AOI22xp5_ASAP7_75t_L g1298 ( .A1(n_28), .A2(n_128), .B1(n_1267), .B2(n_1270), .Y(n_1298) );
INVx1_ASAP7_75t_L g1140 ( .A(n_29), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_30), .A2(n_76), .B1(n_336), .B2(n_337), .C(n_339), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_30), .A2(n_33), .B1(n_461), .B2(n_462), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_31), .Y(n_523) );
INVx1_ASAP7_75t_L g1126 ( .A(n_32), .Y(n_1126) );
AOI22xp33_ASAP7_75t_SL g304 ( .A1(n_33), .A2(n_141), .B1(n_305), .B2(n_314), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_34), .Y(n_1024) );
CKINVDCx5p33_ASAP7_75t_R g870 ( .A(n_35), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_36), .B(n_1163), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_36), .A2(n_260), .B1(n_635), .B2(n_785), .Y(n_1197) );
INVx1_ASAP7_75t_L g1484 ( .A(n_38), .Y(n_1484) );
INVx1_ASAP7_75t_L g353 ( .A(n_39), .Y(n_353) );
OA222x2_ASAP7_75t_L g400 ( .A1(n_39), .A2(n_175), .B1(n_259), .B2(n_401), .C1(n_408), .C2(n_416), .Y(n_400) );
INVx1_ASAP7_75t_L g769 ( .A(n_40), .Y(n_769) );
OAI211xp5_ASAP7_75t_L g1204 ( .A1(n_41), .A2(n_387), .B(n_1205), .C(n_1222), .Y(n_1204) );
INVx1_ASAP7_75t_L g764 ( .A(n_42), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_42), .A2(n_184), .B1(n_782), .B2(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_43), .A2(n_104), .B1(n_1260), .B2(n_1335), .Y(n_1334) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_44), .A2(n_208), .B1(n_321), .B2(n_323), .C(n_328), .Y(n_320) );
INVx1_ASAP7_75t_L g455 ( .A(n_44), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g1274 ( .A1(n_45), .A2(n_96), .B1(n_1260), .B2(n_1275), .Y(n_1274) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_46), .A2(n_125), .B1(n_636), .B2(n_843), .C(n_1131), .Y(n_1130) );
AOI211xp5_ASAP7_75t_L g676 ( .A1(n_47), .A2(n_336), .B(n_677), .C(n_681), .Y(n_676) );
INVx1_ASAP7_75t_L g729 ( .A(n_47), .Y(n_729) );
INVx1_ASAP7_75t_L g788 ( .A(n_48), .Y(n_788) );
INVx1_ASAP7_75t_L g972 ( .A(n_49), .Y(n_972) );
INVxp67_ASAP7_75t_SL g1473 ( .A(n_50), .Y(n_1473) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_50), .A2(n_85), .B1(n_321), .B2(n_497), .Y(n_1498) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_51), .A2(n_177), .B1(n_671), .B2(n_672), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_51), .A2(n_81), .B1(n_877), .B2(n_879), .Y(n_947) );
INVx1_ASAP7_75t_L g1471 ( .A(n_52), .Y(n_1471) );
AOI22xp33_ASAP7_75t_L g1499 ( .A1(n_52), .A2(n_238), .B1(n_695), .B2(n_911), .Y(n_1499) );
AOI22xp33_ASAP7_75t_SL g1123 ( .A1(n_53), .A2(n_116), .B1(n_307), .B2(n_378), .Y(n_1123) );
AOI221xp5_ASAP7_75t_L g1134 ( .A1(n_53), .A2(n_80), .B1(n_429), .B2(n_637), .C(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g313 ( .A(n_54), .Y(n_313) );
INVx1_ASAP7_75t_L g319 ( .A(n_54), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g1286 ( .A1(n_55), .A2(n_136), .B1(n_1260), .B2(n_1275), .Y(n_1286) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_57), .A2(n_246), .B1(n_355), .B2(n_671), .C(n_672), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_57), .A2(n_132), .B1(n_472), .B2(n_476), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_58), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_59), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_60), .A2(n_225), .B1(n_1267), .B2(n_1270), .Y(n_1336) );
OAI221xp5_ASAP7_75t_L g744 ( .A1(n_61), .A2(n_110), .B1(n_516), .B2(n_674), .C(n_745), .Y(n_744) );
INVxp67_ASAP7_75t_SL g776 ( .A(n_61), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_62), .A2(n_242), .B1(n_516), .B2(n_674), .Y(n_1229) );
INVxp67_ASAP7_75t_SL g1244 ( .A(n_62), .Y(n_1244) );
INVx1_ASAP7_75t_L g274 ( .A(n_63), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_64), .A2(n_220), .B1(n_323), .B2(n_608), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_64), .A2(n_170), .B1(n_646), .B2(n_649), .C(n_650), .Y(n_645) );
INVx2_ASAP7_75t_L g331 ( .A(n_65), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g1019 ( .A(n_66), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_67), .A2(n_238), .B1(n_412), .B2(n_845), .Y(n_1481) );
AOI22xp5_ASAP7_75t_L g1500 ( .A1(n_67), .A2(n_160), .B1(n_911), .B2(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g919 ( .A(n_68), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_68), .A2(n_224), .B1(n_412), .B2(n_461), .Y(n_941) );
INVxp67_ASAP7_75t_SL g955 ( .A(n_69), .Y(n_955) );
OAI211xp5_ASAP7_75t_L g996 ( .A1(n_69), .A2(n_355), .B(n_997), .C(n_998), .Y(n_996) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_70), .Y(n_929) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_71), .Y(n_459) );
INVx1_ASAP7_75t_L g882 ( .A(n_72), .Y(n_882) );
INVx1_ASAP7_75t_L g1105 ( .A(n_73), .Y(n_1105) );
OAI221xp5_ASAP7_75t_L g1228 ( .A1(n_74), .A2(n_126), .B1(n_355), .B2(n_671), .C(n_672), .Y(n_1228) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_75), .A2(n_119), .B1(n_606), .B2(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_75), .A2(n_146), .B1(n_639), .B2(n_640), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_76), .A2(n_208), .B1(n_429), .B2(n_431), .C(n_434), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_77), .Y(n_582) );
INVx1_ASAP7_75t_L g957 ( .A(n_78), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_79), .A2(n_249), .B1(n_1047), .B2(n_1050), .Y(n_1046) );
OAI22xp33_ASAP7_75t_L g1094 ( .A1(n_79), .A2(n_249), .B1(n_1095), .B2(n_1097), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_80), .A2(n_226), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
OAI221xp5_ASAP7_75t_L g926 ( .A1(n_81), .A2(n_176), .B1(n_505), .B2(n_927), .C(n_928), .Y(n_926) );
INVx1_ASAP7_75t_L g374 ( .A(n_82), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_82), .B(n_387), .Y(n_386) );
OAI222xp33_ASAP7_75t_L g888 ( .A1(n_83), .A2(n_133), .B1(n_239), .B2(n_518), .C1(n_682), .C2(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g903 ( .A(n_83), .Y(n_903) );
INVx1_ASAP7_75t_L g767 ( .A(n_84), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_84), .A2(n_229), .B1(n_412), .B2(n_461), .Y(n_783) );
XOR2x2_ASAP7_75t_L g665 ( .A(n_86), .B(n_666), .Y(n_665) );
XOR2x1_ASAP7_75t_L g1148 ( .A(n_87), .B(n_1149), .Y(n_1148) );
AOI22xp5_ASAP7_75t_L g1321 ( .A1(n_87), .A2(n_131), .B1(n_1267), .B2(n_1270), .Y(n_1321) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_88), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_89), .A2(n_113), .B1(n_1260), .B2(n_1264), .Y(n_1259) );
INVx1_ASAP7_75t_L g1218 ( .A(n_90), .Y(n_1218) );
INVx1_ASAP7_75t_L g1150 ( .A(n_91), .Y(n_1150) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_92), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_93), .A2(n_234), .B1(n_646), .B2(n_960), .Y(n_959) );
AOI21xp33_ASAP7_75t_L g991 ( .A1(n_93), .A2(n_328), .B(n_992), .Y(n_991) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_94), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_95), .A2(n_132), .B1(n_687), .B2(n_690), .Y(n_686) );
OAI211xp5_ASAP7_75t_L g702 ( .A1(n_95), .A2(n_387), .B(n_703), .C(n_711), .Y(n_702) );
INVx1_ASAP7_75t_L g377 ( .A(n_97), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_97), .A2(n_191), .B1(n_472), .B2(n_476), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_98), .A2(n_123), .B1(n_378), .B2(n_497), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_98), .A2(n_265), .B1(n_431), .B2(n_823), .C(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g874 ( .A(n_99), .Y(n_874) );
AOI221xp5_ASAP7_75t_L g893 ( .A1(n_99), .A2(n_155), .B1(n_608), .B2(n_894), .C(n_896), .Y(n_893) );
INVx1_ASAP7_75t_L g685 ( .A(n_100), .Y(n_685) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_101), .Y(n_276) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_101), .B(n_274), .Y(n_1261) );
INVx1_ASAP7_75t_L g699 ( .A(n_102), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_103), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_105), .A2(n_166), .B1(n_337), .B2(n_513), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_105), .A2(n_106), .B1(n_462), .B2(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g535 ( .A(n_106), .Y(n_535) );
INVx1_ASAP7_75t_L g1245 ( .A(n_107), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_108), .B(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1269 ( .A(n_108), .Y(n_1269) );
XOR2x2_ASAP7_75t_L g789 ( .A(n_109), .B(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g787 ( .A(n_110), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_111), .A2(n_483), .B1(n_484), .B2(n_574), .Y(n_482) );
INVx1_ASAP7_75t_L g574 ( .A(n_111), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g1285 ( .A1(n_111), .A2(n_178), .B1(n_1267), .B2(n_1270), .Y(n_1285) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_112), .A2(n_260), .B1(n_990), .B2(n_1169), .C(n_1172), .Y(n_1168) );
INVx1_ASAP7_75t_L g1195 ( .A(n_112), .Y(n_1195) );
INVx1_ASAP7_75t_L g697 ( .A(n_114), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_115), .A2(n_146), .B1(n_604), .B2(n_606), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_115), .A2(n_119), .B1(n_631), .B2(n_635), .C(n_637), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_116), .A2(n_226), .B1(n_462), .B2(n_845), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_117), .A2(n_256), .B1(n_516), .B2(n_674), .Y(n_1155) );
INVxp33_ASAP7_75t_L g1200 ( .A(n_117), .Y(n_1200) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_118), .Y(n_588) );
INVx2_ASAP7_75t_L g330 ( .A(n_120), .Y(n_330) );
INVx1_ASAP7_75t_L g342 ( .A(n_120), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_120), .B(n_331), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_121), .Y(n_914) );
INVx1_ASAP7_75t_L g883 ( .A(n_122), .Y(n_883) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_122), .A2(n_163), .B1(n_671), .B2(n_672), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_123), .A2(n_257), .B1(n_826), .B2(n_845), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_124), .A2(n_156), .B1(n_488), .B2(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_125), .A2(n_212), .B1(n_804), .B2(n_808), .Y(n_1121) );
INVxp67_ASAP7_75t_SL g1224 ( .A(n_126), .Y(n_1224) );
OAI221xp5_ASAP7_75t_L g1154 ( .A1(n_127), .A2(n_161), .B1(n_355), .B2(n_671), .C(n_672), .Y(n_1154) );
NOR2xp33_ASAP7_75t_L g1185 ( .A(n_127), .B(n_709), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_129), .A2(n_189), .B1(n_804), .B2(n_806), .Y(n_803) );
AOI21xp33_ASAP7_75t_L g842 ( .A1(n_129), .A2(n_823), .B(n_843), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_130), .A2(n_152), .B1(n_545), .B2(n_1214), .C(n_1220), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1236 ( .A1(n_130), .A2(n_162), .B1(n_314), .B2(n_497), .C(n_1237), .Y(n_1236) );
OAI221xp5_ASAP7_75t_L g876 ( .A1(n_133), .A2(n_163), .B1(n_467), .B2(n_877), .C(n_879), .Y(n_876) );
INVx1_ASAP7_75t_L g853 ( .A(n_134), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_135), .A2(n_240), .B1(n_1267), .B2(n_1270), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_137), .A2(n_140), .B1(n_1260), .B2(n_1264), .Y(n_1320) );
INVx1_ASAP7_75t_L g770 ( .A(n_138), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_138), .A2(n_193), .B1(n_639), .B2(n_640), .Y(n_786) );
INVx1_ASAP7_75t_L g1217 ( .A(n_139), .Y(n_1217) );
AOI221xp5_ASAP7_75t_L g1231 ( .A1(n_139), .A2(n_264), .B1(n_314), .B2(n_1015), .C(n_1232), .Y(n_1231) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_141), .Y(n_435) );
INVxp67_ASAP7_75t_SL g1474 ( .A(n_142), .Y(n_1474) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_143), .A2(n_147), .B1(n_1267), .B2(n_1270), .Y(n_1288) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_144), .Y(n_792) );
OAI211xp5_ASAP7_75t_SL g1475 ( .A1(n_145), .A2(n_1476), .B(n_1477), .C(n_1482), .Y(n_1475) );
INVx1_ASAP7_75t_L g1496 ( .A(n_145), .Y(n_1496) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_148), .A2(n_154), .B1(n_516), .B2(n_674), .Y(n_673) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_148), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_149), .A2(n_674), .B1(n_917), .B2(n_920), .Y(n_916) );
INVx1_ASAP7_75t_L g936 ( .A(n_149), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_150), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g1114 ( .A(n_151), .Y(n_1114) );
INVx1_ASAP7_75t_L g1235 ( .A(n_152), .Y(n_1235) );
INVx1_ASAP7_75t_L g969 ( .A(n_153), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_153), .A2(n_219), .B1(n_911), .B2(n_994), .Y(n_993) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_154), .Y(n_707) );
INVx1_ASAP7_75t_L g860 ( .A(n_155), .Y(n_860) );
OAI211xp5_ASAP7_75t_L g819 ( .A1(n_156), .A2(n_820), .B(n_821), .C(n_827), .Y(n_819) );
INVx1_ASAP7_75t_L g1492 ( .A(n_158), .Y(n_1492) );
BUFx3_ASAP7_75t_L g310 ( .A(n_159), .Y(n_310) );
INVx1_ASAP7_75t_L g1470 ( .A(n_160), .Y(n_1470) );
INVxp67_ASAP7_75t_SL g1180 ( .A(n_161), .Y(n_1180) );
AOI221xp5_ASAP7_75t_L g1212 ( .A1(n_162), .A2(n_209), .B1(n_942), .B2(n_1213), .C(n_1214), .Y(n_1212) );
AOI22xp5_ASAP7_75t_L g1276 ( .A1(n_164), .A2(n_168), .B1(n_1267), .B2(n_1270), .Y(n_1276) );
XNOR2x1_ASAP7_75t_L g1462 ( .A(n_164), .B(n_1463), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_164), .A2(n_1509), .B1(n_1512), .B2(n_1516), .Y(n_1508) );
INVx1_ASAP7_75t_L g798 ( .A(n_165), .Y(n_798) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_166), .A2(n_236), .B1(n_552), .B2(n_554), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_167), .A2(n_170), .B1(n_511), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_167), .A2(n_220), .B1(n_639), .B2(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g679 ( .A(n_169), .Y(n_679) );
OAI21xp5_ASAP7_75t_SL g658 ( .A1(n_171), .A2(n_659), .B(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g974 ( .A(n_172), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g1282 ( .A1(n_173), .A2(n_230), .B1(n_1260), .B2(n_1264), .Y(n_1282) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_174), .Y(n_288) );
INVx1_ASAP7_75t_L g379 ( .A(n_175), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g933 ( .A1(n_176), .A2(n_934), .B(n_935), .C(n_938), .Y(n_933) );
INVx1_ASAP7_75t_L g937 ( .A(n_177), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_179), .Y(n_913) );
INVx1_ASAP7_75t_L g1139 ( .A(n_180), .Y(n_1139) );
INVx1_ASAP7_75t_L g1125 ( .A(n_181), .Y(n_1125) );
OAI21xp5_ASAP7_75t_L g1485 ( .A1(n_182), .A2(n_794), .B(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g956 ( .A(n_183), .Y(n_956) );
INVx1_ASAP7_75t_L g755 ( .A(n_184), .Y(n_755) );
INVx1_ASAP7_75t_L g1068 ( .A(n_185), .Y(n_1068) );
OAI211xp5_ASAP7_75t_L g1080 ( .A1(n_185), .A2(n_1081), .B(n_1083), .C(n_1085), .Y(n_1080) );
INVx1_ASAP7_75t_L g501 ( .A(n_186), .Y(n_501) );
OAI221xp5_ASAP7_75t_L g556 ( .A1(n_186), .A2(n_416), .B1(n_557), .B2(n_565), .C(n_566), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_187), .Y(n_868) );
INVx1_ASAP7_75t_L g923 ( .A(n_188), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_188), .A2(n_194), .B1(n_461), .B2(n_555), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g812 ( .A1(n_190), .A2(n_245), .B1(n_813), .B2(n_817), .Y(n_812) );
INVx1_ASAP7_75t_L g828 ( .A(n_190), .Y(n_828) );
INVx1_ASAP7_75t_L g350 ( .A(n_191), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_192), .Y(n_1011) );
INVx1_ASAP7_75t_L g761 ( .A(n_193), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_194), .A2(n_224), .B1(n_338), .B2(n_911), .C(n_912), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_195), .Y(n_491) );
INVx1_ASAP7_75t_L g721 ( .A(n_196), .Y(n_721) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_197), .Y(n_287) );
INVx1_ASAP7_75t_L g747 ( .A(n_198), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_198), .A2(n_200), .B1(n_472), .B2(n_476), .Y(n_779) );
OAI211xp5_ASAP7_75t_L g1056 ( .A1(n_199), .A2(n_1057), .B(n_1059), .C(n_1062), .Y(n_1056) );
INVx1_ASAP7_75t_L g1093 ( .A(n_199), .Y(n_1093) );
INVx1_ASAP7_75t_L g750 ( .A(n_200), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_201), .Y(n_591) );
INVx1_ASAP7_75t_L g683 ( .A(n_202), .Y(n_683) );
CKINVDCx5p33_ASAP7_75t_R g918 ( .A(n_203), .Y(n_918) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_204), .Y(n_1026) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_206), .Y(n_866) );
INVxp67_ASAP7_75t_SL g881 ( .A(n_207), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_207), .A2(n_674), .B1(n_900), .B2(n_901), .Y(n_899) );
INVx1_ASAP7_75t_L g1233 ( .A(n_209), .Y(n_1233) );
INVx1_ASAP7_75t_L g1223 ( .A(n_210), .Y(n_1223) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_211), .Y(n_1016) );
INVx1_ASAP7_75t_L g1159 ( .A(n_213), .Y(n_1159) );
OAI21xp5_ASAP7_75t_L g977 ( .A1(n_214), .A2(n_978), .B(n_979), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_214), .A2(n_232), .B1(n_516), .B2(n_674), .Y(n_980) );
INVx1_ASAP7_75t_L g840 ( .A(n_215), .Y(n_840) );
OAI211xp5_ASAP7_75t_L g748 ( .A1(n_216), .A2(n_355), .B(n_381), .C(n_749), .Y(n_748) );
INVxp33_ASAP7_75t_SL g778 ( .A(n_216), .Y(n_778) );
INVx1_ASAP7_75t_L g669 ( .A(n_217), .Y(n_669) );
INVx1_ASAP7_75t_L g952 ( .A(n_218), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_219), .A2(n_251), .B1(n_412), .B2(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g486 ( .A(n_221), .Y(n_486) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_222), .Y(n_492) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_222), .A2(n_355), .B1(n_516), .B2(n_519), .C(n_529), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_223), .Y(n_862) );
INVx1_ASAP7_75t_L g1001 ( .A(n_225), .Y(n_1001) );
BUFx3_ASAP7_75t_L g291 ( .A(n_227), .Y(n_291) );
INVx1_ASAP7_75t_L g395 ( .A(n_227), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_228), .Y(n_1013) );
INVx1_ASAP7_75t_L g758 ( .A(n_229), .Y(n_758) );
INVx1_ASAP7_75t_L g480 ( .A(n_231), .Y(n_480) );
INVxp33_ASAP7_75t_L g976 ( .A(n_232), .Y(n_976) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_233), .A2(n_328), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g549 ( .A(n_233), .Y(n_549) );
INVx1_ASAP7_75t_L g983 ( .A(n_234), .Y(n_983) );
XOR2xp5_ASAP7_75t_L g577 ( .A(n_235), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g528 ( .A(n_236), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_237), .Y(n_498) );
INVx1_ASAP7_75t_L g885 ( .A(n_239), .Y(n_885) );
INVx2_ASAP7_75t_L g385 ( .A(n_241), .Y(n_385) );
INVx1_ASAP7_75t_L g392 ( .A(n_241), .Y(n_392) );
INVx1_ASAP7_75t_L g405 ( .A(n_241), .Y(n_405) );
INVxp67_ASAP7_75t_SL g1225 ( .A(n_242), .Y(n_1225) );
AOI221xp5_ASAP7_75t_L g984 ( .A1(n_243), .A2(n_251), .B1(n_339), .B2(n_616), .C(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1113 ( .A(n_244), .Y(n_1113) );
INVx1_ASAP7_75t_L g829 ( .A(n_245), .Y(n_829) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_246), .Y(n_710) );
INVx1_ASAP7_75t_L g906 ( .A(n_247), .Y(n_906) );
INVx1_ASAP7_75t_L g925 ( .A(n_248), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_250), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_252), .B(n_570), .Y(n_569) );
XNOR2xp5_ASAP7_75t_L g1513 ( .A(n_253), .B(n_1514), .Y(n_1513) );
OAI21xp33_ASAP7_75t_SL g742 ( .A1(n_255), .A2(n_387), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g746 ( .A(n_255), .Y(n_746) );
INVxp67_ASAP7_75t_SL g1175 ( .A(n_256), .Y(n_1175) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_257), .A2(n_265), .B1(n_378), .B2(n_497), .Y(n_811) );
NAND2xp33_ASAP7_75t_SL g1211 ( .A(n_258), .B(n_452), .Y(n_1211) );
INVx1_ASAP7_75t_L g1238 ( .A(n_258), .Y(n_1238) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_259), .A2(n_263), .B1(n_367), .B2(n_368), .C(n_373), .Y(n_366) );
INVx1_ASAP7_75t_L g500 ( .A(n_261), .Y(n_500) );
INVx1_ASAP7_75t_L g1483 ( .A(n_262), .Y(n_1483) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_263), .Y(n_420) );
INVx1_ASAP7_75t_L g1209 ( .A(n_264), .Y(n_1209) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_292), .B(n_1248), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_277), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g1507 ( .A(n_271), .B(n_280), .Y(n_1507) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g1511 ( .A(n_273), .B(n_276), .Y(n_1511) );
INVx1_ASAP7_75t_L g1519 ( .A(n_273), .Y(n_1519) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g1521 ( .A(n_276), .B(n_1519), .Y(n_1521) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g1070 ( .A(n_280), .B(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g445 ( .A(n_281), .B(n_291), .Y(n_445) );
AND2x4_ASAP7_75t_L g651 ( .A(n_281), .B(n_290), .Y(n_651) );
AND2x4_ASAP7_75t_SL g1506 ( .A(n_282), .B(n_1507), .Y(n_1506) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_284), .B(n_289), .Y(n_283) );
BUFx4f_ASAP7_75t_L g861 ( .A(n_284), .Y(n_861) );
INVxp67_ASAP7_75t_L g873 ( .A(n_284), .Y(n_873) );
INVx1_ASAP7_75t_L g971 ( .A(n_284), .Y(n_971) );
OR2x6_ASAP7_75t_L g1049 ( .A(n_284), .B(n_1045), .Y(n_1049) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx4f_ASAP7_75t_L g437 ( .A(n_285), .Y(n_437) );
INVx3_ASAP7_75t_L g735 ( .A(n_285), .Y(n_735) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g397 ( .A(n_287), .Y(n_397) );
INVx2_ASAP7_75t_L g415 ( .A(n_287), .Y(n_415) );
NAND2x1_ASAP7_75t_L g418 ( .A(n_287), .B(n_288), .Y(n_418) );
AND2x2_ASAP7_75t_L g425 ( .A(n_287), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g433 ( .A(n_287), .B(n_288), .Y(n_433) );
INVx1_ASAP7_75t_L g479 ( .A(n_287), .Y(n_479) );
INVx1_ASAP7_75t_L g398 ( .A(n_288), .Y(n_398) );
AND2x2_ASAP7_75t_L g414 ( .A(n_288), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g426 ( .A(n_288), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_288), .B(n_415), .Y(n_443) );
OR2x2_ASAP7_75t_L g454 ( .A(n_288), .B(n_397), .Y(n_454) );
BUFx2_ASAP7_75t_L g475 ( .A(n_288), .Y(n_475) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g1061 ( .A(n_290), .Y(n_1061) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_L g1055 ( .A(n_291), .Y(n_1055) );
AND2x4_ASAP7_75t_L g1067 ( .A(n_291), .B(n_478), .Y(n_1067) );
OAI22xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B1(n_1106), .B2(n_1107), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
XNOR2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_848), .Y(n_294) );
XOR2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_575), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
XNOR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_482), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_480), .B(n_481), .Y(n_299) );
AND3x1_ASAP7_75t_L g300 ( .A(n_301), .B(n_399), .C(n_427), .Y(n_300) );
AOI31xp33_ASAP7_75t_L g481 ( .A1(n_301), .A2(n_399), .A3(n_427), .B(n_480), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_382), .B(n_386), .Y(n_301) );
NAND3xp33_ASAP7_75t_SL g302 ( .A(n_303), .B(n_344), .C(n_360), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_320), .B1(n_332), .B2(n_335), .Y(n_303) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g605 ( .A(n_307), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_307), .B(n_929), .Y(n_928) );
BUFx3_ASAP7_75t_L g994 ( .A(n_307), .Y(n_994) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
INVx8_ASAP7_75t_L g376 ( .A(n_308), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g381 ( .A(n_308), .B(n_348), .Y(n_381) );
AND2x2_ASAP7_75t_L g688 ( .A(n_308), .B(n_689), .Y(n_688) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_308), .Y(n_1119) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
AND2x4_ASAP7_75t_L g326 ( .A(n_309), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_310), .Y(n_316) );
AND2x4_ASAP7_75t_L g322 ( .A(n_310), .B(n_318), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_310), .B(n_319), .Y(n_372) );
OR2x2_ASAP7_75t_L g527 ( .A(n_310), .B(n_312), .Y(n_527) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_L g327 ( .A(n_313), .Y(n_327) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx5_ASAP7_75t_L g514 ( .A(n_315), .Y(n_514) );
AND2x4_ASAP7_75t_L g573 ( .A(n_315), .B(n_364), .Y(n_573) );
BUFx3_ASAP7_75t_L g608 ( .A(n_315), .Y(n_608) );
BUFx3_ASAP7_75t_L g610 ( .A(n_315), .Y(n_610) );
BUFx12f_ASAP7_75t_L g911 ( .A(n_315), .Y(n_911) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_316), .B(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g1089 ( .A(n_316), .Y(n_1089) );
INVx1_ASAP7_75t_L g352 ( .A(n_317), .Y(n_352) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g358 ( .A(n_319), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_321), .A2(n_491), .B1(n_497), .B2(n_498), .Y(n_496) );
BUFx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g336 ( .A(n_322), .Y(n_336) );
BUFx2_ASAP7_75t_L g378 ( .A(n_322), .Y(n_378) );
BUFx2_ASAP7_75t_L g606 ( .A(n_322), .Y(n_606) );
BUFx2_ASAP7_75t_L g619 ( .A(n_322), .Y(n_619) );
AND2x2_ASAP7_75t_L g691 ( .A(n_322), .B(n_689), .Y(n_691) );
INVx2_ASAP7_75t_L g986 ( .A(n_322), .Y(n_986) );
AND2x4_ASAP7_75t_L g1084 ( .A(n_322), .B(n_343), .Y(n_1084) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_SL g334 ( .A(n_325), .Y(n_334) );
INVx3_ASAP7_75t_L g367 ( .A(n_325), .Y(n_367) );
INVx5_ASAP7_75t_L g805 ( .A(n_325), .Y(n_805) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx8_ASAP7_75t_L g511 ( .A(n_326), .Y(n_511) );
INVx2_ASAP7_75t_L g518 ( .A(n_326), .Y(n_518) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_326), .Y(n_695) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g1008 ( .A(n_329), .B(n_448), .Y(n_1008) );
NAND2xp33_ASAP7_75t_SL g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g349 ( .A(n_330), .Y(n_349) );
AND3x4_ASAP7_75t_L g601 ( .A(n_330), .B(n_539), .C(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g680 ( .A(n_330), .B(n_602), .Y(n_680) );
HB1xp67_ASAP7_75t_L g1102 ( .A(n_330), .Y(n_1102) );
INVx3_ASAP7_75t_L g343 ( .A(n_331), .Y(n_343) );
BUFx3_ASAP7_75t_L g602 ( .A(n_331), .Y(n_602) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g895 ( .A(n_338), .Y(n_895) );
INVx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_340), .A2(n_520), .B1(n_523), .B2(n_524), .C(n_528), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_340), .A2(n_522), .B1(n_697), .B2(n_698), .C(n_699), .Y(n_696) );
OAI221xp5_ASAP7_75t_L g763 ( .A1(n_340), .A2(n_698), .B1(n_764), .B2(n_765), .C(n_767), .Y(n_763) );
OAI221xp5_ASAP7_75t_L g900 ( .A1(n_340), .A2(n_522), .B1(n_698), .B2(n_862), .C(n_870), .Y(n_900) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_340), .A2(n_356), .B1(n_526), .B2(n_918), .C(n_919), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_340), .B(n_1173), .Y(n_1172) );
OAI221xp5_ASAP7_75t_L g1232 ( .A1(n_340), .A2(n_524), .B1(n_1233), .B2(n_1234), .C(n_1235), .Y(n_1232) );
INVx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x6_ASAP7_75t_L g810 ( .A(n_341), .B(n_384), .Y(n_810) );
NAND2x1p5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND3x1_ASAP7_75t_L g613 ( .A(n_342), .B(n_343), .C(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_L g348 ( .A(n_343), .B(n_349), .Y(n_348) );
OR2x4_ASAP7_75t_L g1076 ( .A(n_343), .B(n_527), .Y(n_1076) );
INVx1_ASAP7_75t_L g1079 ( .A(n_343), .Y(n_1079) );
OR2x6_ASAP7_75t_L g1099 ( .A(n_343), .B(n_371), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_350), .B1(n_351), .B2(n_353), .C(n_354), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_345), .A2(n_351), .B1(n_500), .B2(n_501), .Y(n_499) );
INVx4_ASAP7_75t_L g671 ( .A(n_345), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_345), .A2(n_351), .B1(n_750), .B2(n_751), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_345), .A2(n_351), .B1(n_956), .B2(n_974), .Y(n_998) );
AND2x6_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
NAND2x1_ASAP7_75t_L g593 ( .A(n_346), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g799 ( .A(n_346), .B(n_594), .Y(n_799) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g351 ( .A(n_348), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g359 ( .A(n_348), .Y(n_359) );
AND2x4_ASAP7_75t_L g594 ( .A(n_348), .B(n_404), .Y(n_594) );
INVx2_ASAP7_75t_L g672 ( .A(n_351), .Y(n_672) );
INVx1_ASAP7_75t_L g598 ( .A(n_352), .Y(n_598) );
NOR3xp33_ASAP7_75t_L g892 ( .A(n_354), .B(n_893), .C(n_899), .Y(n_892) );
NOR3xp33_ASAP7_75t_L g909 ( .A(n_354), .B(n_910), .C(n_916), .Y(n_909) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_355), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
INVx1_ASAP7_75t_L g990 ( .A(n_356), .Y(n_990) );
INVx1_ASAP7_75t_L g1082 ( .A(n_356), .Y(n_1082) );
BUFx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_357), .Y(n_507) );
BUFx3_ASAP7_75t_L g522 ( .A(n_357), .Y(n_522) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_358), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_366), .B1(n_379), .B2(n_380), .Y(n_360) );
INVxp67_ASAP7_75t_L g495 ( .A(n_361), .Y(n_495) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g890 ( .A(n_363), .Y(n_890) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g517 ( .A(n_364), .Y(n_517) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g587 ( .A(n_365), .B(n_448), .Y(n_587) );
INVx1_ASAP7_75t_L g689 ( .A(n_365), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_367), .A2(n_921), .B1(n_922), .B2(n_923), .Y(n_920) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g1020 ( .A(n_371), .Y(n_1020) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g534 ( .A(n_372), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_377), .B2(n_378), .Y(n_373) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx8_ASAP7_75t_L g497 ( .A(n_376), .Y(n_497) );
INVx2_ASAP7_75t_L g616 ( .A(n_376), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_380), .A2(n_669), .B(n_670), .C(n_673), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g887 ( .A1(n_380), .A2(n_882), .B1(n_888), .B2(n_890), .C(n_891), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_380), .A2(n_890), .B1(n_925), .B2(n_926), .C(n_930), .Y(n_924) );
INVx2_ASAP7_75t_L g997 ( .A(n_380), .Y(n_997) );
AOI211xp5_ASAP7_75t_SL g1152 ( .A1(n_380), .A2(n_1153), .B(n_1154), .C(n_1155), .Y(n_1152) );
AOI211xp5_ASAP7_75t_SL g1227 ( .A1(n_380), .A2(n_1223), .B(n_1228), .C(n_1229), .Y(n_1227) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g488 ( .A(n_381), .B(n_489), .Y(n_488) );
OR2x6_ASAP7_75t_L g581 ( .A(n_381), .B(n_489), .Y(n_581) );
INVx1_ASAP7_75t_L g657 ( .A(n_382), .Y(n_657) );
INVx2_ASAP7_75t_L g701 ( .A(n_382), .Y(n_701) );
BUFx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_383), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g1000 ( .A(n_383), .Y(n_1000) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g465 ( .A(n_384), .B(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_385), .B(n_407), .Y(n_470) );
INVx2_ASAP7_75t_L g539 ( .A(n_385), .Y(n_539) );
INVx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI222xp33_ASAP7_75t_L g485 ( .A1(n_388), .A2(n_422), .B1(n_486), .B2(n_487), .C1(n_491), .C2(n_492), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_388), .B(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_388), .B(n_929), .Y(n_932) );
AOI211x1_ASAP7_75t_L g951 ( .A1(n_388), .A2(n_952), .B(n_953), .C(n_977), .Y(n_951) );
AO211x2_ASAP7_75t_L g1149 ( .A1(n_388), .A2(n_1150), .B(n_1151), .C(n_1176), .Y(n_1149) );
AND2x4_ASAP7_75t_L g388 ( .A(n_389), .B(n_393), .Y(n_388) );
AND2x4_ASAP7_75t_L g422 ( .A(n_389), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g476 ( .A(n_390), .B(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_L g489 ( .A(n_390), .Y(n_489) );
OR2x2_ASAP7_75t_L g879 ( .A(n_390), .B(n_477), .Y(n_879) );
INVx1_ASAP7_75t_L g1071 ( .A(n_390), .Y(n_1071) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g448 ( .A(n_391), .Y(n_448) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_393), .Y(n_624) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_394), .B(n_405), .Y(n_411) );
AND2x2_ASAP7_75t_L g423 ( .A(n_394), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g627 ( .A(n_394), .B(n_424), .Y(n_627) );
AND2x4_ASAP7_75t_L g629 ( .A(n_394), .B(n_555), .Y(n_629) );
AND2x4_ASAP7_75t_SL g644 ( .A(n_394), .B(n_432), .Y(n_644) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_395), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_396), .B(n_407), .Y(n_406) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_396), .Y(n_461) );
INVx3_ASAP7_75t_L g553 ( .A(n_396), .Y(n_553) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_419), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_403), .B(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g584 ( .A(n_403), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g705 ( .A(n_404), .Y(n_705) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g614 ( .A(n_405), .Y(n_614) );
INVx1_ASAP7_75t_L g706 ( .A(n_406), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_407), .B(n_478), .Y(n_477) );
AND2x6_ASAP7_75t_L g641 ( .A(n_407), .B(n_432), .Y(n_641) );
AND2x2_ASAP7_75t_L g655 ( .A(n_407), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g838 ( .A(n_407), .Y(n_838) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g490 ( .A(n_409), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g703 ( .A1(n_409), .A2(n_669), .B1(n_704), .B2(n_707), .C1(n_708), .C2(n_710), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g777 ( .A1(n_409), .A2(n_778), .B(n_779), .Y(n_777) );
AOI222xp33_ASAP7_75t_L g880 ( .A1(n_409), .A2(n_704), .B1(n_708), .B2(n_881), .C1(n_882), .C2(n_883), .Y(n_880) );
AOI222xp33_ASAP7_75t_L g954 ( .A1(n_409), .A2(n_567), .B1(n_568), .B2(n_955), .C1(n_956), .C2(n_957), .Y(n_954) );
INVx1_ASAP7_75t_L g1179 ( .A(n_409), .Y(n_1179) );
AOI222xp33_ASAP7_75t_L g1222 ( .A1(n_409), .A2(n_704), .B1(n_708), .B2(n_1223), .C1(n_1224), .C2(n_1225), .Y(n_1222) );
AND2x4_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
AOI332xp33_ASAP7_75t_L g935 ( .A1(n_410), .A2(n_412), .A3(n_705), .B1(n_706), .B2(n_708), .B3(n_925), .C1(n_936), .C2(n_937), .Y(n_935) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g416 ( .A(n_411), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g709 ( .A(n_411), .B(n_417), .Y(n_709) );
INVx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_414), .Y(n_555) );
BUFx3_ASAP7_75t_L g640 ( .A(n_414), .Y(n_640) );
BUFx3_ASAP7_75t_L g869 ( .A(n_417), .Y(n_869) );
INVx2_ASAP7_75t_SL g1036 ( .A(n_417), .Y(n_1036) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_418), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_421), .B(n_1244), .Y(n_1243) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_422), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_422), .B(n_776), .Y(n_775) );
NAND2xp33_ASAP7_75t_SL g902 ( .A(n_422), .B(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g934 ( .A(n_422), .Y(n_934) );
INVx1_ASAP7_75t_L g978 ( .A(n_422), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_422), .B(n_1175), .Y(n_1174) );
BUFx6f_ASAP7_75t_L g782 ( .A(n_424), .Y(n_782) );
INVx2_ASAP7_75t_L g1192 ( .A(n_424), .Y(n_1192) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g430 ( .A(n_425), .Y(n_430) );
BUFx3_ASAP7_75t_L g636 ( .A(n_425), .Y(n_636) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_425), .B(n_1045), .Y(n_1044) );
AOI211xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_444), .B(n_449), .C(n_471), .Y(n_427) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g648 ( .A(n_430), .Y(n_648) );
BUFx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx3_ASAP7_75t_L g649 ( .A(n_432), .Y(n_649) );
BUFx3_ASAP7_75t_L g785 ( .A(n_432), .Y(n_785) );
INVx1_ASAP7_75t_L g967 ( .A(n_432), .Y(n_967) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_432), .B(n_1061), .Y(n_1060) );
BUFx6f_ASAP7_75t_L g1131 ( .A(n_432), .Y(n_1131) );
BUFx3_ASAP7_75t_L g1135 ( .A(n_432), .Y(n_1135) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g634 ( .A(n_433), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_438), .B2(n_439), .Y(n_434) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_437), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_439), .A2(n_1010), .B1(n_1024), .B2(n_1030), .Y(n_1029) );
INVx6_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx5_ASAP7_75t_L g1196 ( .A(n_440), .Y(n_1196) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g725 ( .A(n_441), .Y(n_725) );
INVx2_ASAP7_75t_SL g736 ( .A(n_441), .Y(n_736) );
INVx4_ASAP7_75t_L g973 ( .A(n_441), .Y(n_973) );
INVx1_ASAP7_75t_L g1040 ( .A(n_441), .Y(n_1040) );
INVx2_ASAP7_75t_L g1221 ( .A(n_441), .Y(n_1221) );
INVx8_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_442), .B(n_1055), .Y(n_1054) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_444), .Y(n_565) );
AOI332xp33_ASAP7_75t_L g780 ( .A1(n_444), .A2(n_544), .A3(n_704), .B1(n_781), .B2(n_783), .B3(n_784), .C1(n_786), .C2(n_787), .Y(n_780) );
AOI322xp5_ASAP7_75t_L g958 ( .A1(n_444), .A2(n_708), .A3(n_959), .B1(n_962), .B2(n_964), .C1(n_965), .C2(n_974), .Y(n_958) );
INVx2_ASAP7_75t_L g1037 ( .A(n_444), .Y(n_1037) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx4_ASAP7_75t_L g637 ( .A(n_445), .Y(n_637) );
AND2x2_ASAP7_75t_SL g732 ( .A(n_445), .B(n_448), .Y(n_732) );
INVx1_ASAP7_75t_SL g824 ( .A(n_445), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_445), .B(n_446), .Y(n_942) );
INVx4_ASAP7_75t_L g1480 ( .A(n_445), .Y(n_1480) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_448), .Y(n_1104) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_463), .B(n_467), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_455), .B1(n_456), .B2(n_459), .C(n_460), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g1216 ( .A1(n_451), .A2(n_550), .B1(n_1217), .B2(n_1218), .C(n_1219), .Y(n_1216) );
OAI221xp5_ASAP7_75t_L g1468 ( .A1(n_451), .A2(n_651), .B1(n_1469), .B2(n_1470), .C(n_1471), .Y(n_1468) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g940 ( .A1(n_453), .A2(n_550), .B1(n_914), .B2(n_921), .C(n_941), .Y(n_940) );
BUFx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g548 ( .A(n_454), .Y(n_548) );
BUFx2_ASAP7_75t_L g560 ( .A(n_454), .Y(n_560) );
INVx1_ASAP7_75t_L g1213 ( .A(n_456), .Y(n_1213) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g730 ( .A(n_457), .Y(n_730) );
INVx2_ASAP7_75t_L g841 ( .A(n_457), .Y(n_841) );
INVx4_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x6_ASAP7_75t_L g467 ( .A(n_458), .B(n_468), .Y(n_467) );
BUFx4f_ASAP7_75t_L g550 ( .A(n_458), .Y(n_550) );
BUFx4f_ASAP7_75t_L g561 ( .A(n_458), .Y(n_561) );
BUFx4f_ASAP7_75t_L g720 ( .A(n_458), .Y(n_720) );
BUFx6f_ASAP7_75t_L g945 ( .A(n_458), .Y(n_945) );
BUFx4f_ASAP7_75t_L g1469 ( .A(n_458), .Y(n_1469) );
INVx3_ASAP7_75t_L g564 ( .A(n_461), .Y(n_564) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_461), .Y(n_845) );
INVx1_ASAP7_75t_L g964 ( .A(n_463), .Y(n_964) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx4_ASAP7_75t_L g545 ( .A(n_465), .Y(n_545) );
INVx2_ASAP7_75t_L g717 ( .A(n_465), .Y(n_717) );
INVx2_ASAP7_75t_L g858 ( .A(n_465), .Y(n_858) );
INVx1_ASAP7_75t_L g1028 ( .A(n_465), .Y(n_1028) );
OAI21xp5_ASAP7_75t_SL g541 ( .A1(n_467), .A2(n_542), .B(n_546), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_467), .Y(n_714) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2x2_ASAP7_75t_L g472 ( .A(n_469), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g567 ( .A(n_472), .Y(n_567) );
INVx2_ASAP7_75t_SL g878 ( .A(n_472), .Y(n_878) );
INVx2_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g656 ( .A(n_475), .Y(n_656) );
INVx1_ASAP7_75t_L g837 ( .A(n_475), .Y(n_837) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_475), .B(n_1055), .Y(n_1063) );
INVx2_ASAP7_75t_SL g568 ( .A(n_476), .Y(n_568) );
AND2x4_ASAP7_75t_L g659 ( .A(n_476), .B(n_660), .Y(n_659) );
AND2x4_ASAP7_75t_L g794 ( .A(n_476), .B(n_660), .Y(n_794) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .C(n_540), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_515), .B(n_536), .Y(n_493) );
OAI211xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_499), .C(n_502), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_498), .A2(n_500), .B1(n_567), .B2(n_568), .Y(n_566) );
OAI211xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_508), .C(n_512), .Y(n_502) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_503), .A2(n_523), .B1(n_558), .B2(n_561), .C(n_562), .Y(n_557) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g889 ( .A(n_506), .Y(n_889) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g660 ( .A(n_507), .B(n_587), .Y(n_660) );
BUFx6f_ASAP7_75t_L g754 ( .A(n_507), .Y(n_754) );
INVx4_ASAP7_75t_L g766 ( .A(n_507), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g912 ( .A1(n_507), .A2(n_680), .B1(n_913), .B2(n_914), .C(n_915), .Y(n_912) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_507), .Y(n_1025) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_510), .A2(n_762), .B1(n_864), .B2(n_875), .Y(n_901) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_SL g530 ( .A(n_511), .Y(n_530) );
AND2x4_ASAP7_75t_L g664 ( .A(n_511), .B(n_663), .Y(n_664) );
INVx3_ASAP7_75t_L g678 ( .A(n_511), .Y(n_678) );
INVx2_ASAP7_75t_SL g1239 ( .A(n_511), .Y(n_1239) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g806 ( .A(n_514), .Y(n_806) );
INVx2_ASAP7_75t_R g808 ( .A(n_514), .Y(n_808) );
OR2x6_ASAP7_75t_SL g516 ( .A(n_517), .B(n_518), .Y(n_516) );
INVx3_ASAP7_75t_L g898 ( .A(n_518), .Y(n_898) );
OAI22xp33_ASAP7_75t_L g1009 ( .A1(n_520), .A2(n_682), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g896 ( .A1(n_522), .A2(n_680), .B1(n_866), .B2(n_868), .C(n_897), .Y(n_896) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx4f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g682 ( .A(n_527), .Y(n_682) );
BUFx3_ASAP7_75t_L g698 ( .A(n_527), .Y(n_698) );
INVx2_ASAP7_75t_L g760 ( .A(n_527), .Y(n_760) );
OR2x4_ASAP7_75t_L g1096 ( .A(n_527), .B(n_1079), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_532), .B2(n_535), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g546 ( .A1(n_531), .A2(n_547), .B1(n_549), .B2(n_550), .C(n_551), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g982 ( .A1(n_532), .A2(n_927), .B1(n_972), .B2(n_983), .C(n_984), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_532), .A2(n_1013), .B1(n_1014), .B2(n_1016), .Y(n_1012) );
CKINVDCx8_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g684 ( .A(n_533), .Y(n_684) );
INVx3_ASAP7_75t_L g762 ( .A(n_533), .Y(n_762) );
INVx3_ASAP7_75t_L g922 ( .A(n_533), .Y(n_922) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g586 ( .A(n_534), .Y(n_586) );
INVx1_ASAP7_75t_L g846 ( .A(n_536), .Y(n_846) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g1242 ( .A(n_537), .Y(n_1242) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_538), .Y(n_931) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI31xp33_ASAP7_75t_SL g743 ( .A1(n_539), .A2(n_744), .A3(n_748), .B(n_752), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_556), .C(n_569), .Y(n_540) );
INVxp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g1187 ( .A(n_545), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_547), .A2(n_550), .B1(n_1013), .B2(n_1018), .Y(n_1031) );
INVx1_ASAP7_75t_L g1034 ( .A(n_547), .Y(n_1034) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g728 ( .A(n_548), .Y(n_728) );
INVx2_ASAP7_75t_L g944 ( .A(n_548), .Y(n_944) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g639 ( .A(n_553), .Y(n_639) );
INVx2_ASAP7_75t_L g963 ( .A(n_553), .Y(n_963) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_555), .Y(n_826) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g719 ( .A(n_559), .Y(n_719) );
INVx4_ASAP7_75t_L g865 ( .A(n_559), .Y(n_865) );
INVx4_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g1137 ( .A(n_564), .Y(n_1137) );
AOI222xp33_ASAP7_75t_L g1177 ( .A1(n_567), .A2(n_568), .B1(n_1153), .B2(n_1178), .C1(n_1180), .C2(n_1181), .Y(n_1177) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx3_ASAP7_75t_L g674 ( .A(n_573), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_738), .B1(n_739), .B2(n_847), .Y(n_575) );
INVx1_ASAP7_75t_L g847 ( .A(n_576), .Y(n_847) );
XNOR2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_665), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_620), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_582), .B1(n_583), .B2(n_588), .C(n_589), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g1112 ( .A1(n_580), .A2(n_583), .B1(n_1113), .B2(n_1114), .C(n_1115), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_580), .B(n_1496), .Y(n_1495) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_582), .A2(n_629), .B1(n_630), .B2(n_638), .C(n_641), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g791 ( .A1(n_583), .A2(n_792), .B(n_793), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_583), .B(n_1489), .Y(n_1488) );
INVx8_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g772 ( .A(n_586), .Y(n_772) );
INVx1_ASAP7_75t_L g663 ( .A(n_587), .Y(n_663) );
INVx1_ASAP7_75t_L g816 ( .A(n_587), .Y(n_816) );
NAND3xp33_ASAP7_75t_SL g589 ( .A(n_590), .B(n_599), .C(n_617), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_595), .B2(n_596), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g642 ( .A1(n_591), .A2(n_595), .B1(n_643), .B2(n_645), .C1(n_652), .C2(n_653), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g1491 ( .A1(n_592), .A2(n_1492), .B1(n_1493), .B2(n_1494), .Y(n_1491) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g596 ( .A(n_594), .B(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g618 ( .A(n_594), .B(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_SL g1494 ( .A(n_594), .B(n_597), .Y(n_1494) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_596), .A2(n_798), .B1(n_799), .B2(n_800), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_596), .A2(n_799), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AOI33xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .A3(n_607), .B1(n_609), .B2(n_611), .B3(n_615), .Y(n_599) );
BUFx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI33xp33_ASAP7_75t_L g801 ( .A1(n_601), .A2(n_802), .A3(n_803), .B1(n_807), .B2(n_809), .B3(n_811), .Y(n_801) );
AOI33xp33_ASAP7_75t_L g1117 ( .A1(n_601), .A2(n_809), .A3(n_1118), .B1(n_1121), .B2(n_1122), .B3(n_1123), .Y(n_1117) );
AOI33xp33_ASAP7_75t_L g1497 ( .A1(n_601), .A2(n_1498), .A3(n_1499), .B1(n_1500), .B2(n_1502), .B3(n_1503), .Y(n_1497) );
INVx3_ASAP7_75t_L g1088 ( .A(n_602), .Y(n_1088) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx2_ASAP7_75t_L g1503 ( .A(n_612), .Y(n_1503) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx3_ASAP7_75t_L g1022 ( .A(n_613), .Y(n_1022) );
AND2x4_ASAP7_75t_L g662 ( .A(n_616), .B(n_663), .Y(n_662) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_616), .B(n_663), .Y(n_1143) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_618), .B(n_796), .C(n_812), .Y(n_795) );
INVx3_ASAP7_75t_L g1116 ( .A(n_618), .Y(n_1116) );
AOI21xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_657), .B(n_658), .Y(n_620) );
NAND3xp33_ASAP7_75t_SL g621 ( .A(n_622), .B(n_628), .C(n_642), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_625), .B2(n_626), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_623), .A2(n_625), .B1(n_662), .B2(n_664), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_624), .A2(n_627), .B1(n_828), .B2(n_829), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_624), .A2(n_627), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_624), .A2(n_627), .B1(n_1483), .B2(n_1484), .Y(n_1482) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_SL g820 ( .A(n_629), .Y(n_820) );
AOI221xp5_ASAP7_75t_L g1133 ( .A1(n_629), .A2(n_641), .B1(n_1113), .B2(n_1134), .C(n_1136), .Y(n_1133) );
INVx3_ASAP7_75t_L g1476 ( .A(n_629), .Y(n_1476) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx2_ASAP7_75t_L g961 ( .A(n_634), .Y(n_961) );
BUFx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_641), .A2(n_822), .B(n_825), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g1477 ( .A1(n_641), .A2(n_1478), .B(n_1481), .Y(n_1477) );
AOI222xp33_ASAP7_75t_L g1129 ( .A1(n_643), .A2(n_655), .B1(n_1125), .B2(n_1126), .C1(n_1130), .C2(n_1132), .Y(n_1129) );
BUFx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g833 ( .A(n_644), .Y(n_833) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g823 ( .A(n_647), .Y(n_823) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx3_ASAP7_75t_L g843 ( .A(n_651), .Y(n_843) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_SL g1465 ( .A1(n_657), .A2(n_1466), .B(n_1475), .C(n_1485), .Y(n_1465) );
INVx2_ASAP7_75t_L g817 ( .A(n_664), .Y(n_817) );
AOI211x1_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_700), .B(n_702), .C(n_713), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_675), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_686), .C(n_692), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B(n_680), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g753 ( .A1(n_678), .A2(n_680), .B1(n_754), .B2(n_755), .C(n_756), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_678), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
INVx1_ASAP7_75t_L g1501 ( .A(n_678), .Y(n_1501) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_679), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g1165 ( .A(n_680), .Y(n_1165) );
OAI221xp5_ASAP7_75t_L g1237 ( .A1(n_680), .A2(n_1218), .B1(n_1234), .B2(n_1238), .C(n_1239), .Y(n_1237) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_682), .A2(n_1024), .B1(n_1025), .B2(n_1026), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_683), .A2(n_699), .B1(n_723), .B2(n_725), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_685), .A2(n_734), .B1(n_736), .B2(n_737), .Y(n_733) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_688), .A2(n_691), .B1(n_746), .B2(n_747), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_688), .A2(n_691), .B1(n_952), .B2(n_957), .Y(n_995) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g915 ( .A(n_695), .Y(n_915) );
BUFx6f_ASAP7_75t_L g992 ( .A(n_695), .Y(n_992) );
BUFx6f_ASAP7_75t_L g1015 ( .A(n_695), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1078 ( .A(n_695), .B(n_1079), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_697), .A2(n_727), .B1(n_729), .B2(n_730), .Y(n_726) );
INVx1_ASAP7_75t_L g1171 ( .A(n_698), .Y(n_1171) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g886 ( .A1(n_701), .A2(n_887), .B(n_892), .C(n_902), .Y(n_886) );
AOI21xp33_ASAP7_75t_L g975 ( .A1(n_704), .A2(n_714), .B(n_976), .Y(n_975) );
AOI21xp33_ASAP7_75t_L g1199 ( .A1(n_704), .A2(n_714), .B(n_1200), .Y(n_1199) );
AND2x4_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_708), .A2(n_714), .B(n_751), .Y(n_774) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR3x1_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .C(n_716), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g938 ( .A(n_714), .B(n_939), .C(n_947), .Y(n_938) );
NOR3xp33_ASAP7_75t_L g1205 ( .A(n_714), .B(n_1206), .C(n_1207), .Y(n_1205) );
OAI33xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .A3(n_722), .B1(n_726), .B2(n_731), .B3(n_733), .Y(n_716) );
INVx1_ASAP7_75t_L g1058 ( .A(n_720), .Y(n_1058) );
INVx3_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g1030 ( .A(n_724), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_727), .A2(n_868), .B1(n_869), .B2(n_870), .Y(n_867) );
INVx4_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI33xp33_ASAP7_75t_L g857 ( .A1(n_731), .A2(n_858), .A3(n_859), .B1(n_863), .B2(n_867), .B3(n_871), .Y(n_857) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx6f_ASAP7_75t_L g1215 ( .A(n_735), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_736), .A2(n_860), .B1(n_861), .B2(n_862), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_736), .A2(n_872), .B1(n_874), .B2(n_875), .Y(n_871) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
XNOR2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_789), .Y(n_739) );
XOR2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_788), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_773), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_757), .B1(n_763), .B2(n_768), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B1(n_761), .B2(n_762), .Y(n_757) );
INVx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_SL g814 ( .A(n_760), .Y(n_814) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g1234 ( .A(n_766), .Y(n_1234) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND4xp25_ASAP7_75t_SL g773 ( .A(n_774), .B(n_775), .C(n_777), .D(n_780), .Y(n_773) );
NAND3xp33_ASAP7_75t_SL g790 ( .A(n_791), .B(n_795), .C(n_818), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_801), .Y(n_796) );
INVx8_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
OR2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVxp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_816), .B(n_898), .Y(n_1144) );
OAI21xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_830), .B(n_846), .Y(n_818) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g1467 ( .A(n_832), .Y(n_1467) );
INVx4_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
BUFx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NOR2x1_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
OAI211xp5_ASAP7_75t_SL g839 ( .A1(n_840), .A2(n_841), .B(n_842), .C(n_844), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_841), .A2(n_864), .B1(n_865), .B2(n_866), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g1127 ( .A1(n_846), .A2(n_1128), .B(n_1141), .Y(n_1127) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
XNOR2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_948), .Y(n_849) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
XNOR2x1_ASAP7_75t_L g851 ( .A(n_852), .B(n_904), .Y(n_851) );
XNOR2x1_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .Y(n_852) );
NOR2x1_ASAP7_75t_L g854 ( .A(n_855), .B(n_886), .Y(n_854) );
NAND3xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_880), .C(n_884), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_876), .Y(n_856) );
OAI22xp5_ASAP7_75t_SL g939 ( .A1(n_858), .A2(n_940), .B1(n_942), .B2(n_943), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_861), .A2(n_1194), .B1(n_1195), .B2(n_1196), .Y(n_1193) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_897), .A2(n_1018), .B1(n_1019), .B2(n_1020), .Y(n_1017) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g927 ( .A(n_898), .Y(n_927) );
INVx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
XNOR2x1_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
OR2x2_ASAP7_75t_L g907 ( .A(n_908), .B(n_933), .Y(n_907) );
A2O1A1Ixp33_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_924), .B(n_931), .C(n_932), .Y(n_908) );
OAI221xp5_ASAP7_75t_L g943 ( .A1(n_913), .A2(n_918), .B1(n_944), .B2(n_945), .C(n_946), .Y(n_943) );
A2O1A1Ixp33_ASAP7_75t_SL g1151 ( .A1(n_931), .A2(n_1152), .B(n_1156), .C(n_1174), .Y(n_1151) );
OAI22xp33_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_950), .B1(n_1002), .B2(n_1003), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
XOR2x2_ASAP7_75t_L g950 ( .A(n_951), .B(n_1001), .Y(n_950) );
NAND3xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_958), .C(n_975), .Y(n_953) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g1479 ( .A(n_967), .Y(n_1479) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_969), .A2(n_970), .B1(n_972), .B2(n_973), .Y(n_968) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
HB1xp67_ASAP7_75t_L g1210 ( .A(n_973), .Y(n_1210) );
OAI31xp33_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_981), .A3(n_996), .B(n_999), .Y(n_979) );
NAND3xp33_ASAP7_75t_L g981 ( .A(n_982), .B(n_987), .C(n_995), .Y(n_981) );
INVx2_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx2_ASAP7_75t_L g1120 ( .A(n_986), .Y(n_1120) );
OAI211xp5_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_989), .B(n_991), .C(n_993), .Y(n_987) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
XOR2x2_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1105), .Y(n_1003) );
AND3x1_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1041), .C(n_1072), .Y(n_1004) );
NOR2xp33_ASAP7_75t_SL g1005 ( .A(n_1006), .B(n_1027), .Y(n_1005) );
OAI33xp33_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1009), .A3(n_1012), .B1(n_1017), .B2(n_1021), .B3(n_1023), .Y(n_1006) );
BUFx8_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_1011), .A2(n_1026), .B1(n_1033), .B2(n_1035), .Y(n_1032) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1015), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_1016), .A2(n_1019), .B1(n_1030), .B2(n_1039), .Y(n_1038) );
INVx2_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1025), .Y(n_1163) );
OAI33xp33_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1029), .A3(n_1031), .B1(n_1032), .B2(n_1037), .B3(n_1038), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1472 ( .A1(n_1030), .A2(n_1039), .B1(n_1473), .B2(n_1474), .Y(n_1472) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx5_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
BUFx3_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
OAI31xp33_ASAP7_75t_L g1041 ( .A1(n_1042), .A2(n_1046), .A3(n_1056), .B(n_1069), .Y(n_1041) );
INVx4_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVx2_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx3_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1064), .B1(n_1065), .B2(n_1068), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_1064), .A2(n_1086), .B1(n_1090), .B2(n_1093), .Y(n_1085) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
BUFx3_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
OAI31xp33_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1080), .A3(n_1094), .B(n_1100), .Y(n_1072) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx2_ASAP7_75t_SL g1075 ( .A(n_1076), .Y(n_1075) );
INVx2_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVxp67_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
CKINVDCx8_ASAP7_75t_R g1083 ( .A(n_1084), .Y(n_1083) );
BUFx3_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1089), .Y(n_1087) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_1088), .B(n_1092), .Y(n_1091) );
BUFx6f_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
BUFx2_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
AND2x2_ASAP7_75t_SL g1100 ( .A(n_1101), .B(n_1103), .Y(n_1100) );
INVx1_ASAP7_75t_SL g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_1108), .A2(n_1109), .B1(n_1145), .B2(n_1146), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
HB1xp67_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1127), .Y(n_1111) );
NAND3xp33_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1117), .C(n_1124), .Y(n_1115) );
AND4x1_ASAP7_75t_L g1490 ( .A(n_1116), .B(n_1491), .C(n_1495), .D(n_1497), .Y(n_1490) );
NAND3xp33_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1133), .C(n_1138), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_1139), .A2(n_1140), .B1(n_1143), .B2(n_1144), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1486 ( .A1(n_1143), .A2(n_1144), .B1(n_1483), .B2(n_1484), .Y(n_1486) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
AOI22xp5_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1201), .B1(n_1246), .B2(n_1247), .Y(n_1146) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1147), .Y(n_1246) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
NOR3xp33_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1167), .C(n_1168), .Y(n_1156) );
NOR3xp33_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1161), .C(n_1166), .Y(n_1157) );
NOR2xp33_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1160), .Y(n_1158) );
NOR2xp33_ASAP7_75t_L g1189 ( .A(n_1159), .B(n_1185), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1164), .Y(n_1161) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
NAND3xp33_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1182), .C(n_1199), .Y(n_1176) );
INVxp67_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
AOI22xp5_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1188), .B1(n_1197), .B2(n_1198), .Y(n_1182) );
AOI22xp5_ASAP7_75t_L g1188 ( .A1(n_1184), .A2(n_1189), .B1(n_1190), .B2(n_1193), .Y(n_1188) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
HB1xp67_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx2_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
HB1xp67_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1202), .Y(n_1247) );
XOR2x2_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1245), .Y(n_1202) );
NOR2x1_ASAP7_75t_SL g1203 ( .A(n_1204), .B(n_1226), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1216), .Y(n_1207) );
OAI211xp5_ASAP7_75t_L g1208 ( .A1(n_1209), .A2(n_1210), .B(n_1211), .C(n_1212), .Y(n_1208) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVxp33_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
A2O1A1Ixp33_ASAP7_75t_SL g1226 ( .A1(n_1227), .A2(n_1230), .B(n_1241), .C(n_1243), .Y(n_1226) );
NOR3xp33_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1236), .C(n_1240), .Y(n_1230) );
INVx2_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
OAI221xp5_ASAP7_75t_L g1248 ( .A1(n_1249), .A2(n_1458), .B1(n_1461), .B2(n_1504), .C(n_1508), .Y(n_1248) );
AND4x1_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1376), .C(n_1406), .D(n_1435), .Y(n_1249) );
AOI211xp5_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1318), .B(n_1322), .C(n_1361), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
A2O1A1Ixp33_ASAP7_75t_L g1389 ( .A1(n_1252), .A2(n_1347), .B(n_1351), .C(n_1390), .Y(n_1389) );
NOR2xp33_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1306), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1300), .Y(n_1253) );
AOI22xp5_ASAP7_75t_L g1254 ( .A1(n_1255), .A2(n_1277), .B1(n_1290), .B2(n_1293), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1255), .B(n_1301), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_1255), .B(n_1279), .Y(n_1400) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
OR2x2_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1272), .Y(n_1256) );
OAI32xp33_ASAP7_75t_L g1329 ( .A1(n_1257), .A2(n_1330), .A3(n_1332), .B1(n_1337), .B2(n_1339), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1257), .B(n_1279), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1257), .B(n_1415), .Y(n_1414) );
INVx2_ASAP7_75t_L g1433 ( .A(n_1257), .Y(n_1433) );
INVx2_ASAP7_75t_SL g1257 ( .A(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1258), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1258), .B(n_1279), .Y(n_1338) );
OR2x2_ASAP7_75t_L g1346 ( .A(n_1258), .B(n_1273), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1258), .B(n_1272), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1266), .Y(n_1258) );
AND2x6_ASAP7_75t_L g1260 ( .A(n_1261), .B(n_1262), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1261), .B(n_1265), .Y(n_1264) );
AND2x4_ASAP7_75t_L g1267 ( .A(n_1261), .B(n_1268), .Y(n_1267) );
AND2x6_ASAP7_75t_L g1270 ( .A(n_1261), .B(n_1271), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1261), .B(n_1265), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1261), .B(n_1265), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1263), .B(n_1269), .Y(n_1268) );
INVx2_ASAP7_75t_L g1460 ( .A(n_1270), .Y(n_1460) );
HB1xp67_ASAP7_75t_L g1518 ( .A(n_1271), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1272), .B(n_1318), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1272), .B(n_1333), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1272), .B(n_1350), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1272), .B(n_1319), .Y(n_1397) );
OAI32xp33_ASAP7_75t_L g1411 ( .A1(n_1272), .A2(n_1273), .A3(n_1344), .B1(n_1412), .B2(n_1414), .Y(n_1411) );
HB1xp67_ASAP7_75t_SL g1436 ( .A(n_1272), .Y(n_1436) );
CKINVDCx5p33_ASAP7_75t_R g1272 ( .A(n_1273), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1273), .B(n_1292), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1273), .B(n_1356), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1273), .B(n_1319), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1273), .B(n_1280), .Y(n_1445) );
AND2x4_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1276), .Y(n_1273) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1351 ( .A(n_1278), .B(n_1315), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1283), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1279), .B(n_1340), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1279), .B(n_1315), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1279), .B(n_1345), .Y(n_1418) );
CKINVDCx14_ASAP7_75t_R g1425 ( .A(n_1279), .Y(n_1425) );
INVx3_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
CKINVDCx5p33_ASAP7_75t_R g1294 ( .A(n_1280), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1280), .B(n_1297), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1280), .B(n_1283), .Y(n_1396) );
OR2x2_ASAP7_75t_L g1401 ( .A(n_1280), .B(n_1402), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1280), .B(n_1312), .Y(n_1410) );
NOR2xp33_ASAP7_75t_L g1422 ( .A(n_1280), .B(n_1303), .Y(n_1422) );
AND2x4_ASAP7_75t_SL g1280 ( .A(n_1281), .B(n_1282), .Y(n_1280) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1283), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1283), .B(n_1315), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1283), .B(n_1305), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_1283), .B(n_1418), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1287), .Y(n_1283) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1284), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_1284), .B(n_1304), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1284), .B(n_1315), .Y(n_1314) );
NOR2xp33_ASAP7_75t_L g1342 ( .A(n_1284), .B(n_1343), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1284), .B(n_1297), .Y(n_1378) );
OR2x2_ASAP7_75t_L g1402 ( .A(n_1284), .B(n_1297), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1286), .Y(n_1284) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1287), .Y(n_1304) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1287), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1287), .B(n_1315), .Y(n_1331) );
OR2x2_ASAP7_75t_L g1367 ( .A(n_1287), .B(n_1296), .Y(n_1367) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1287), .Y(n_1399) );
NAND2x1_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1289), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1290), .B(n_1356), .Y(n_1375) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1291), .B(n_1294), .Y(n_1317) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1291), .Y(n_1420) );
OAI21xp33_ASAP7_75t_L g1307 ( .A1(n_1292), .A2(n_1308), .B(n_1311), .Y(n_1307) );
INVx2_ASAP7_75t_L g1325 ( .A(n_1292), .Y(n_1325) );
OAI21xp5_ASAP7_75t_L g1419 ( .A1(n_1293), .A2(n_1308), .B(n_1420), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1295), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1294), .B(n_1309), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1294), .B(n_1312), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1294), .B(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1294), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1294), .B(n_1432), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1451 ( .A(n_1294), .B(n_1423), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1296), .B(n_1297), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1296), .B(n_1310), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1297), .B(n_1310), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1297), .B(n_1312), .Y(n_1311) );
INVx2_ASAP7_75t_L g1315 ( .A(n_1297), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1297), .B(n_1328), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1409 ( .A(n_1297), .B(n_1410), .Y(n_1409) );
OR2x2_ASAP7_75t_L g1427 ( .A(n_1297), .B(n_1367), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1299), .Y(n_1297) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1301), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1305), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1302), .B(n_1315), .Y(n_1340) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1408 ( .A(n_1303), .B(n_1315), .Y(n_1408) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1305), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1305), .B(n_1312), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1313), .Y(n_1306) );
AOI221xp5_ASAP7_75t_L g1362 ( .A1(n_1308), .A2(n_1311), .B1(n_1326), .B2(n_1363), .C(n_1364), .Y(n_1362) );
NOR2xp33_ASAP7_75t_SL g1444 ( .A(n_1309), .B(n_1340), .Y(n_1444) );
OAI21xp5_ASAP7_75t_L g1313 ( .A1(n_1312), .A2(n_1314), .B(n_1316), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1312), .B(n_1385), .Y(n_1384) );
OAI221xp5_ASAP7_75t_L g1394 ( .A1(n_1312), .A2(n_1343), .B1(n_1367), .B2(n_1395), .C(n_1396), .Y(n_1394) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1312), .Y(n_1457) );
A2O1A1Ixp33_ASAP7_75t_L g1369 ( .A1(n_1314), .A2(n_1370), .B(n_1371), .C(n_1372), .Y(n_1369) );
OR2x2_ASAP7_75t_L g1359 ( .A(n_1315), .B(n_1360), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1315), .B(n_1399), .Y(n_1453) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
AOI21xp33_ASAP7_75t_L g1455 ( .A1(n_1317), .A2(n_1456), .B(n_1457), .Y(n_1455) );
OAI221xp5_ASAP7_75t_L g1448 ( .A1(n_1318), .A2(n_1354), .B1(n_1409), .B2(n_1449), .C(n_1452), .Y(n_1448) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1319), .B(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1319), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1321), .Y(n_1319) );
NAND4xp25_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1341), .C(n_1349), .D(n_1352), .Y(n_1322) );
O2A1O1Ixp33_ASAP7_75t_L g1323 ( .A1(n_1324), .A2(n_1326), .B(n_1327), .C(n_1329), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1325), .B(n_1356), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1325), .B(n_1392), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1325), .B(n_1413), .Y(n_1440) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1326), .Y(n_1382) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1331), .Y(n_1432) );
INVxp67_ASAP7_75t_SL g1434 ( .A(n_1332), .Y(n_1434) );
INVx3_ASAP7_75t_L g1348 ( .A(n_1333), .Y(n_1348) );
NAND3xp33_ASAP7_75t_SL g1391 ( .A(n_1333), .B(n_1351), .C(n_1392), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1333), .B(n_1356), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1336), .Y(n_1333) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1338), .Y(n_1395) );
INVx2_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
OAI211xp5_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1344), .B(n_1345), .C(n_1347), .Y(n_1341) );
INVx2_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
A2O1A1Ixp33_ASAP7_75t_L g1383 ( .A1(n_1346), .A2(n_1347), .B(n_1384), .C(n_1387), .Y(n_1383) );
A2O1A1Ixp33_ASAP7_75t_L g1407 ( .A1(n_1346), .A2(n_1408), .B(n_1409), .C(n_1411), .Y(n_1407) );
NOR2xp33_ASAP7_75t_L g1447 ( .A(n_1346), .B(n_1427), .Y(n_1447) );
AOI21xp33_ASAP7_75t_L g1421 ( .A1(n_1347), .A2(n_1422), .B(n_1423), .Y(n_1421) );
CKINVDCx14_ASAP7_75t_R g1347 ( .A(n_1348), .Y(n_1347) );
AOI31xp33_ASAP7_75t_L g1361 ( .A1(n_1348), .A2(n_1362), .A3(n_1369), .B(n_1373), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1348), .B(n_1355), .Y(n_1388) );
AOI21xp5_ASAP7_75t_L g1429 ( .A1(n_1348), .A2(n_1430), .B(n_1433), .Y(n_1429) );
A2O1A1Ixp33_ASAP7_75t_L g1452 ( .A1(n_1348), .A2(n_1453), .B(n_1454), .C(n_1455), .Y(n_1452) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1358), .Y(n_1352) );
A2O1A1Ixp33_ASAP7_75t_L g1376 ( .A1(n_1353), .A2(n_1377), .B(n_1379), .C(n_1389), .Y(n_1376) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1357), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
NAND3xp33_ASAP7_75t_L g1365 ( .A(n_1356), .B(n_1366), .C(n_1368), .Y(n_1365) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1356), .Y(n_1392) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1357), .Y(n_1423) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
OAI221xp5_ASAP7_75t_L g1379 ( .A1(n_1359), .A2(n_1380), .B1(n_1381), .B2(n_1382), .C(n_1383), .Y(n_1379) );
OR2x2_ASAP7_75t_L g1443 ( .A(n_1360), .B(n_1386), .Y(n_1443) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
NOR2xp33_ASAP7_75t_L g1374 ( .A(n_1367), .B(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1371), .Y(n_1456) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1372), .Y(n_1381) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
NOR2xp33_ASAP7_75t_L g1450 ( .A(n_1378), .B(n_1451), .Y(n_1450) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
CKINVDCx14_ASAP7_75t_R g1387 ( .A(n_1388), .Y(n_1387) );
A2O1A1O1Ixp25_ASAP7_75t_L g1435 ( .A1(n_1388), .A2(n_1436), .B(n_1437), .C(n_1438), .D(n_1448), .Y(n_1435) );
AOI221xp5_ASAP7_75t_L g1390 ( .A1(n_1391), .A2(n_1393), .B1(n_1394), .B2(n_1397), .C(n_1398), .Y(n_1390) );
AOI21xp5_ASAP7_75t_L g1406 ( .A1(n_1392), .A2(n_1407), .B(n_1416), .Y(n_1406) );
O2A1O1Ixp33_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1400), .B(n_1401), .C(n_1403), .Y(n_1398) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1400), .Y(n_1454) );
NOR2xp33_ASAP7_75t_SL g1403 ( .A(n_1404), .B(n_1405), .Y(n_1403) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1414), .Y(n_1428) );
AOI331xp33_ASAP7_75t_L g1416 ( .A1(n_1417), .A2(n_1419), .A3(n_1421), .B1(n_1424), .B2(n_1428), .B3(n_1429), .C1(n_1434), .Y(n_1416) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1424), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1426), .Y(n_1424) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
NOR2xp33_ASAP7_75t_SL g1441 ( .A(n_1433), .B(n_1442), .Y(n_1441) );
OAI221xp5_ASAP7_75t_L g1438 ( .A1(n_1439), .A2(n_1441), .B1(n_1444), .B2(n_1445), .C(n_1446), .Y(n_1438) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
INVxp67_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
INVxp67_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
CKINVDCx20_ASAP7_75t_R g1458 ( .A(n_1459), .Y(n_1458) );
CKINVDCx20_ASAP7_75t_R g1459 ( .A(n_1460), .Y(n_1459) );
HB1xp67_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVxp33_ASAP7_75t_L g1515 ( .A(n_1463), .Y(n_1515) );
NOR2x1p5_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1487), .Y(n_1463) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1490), .Y(n_1487) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
BUFx3_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
BUFx3_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
BUFx3_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
INVxp33_ASAP7_75t_SL g1512 ( .A(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
HB1xp67_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
OAI21xp5_ASAP7_75t_L g1517 ( .A1(n_1518), .A2(n_1519), .B(n_1520), .Y(n_1517) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
endmodule