module fake_netlist_6_4257_n_1220 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1220);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1220;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_881;
wire n_1199;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_680;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_886;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_1203;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1217;
wire n_751;
wire n_449;
wire n_749;
wire n_1208;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_1209;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_1214;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1204;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_1101;
wire n_1099;
wire n_1026;
wire n_443;
wire n_485;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_1192;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1212;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_963;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_1206;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_1196;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_1205;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_720;
wire n_525;
wire n_842;
wire n_1173;
wire n_1163;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_1219;
wire n_1216;
wire n_843;
wire n_656;
wire n_772;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_953;
wire n_448;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_1213;
wire n_638;
wire n_234;
wire n_1181;
wire n_910;
wire n_1211;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_1215;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_1084;
wire n_460;
wire n_929;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_1195;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_813;
wire n_395;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_1201;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_608;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_1218;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_1198;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_273;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_882;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1207;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_1210;
wire n_679;
wire n_1069;
wire n_1185;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1200;
wire n_1059;
wire n_1197;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_1098;
wire n_391;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_385;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_736;
wire n_613;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_94),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_8),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

BUFx2_ASAP7_75t_R g187 ( 
.A(n_105),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_83),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_34),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_35),
.Y(n_192)
);

BUFx8_ASAP7_75t_SL g193 ( 
.A(n_116),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_15),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_73),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_95),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_107),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_109),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_40),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_144),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_81),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_34),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_164),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_111),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_35),
.Y(n_208)
);

BUFx2_ASAP7_75t_SL g209 ( 
.A(n_48),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_48),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_10),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_152),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_161),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_49),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_128),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_121),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_166),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_14),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_69),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_173),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_51),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_168),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_52),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_39),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_79),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_113),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_80),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_13),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_123),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_101),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_68),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_91),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_7),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_47),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_71),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_63),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_134),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_3),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_60),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_61),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_167),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_70),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_104),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_27),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_93),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_131),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_142),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_49),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_37),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_159),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_37),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_75),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_158),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_24),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_18),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_124),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_86),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_33),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_92),
.Y(n_268)
);

CKINVDCx6p67_ASAP7_75t_R g269 ( 
.A(n_57),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_17),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_119),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_148),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_18),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_4),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_130),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_55),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_66),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_0),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_53),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_38),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_88),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_14),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_120),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_133),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_102),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_22),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_67),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_146),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_58),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_2),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_117),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_57),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_196),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_213),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_232),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_193),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_181),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_197),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_0),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_199),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_196),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_231),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_200),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_202),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_209),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_203),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_189),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_196),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_206),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_192),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_284),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_196),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_207),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_238),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_196),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_209),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_212),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_201),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_201),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_216),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_218),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_221),
.B(n_1),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_182),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_220),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_208),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_221),
.B(n_258),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_224),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_258),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_227),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_285),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_263),
.B(n_1),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_251),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_263),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_186),
.B(n_2),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_267),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_237),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_267),
.Y(n_342)
);

BUFx2_ASAP7_75t_SL g343 ( 
.A(n_182),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_282),
.B(n_3),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_282),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_185),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_245),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_245),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_239),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_242),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_186),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_188),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_244),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_188),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_247),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_190),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_210),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_190),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_211),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_250),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_214),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_253),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_254),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_256),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_191),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_228),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_191),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_230),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_185),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_194),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_259),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_194),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_195),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_229),
.B(n_4),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_195),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_235),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_182),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_261),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_294),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_262),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_303),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_294),
.B(n_271),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_302),
.B(n_217),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_302),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

OA21x2_ASAP7_75t_L g387 ( 
.A1(n_303),
.A2(n_204),
.B(n_198),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_346),
.B(n_217),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_320),
.Y(n_393)
);

AND2x2_ASAP7_75t_SL g394 ( 
.A(n_300),
.B(n_229),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_335),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_215),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_243),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_351),
.B(n_275),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_352),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_315),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_343),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_343),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_361),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g412 ( 
.A1(n_354),
.A2(n_204),
.B(n_198),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_316),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_243),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_283),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_356),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_358),
.B(n_222),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_358),
.B(n_290),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_365),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_365),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_324),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_367),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_370),
.B(n_183),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_372),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_373),
.B(n_265),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_219),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_375),
.B(n_347),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g433 ( 
.A(n_339),
.B(n_265),
.Y(n_433)
);

NOR2x1_ASAP7_75t_L g434 ( 
.A(n_318),
.B(n_287),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_333),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_295),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_333),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_338),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_340),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_347),
.B(n_222),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_348),
.B(n_223),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_368),
.B(n_281),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_340),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_329),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_342),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_304),
.A2(n_264),
.B1(n_205),
.B2(n_225),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_384),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_444),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_408),
.B(n_328),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_389),
.B(n_296),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_408),
.B(n_328),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_327),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_389),
.Y(n_458)
);

OR2x6_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_327),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_409),
.B(n_298),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_394),
.A2(n_307),
.B1(n_319),
.B2(n_344),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_411),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_433),
.B(n_309),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_409),
.B(n_377),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

NOR2x1p5_ASAP7_75t_L g466 ( 
.A(n_426),
.B(n_269),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_410),
.B(n_377),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_426),
.A2(n_269),
.B1(n_307),
.B2(n_331),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_321),
.Y(n_469)
);

OAI22xp33_ASAP7_75t_L g470 ( 
.A1(n_431),
.A2(n_331),
.B1(n_286),
.B2(n_184),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_380),
.B(n_299),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_287),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_427),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_444),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_394),
.A2(n_305),
.B1(n_336),
.B2(n_344),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_384),
.B(n_223),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_394),
.A2(n_336),
.B1(n_330),
.B2(n_357),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_381),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_394),
.A2(n_270),
.B1(n_276),
.B2(n_240),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_381),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_400),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_433),
.A2(n_359),
.B1(n_366),
.B2(n_226),
.Y(n_487)
);

AO21x2_ASAP7_75t_L g488 ( 
.A1(n_431),
.A2(n_233),
.B(n_226),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_384),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_382),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_433),
.B(n_233),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_428),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_399),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_443),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_389),
.B(n_348),
.Y(n_495)
);

BUFx10_ASAP7_75t_L g496 ( 
.A(n_443),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_398),
.A2(n_293),
.B1(n_279),
.B2(n_241),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_410),
.B(n_301),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_428),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_433),
.B(n_234),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_429),
.Y(n_502)
);

AND3x2_ASAP7_75t_L g503 ( 
.A(n_398),
.B(n_410),
.C(n_397),
.Y(n_503)
);

OR2x6_ASAP7_75t_L g504 ( 
.A(n_403),
.B(n_234),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_429),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_382),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_382),
.Y(n_507)
);

INVx6_ASAP7_75t_L g508 ( 
.A(n_384),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_396),
.Y(n_509)
);

OAI21xp33_ASAP7_75t_SL g510 ( 
.A1(n_441),
.A2(n_246),
.B(n_236),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_403),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_396),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_433),
.B(n_236),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_429),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_379),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_400),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_487),
.A2(n_407),
.B1(n_341),
.B2(n_355),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_481),
.A2(n_407),
.B1(n_350),
.B2(n_362),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_449),
.Y(n_519)
);

NAND2x1_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_425),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_465),
.B(n_397),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_471),
.B(n_380),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_462),
.B(n_403),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_458),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_449),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_453),
.B(n_376),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_SL g527 ( 
.A(n_479),
.B(n_248),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_462),
.B(n_433),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_465),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_463),
.B(n_306),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_463),
.B(n_308),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_469),
.B(n_449),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_452),
.Y(n_533)
);

INVx8_ASAP7_75t_L g534 ( 
.A(n_504),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_473),
.Y(n_535)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_460),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_453),
.B(n_413),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_474),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_475),
.B(n_310),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_475),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_458),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_483),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_483),
.B(n_413),
.Y(n_544)
);

NOR2xp67_ASAP7_75t_L g545 ( 
.A(n_454),
.B(n_297),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_494),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_476),
.B(n_314),
.Y(n_547)
);

INVxp33_ASAP7_75t_L g548 ( 
.A(n_495),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_476),
.B(n_322),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_489),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_489),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_469),
.B(n_325),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_489),
.B(n_326),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_494),
.B(n_332),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_495),
.B(n_432),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_493),
.B(n_436),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_477),
.B(n_334),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_494),
.B(n_360),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_494),
.B(n_378),
.Y(n_560)
);

O2A1O1Ixp33_ASAP7_75t_L g561 ( 
.A1(n_510),
.A2(n_419),
.B(n_415),
.C(n_404),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_493),
.B(n_349),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_492),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_456),
.A2(n_313),
.B1(n_364),
.B2(n_363),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_515),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_508),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_515),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_480),
.B(n_432),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_496),
.B(n_353),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_511),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_496),
.B(n_371),
.Y(n_571)
);

NOR2xp67_ASAP7_75t_L g572 ( 
.A(n_464),
.B(n_445),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_499),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_496),
.B(n_425),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_499),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_496),
.B(n_491),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_502),
.B(n_383),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_508),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_502),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_505),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_505),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_511),
.B(n_436),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_461),
.B(n_415),
.C(n_404),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_514),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_514),
.B(n_383),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_498),
.B(n_445),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_504),
.B(n_441),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_508),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_467),
.B(n_419),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_484),
.B(n_448),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_456),
.B(n_448),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_508),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_497),
.Y(n_593)
);

INVx8_ASAP7_75t_L g594 ( 
.A(n_504),
.Y(n_594)
);

NOR3xp33_ASAP7_75t_L g595 ( 
.A(n_470),
.B(n_345),
.C(n_323),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_504),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_480),
.B(n_425),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_480),
.B(n_425),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_456),
.A2(n_459),
.B1(n_504),
.B2(n_480),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_491),
.B(n_425),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_501),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_450),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_488),
.A2(n_412),
.B1(n_387),
.B2(n_430),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_501),
.B(n_285),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_456),
.A2(n_401),
.B1(n_414),
.B2(n_384),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_497),
.B(n_432),
.Y(n_606)
);

AO21x1_ASAP7_75t_L g607 ( 
.A1(n_527),
.A2(n_513),
.B(n_472),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_535),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_527),
.A2(n_522),
.B(n_591),
.C(n_561),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_525),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_599),
.B(n_513),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_536),
.B(n_503),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_605),
.B(n_472),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_577),
.B(n_459),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_532),
.A2(n_585),
.B(n_597),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_526),
.B(n_459),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_537),
.B(n_484),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_535),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_538),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_536),
.B(n_503),
.Y(n_620)
);

BUFx5_ASAP7_75t_L g621 ( 
.A(n_588),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_525),
.Y(n_622)
);

AOI33xp33_ASAP7_75t_L g623 ( 
.A1(n_524),
.A2(n_470),
.A3(n_468),
.B1(n_423),
.B2(n_417),
.B3(n_442),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_538),
.Y(n_624)
);

OAI21xp33_ASAP7_75t_L g625 ( 
.A1(n_548),
.A2(n_542),
.B(n_593),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_539),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_529),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_539),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_523),
.B(n_459),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_583),
.B(n_459),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_598),
.A2(n_478),
.B(n_451),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_543),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_525),
.B(n_451),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_596),
.A2(n_601),
.B1(n_551),
.B2(n_519),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_555),
.B(n_488),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_548),
.B(n_468),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_555),
.B(n_437),
.Y(n_637)
);

AO21x1_ASAP7_75t_L g638 ( 
.A1(n_576),
.A2(n_249),
.B(n_248),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_544),
.B(n_466),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_555),
.B(n_466),
.Y(n_640)
);

OAI21xp33_ASAP7_75t_L g641 ( 
.A1(n_590),
.A2(n_442),
.B(n_441),
.Y(n_641)
);

BUFx12f_ASAP7_75t_L g642 ( 
.A(n_556),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_573),
.B(n_437),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_521),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_581),
.B(n_437),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_529),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_541),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_525),
.Y(n_648)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_606),
.A2(n_442),
.B(n_418),
.C(n_268),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_568),
.B(n_437),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_576),
.A2(n_418),
.B(n_384),
.C(n_414),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_568),
.B(n_417),
.Y(n_652)
);

AO21x1_ASAP7_75t_L g653 ( 
.A1(n_574),
.A2(n_266),
.B(n_249),
.Y(n_653)
);

OA21x2_ASAP7_75t_L g654 ( 
.A1(n_603),
.A2(n_455),
.B(n_450),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_541),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_519),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_562),
.B(n_187),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_519),
.B(n_478),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_570),
.Y(n_659)
);

AOI33xp33_ASAP7_75t_L g660 ( 
.A1(n_570),
.A2(n_423),
.A3(n_435),
.B1(n_438),
.B2(n_440),
.B3(n_418),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_L g661 ( 
.A(n_518),
.B(n_517),
.C(n_559),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_528),
.A2(n_486),
.B(n_457),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_558),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_255),
.C(n_252),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_533),
.Y(n_665)
);

NOR3xp33_ASAP7_75t_L g666 ( 
.A(n_560),
.B(n_272),
.C(n_268),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_520),
.A2(n_486),
.B(n_457),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_569),
.B(n_401),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_558),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_592),
.A2(n_486),
.B(n_457),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_589),
.B(n_540),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_600),
.A2(n_516),
.B(n_486),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_563),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_546),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_L g675 ( 
.A(n_586),
.B(n_277),
.C(n_272),
.Y(n_675)
);

O2A1O1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_574),
.A2(n_552),
.B(n_530),
.C(n_531),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_568),
.B(n_547),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_531),
.A2(n_552),
.B(n_566),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_563),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_566),
.A2(n_516),
.B(n_405),
.Y(n_680)
);

CKINVDCx8_ASAP7_75t_R g681 ( 
.A(n_546),
.Y(n_681)
);

BUFx12f_ASAP7_75t_L g682 ( 
.A(n_587),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_549),
.A2(n_401),
.B1(n_414),
.B2(n_430),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_566),
.A2(n_516),
.B(n_405),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_575),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_575),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_595),
.B(n_414),
.Y(n_687)
);

AO22x1_ASAP7_75t_L g688 ( 
.A1(n_550),
.A2(n_291),
.B1(n_257),
.B2(n_289),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_564),
.B(n_414),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_600),
.A2(n_516),
.B(n_455),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_557),
.B(n_437),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_579),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_551),
.A2(n_405),
.B(n_402),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_551),
.A2(n_405),
.B(n_402),
.Y(n_694)
);

NOR2x1_ASAP7_75t_L g695 ( 
.A(n_554),
.B(n_379),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_579),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_610),
.Y(n_697)
);

O2A1O1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_609),
.A2(n_554),
.B(n_571),
.C(n_553),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_624),
.Y(n_699)
);

AOI21x1_ASAP7_75t_L g700 ( 
.A1(n_678),
.A2(n_567),
.B(n_565),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_671),
.B(n_550),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_624),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_SL g703 ( 
.A(n_674),
.B(n_533),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_671),
.B(n_571),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_661),
.A2(n_572),
.B(n_534),
.C(n_594),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_644),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_614),
.B(n_580),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_664),
.B(n_545),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_610),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_632),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_610),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_642),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_616),
.B(n_584),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_L g714 ( 
.A(n_612),
.B(n_604),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_629),
.B(n_534),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_617),
.B(n_587),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_626),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_636),
.B(n_587),
.Y(n_718)
);

OAI22x1_ASAP7_75t_L g719 ( 
.A1(n_636),
.A2(n_620),
.B1(n_612),
.B2(n_657),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_630),
.B(n_578),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_615),
.A2(n_578),
.B(n_602),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_641),
.B(n_578),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_677),
.B(n_578),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_610),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_668),
.B(n_652),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_675),
.A2(n_412),
.B1(n_277),
.B2(n_288),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_632),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_SL g728 ( 
.A1(n_665),
.A2(n_280),
.B1(n_260),
.B2(n_274),
.Y(n_728)
);

BUFx12f_ASAP7_75t_L g729 ( 
.A(n_646),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_687),
.A2(n_602),
.B1(n_430),
.B2(n_288),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_627),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_676),
.A2(n_430),
.B(n_406),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_658),
.A2(n_406),
.B(n_402),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_640),
.B(n_435),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_658),
.A2(n_406),
.B(n_402),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_626),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_622),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_SL g738 ( 
.A(n_639),
.B(n_273),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_647),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_675),
.A2(n_435),
.B(n_438),
.C(n_440),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_625),
.B(n_438),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_666),
.A2(n_440),
.B(n_406),
.C(n_416),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_633),
.A2(n_420),
.B(n_416),
.Y(n_743)
);

INVxp33_ASAP7_75t_SL g744 ( 
.A(n_620),
.Y(n_744)
);

OR2x6_ASAP7_75t_L g745 ( 
.A(n_682),
.B(n_285),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_659),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_635),
.A2(n_412),
.B1(n_387),
.B2(n_420),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_656),
.B(n_285),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_647),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_690),
.A2(n_387),
.B(n_412),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_666),
.A2(n_412),
.B1(n_182),
.B2(n_387),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_663),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_691),
.A2(n_387),
.B1(n_422),
.B2(n_416),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_627),
.B(n_652),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_623),
.A2(n_651),
.B(n_689),
.C(n_649),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_623),
.B(n_439),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_688),
.B(n_446),
.C(n_439),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_640),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_663),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_656),
.A2(n_611),
.B1(n_683),
.B2(n_634),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_649),
.A2(n_379),
.B(n_386),
.C(n_439),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_699),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_727),
.B(n_622),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_721),
.A2(n_662),
.B(n_631),
.Y(n_764)
);

O2A1O1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_704),
.A2(n_637),
.B(n_650),
.C(n_607),
.Y(n_765)
);

BUFx12f_ASAP7_75t_L g766 ( 
.A(n_729),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_712),
.Y(n_767)
);

OAI21x1_ASAP7_75t_SL g768 ( 
.A1(n_698),
.A2(n_653),
.B(n_638),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_717),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_704),
.B(n_679),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_736),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_701),
.B(n_679),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_706),
.B(n_619),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_707),
.B(n_685),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_754),
.Y(n_775)
);

INVx6_ASAP7_75t_L g776 ( 
.A(n_734),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_713),
.B(n_685),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_749),
.Y(n_778)
);

AO22x2_ASAP7_75t_L g779 ( 
.A1(n_760),
.A2(n_696),
.B1(n_618),
.B2(n_628),
.Y(n_779)
);

AO31x2_ASAP7_75t_L g780 ( 
.A1(n_753),
.A2(n_686),
.A3(n_673),
.B(n_655),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_700),
.A2(n_694),
.B(n_693),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_SL g782 ( 
.A1(n_755),
.A2(n_643),
.B(n_645),
.C(n_608),
.Y(n_782)
);

AOI221xp5_ASAP7_75t_L g783 ( 
.A1(n_719),
.A2(n_669),
.B1(n_446),
.B2(n_692),
.C(n_686),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_744),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_718),
.A2(n_695),
.B(n_660),
.C(n_684),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_718),
.A2(n_660),
.B(n_680),
.C(n_670),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_737),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_716),
.B(n_725),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_758),
.B(n_648),
.Y(n_789)
);

AO21x1_ASAP7_75t_L g790 ( 
.A1(n_720),
.A2(n_672),
.B(n_667),
.Y(n_790)
);

OAI21x1_ASAP7_75t_L g791 ( 
.A1(n_750),
.A2(n_654),
.B(n_648),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_702),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_731),
.B(n_681),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_710),
.Y(n_794)
);

O2A1O1Ixp5_ASAP7_75t_L g795 ( 
.A1(n_720),
.A2(n_390),
.B(n_388),
.C(n_385),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_732),
.A2(n_654),
.B(n_390),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_733),
.A2(n_490),
.B(n_450),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_754),
.B(n_703),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_739),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_726),
.A2(n_613),
.B1(n_446),
.B2(n_420),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_752),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_716),
.A2(n_613),
.B1(n_621),
.B2(n_446),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_723),
.B(n_613),
.Y(n_803)
);

OAI21x1_ASAP7_75t_L g804 ( 
.A1(n_735),
.A2(n_490),
.B(n_455),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_759),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_743),
.A2(n_500),
.B(n_482),
.Y(n_806)
);

OA21x2_ASAP7_75t_L g807 ( 
.A1(n_761),
.A2(n_385),
.B(n_388),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_756),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_758),
.A2(n_613),
.B1(n_444),
.B2(n_447),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_746),
.Y(n_810)
);

AOI31xp67_ASAP7_75t_L g811 ( 
.A1(n_748),
.A2(n_421),
.A3(n_422),
.B(n_424),
.Y(n_811)
);

AO31x2_ASAP7_75t_L g812 ( 
.A1(n_705),
.A2(n_421),
.A3(n_422),
.B(n_424),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_714),
.B(n_613),
.Y(n_813)
);

OR2x6_ASAP7_75t_L g814 ( 
.A(n_709),
.B(n_621),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_715),
.B(n_621),
.Y(n_815)
);

OAI21x1_ASAP7_75t_L g816 ( 
.A1(n_747),
.A2(n_490),
.B(n_512),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_801),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_798),
.A2(n_726),
.B1(n_708),
.B2(n_741),
.Y(n_818)
);

BUFx8_ASAP7_75t_SL g819 ( 
.A(n_767),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_792),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_799),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_788),
.A2(n_728),
.B1(n_738),
.B2(n_813),
.Y(n_822)
);

CKINVDCx6p67_ASAP7_75t_R g823 ( 
.A(n_766),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_788),
.A2(n_741),
.B1(n_722),
.B2(n_751),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_775),
.A2(n_751),
.B1(n_734),
.B2(n_730),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_784),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_805),
.Y(n_827)
);

INVx6_ASAP7_75t_L g828 ( 
.A(n_776),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_762),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_802),
.A2(n_745),
.B1(n_737),
.B2(n_724),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_814),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_769),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_770),
.B(n_740),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_771),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_789),
.B(n_697),
.Y(n_835)
);

INVx6_ASAP7_75t_L g836 ( 
.A(n_776),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_778),
.Y(n_837)
);

BUFx4f_ASAP7_75t_SL g838 ( 
.A(n_794),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_813),
.A2(n_745),
.B1(n_709),
.B2(n_711),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_810),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_803),
.A2(n_757),
.B1(n_745),
.B2(n_748),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_803),
.A2(n_808),
.B1(n_783),
.B2(n_793),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_773),
.A2(n_724),
.B1(n_697),
.B2(n_711),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_772),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_770),
.A2(n_709),
.B1(n_447),
.B2(n_444),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_763),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_815),
.A2(n_709),
.B(n_757),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_789),
.A2(n_621),
.B1(n_386),
.B2(n_422),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_772),
.B(n_742),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_777),
.B(n_621),
.Y(n_850)
);

OAI22xp33_ASAP7_75t_L g851 ( 
.A1(n_763),
.A2(n_447),
.B1(n_444),
.B2(n_386),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_783),
.A2(n_621),
.B1(n_386),
.B2(n_421),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_763),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_777),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_774),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_787),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_774),
.B(n_444),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_791),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_765),
.B(n_444),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_779),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_768),
.A2(n_444),
.B1(n_447),
.B2(n_385),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_787),
.Y(n_862)
);

OAI22xp33_ASAP7_75t_L g863 ( 
.A1(n_815),
.A2(n_447),
.B1(n_392),
.B2(n_393),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_779),
.Y(n_864)
);

CKINVDCx6p67_ASAP7_75t_R g865 ( 
.A(n_814),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_800),
.A2(n_447),
.B1(n_388),
.B2(n_392),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_800),
.A2(n_447),
.B1(n_392),
.B2(n_393),
.Y(n_867)
);

INVx6_ASAP7_75t_L g868 ( 
.A(n_814),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_807),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_790),
.A2(n_447),
.B1(n_393),
.B2(n_395),
.Y(n_870)
);

BUFx4_ASAP7_75t_SL g871 ( 
.A(n_782),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_807),
.Y(n_872)
);

BUFx10_ASAP7_75t_L g873 ( 
.A(n_785),
.Y(n_873)
);

INVx6_ASAP7_75t_L g874 ( 
.A(n_786),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_796),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_780),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_876),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_860),
.B(n_780),
.Y(n_878)
);

INVx6_ASAP7_75t_L g879 ( 
.A(n_831),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_864),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_844),
.B(n_809),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_875),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_875),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_869),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_832),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_858),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_869),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_869),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_872),
.Y(n_889)
);

OAI21xp33_ASAP7_75t_SL g890 ( 
.A1(n_842),
.A2(n_781),
.B(n_764),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_858),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_845),
.A2(n_816),
.B(n_795),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_869),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_832),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_868),
.Y(n_895)
);

AO21x2_ASAP7_75t_L g896 ( 
.A1(n_859),
.A2(n_804),
.B(n_797),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_834),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_868),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_834),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_831),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_829),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_854),
.B(n_812),
.Y(n_902)
);

OA21x2_ASAP7_75t_L g903 ( 
.A1(n_847),
.A2(n_806),
.B(n_812),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_837),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_862),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_874),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_831),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_874),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_874),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_874),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_820),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_820),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_868),
.Y(n_913)
);

HB1xp67_ASAP7_75t_SL g914 ( 
.A(n_835),
.Y(n_914)
);

AO32x1_ASAP7_75t_L g915 ( 
.A1(n_877),
.A2(n_818),
.A3(n_843),
.B1(n_824),
.B2(n_853),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_898),
.B(n_853),
.Y(n_916)
);

OAI211xp5_ASAP7_75t_L g917 ( 
.A1(n_909),
.A2(n_822),
.B(n_839),
.C(n_841),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_909),
.A2(n_846),
.B1(n_825),
.B2(n_840),
.Y(n_918)
);

NOR2x1_ASAP7_75t_SL g919 ( 
.A(n_895),
.B(n_855),
.Y(n_919)
);

NOR2x1_ASAP7_75t_SL g920 ( 
.A(n_895),
.B(n_821),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_904),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_898),
.B(n_827),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_906),
.A2(n_873),
.B1(n_846),
.B2(n_868),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_904),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_898),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_914),
.A2(n_833),
.B1(n_865),
.B2(n_849),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_898),
.B(n_827),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_906),
.Y(n_928)
);

OA21x2_ASAP7_75t_L g929 ( 
.A1(n_892),
.A2(n_870),
.B(n_857),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_895),
.Y(n_930)
);

NAND4xp25_ASAP7_75t_L g931 ( 
.A(n_905),
.B(n_817),
.C(n_861),
.D(n_830),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_913),
.B(n_835),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_905),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_904),
.B(n_850),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_906),
.A2(n_823),
.B1(n_873),
.B2(n_838),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_894),
.B(n_873),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_880),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_913),
.B(n_835),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_SL g939 ( 
.A1(n_895),
.A2(n_881),
.B(n_908),
.Y(n_939)
);

AO21x2_ASAP7_75t_L g940 ( 
.A1(n_892),
.A2(n_902),
.B(n_888),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_901),
.B(n_817),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_908),
.B(n_826),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_880),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_913),
.B(n_856),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_894),
.B(n_865),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_914),
.A2(n_867),
.B1(n_866),
.B2(n_852),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_880),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_901),
.B(n_885),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_879),
.B(n_828),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_908),
.A2(n_910),
.B1(n_823),
.B2(n_895),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_890),
.A2(n_848),
.B(n_851),
.Y(n_951)
);

AOI221xp5_ASAP7_75t_L g952 ( 
.A1(n_908),
.A2(n_863),
.B1(n_395),
.B2(n_826),
.C(n_871),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_889),
.B(n_395),
.Y(n_953)
);

OAI221xp5_ASAP7_75t_L g954 ( 
.A1(n_890),
.A2(n_828),
.B1(n_836),
.B2(n_7),
.C(n_8),
.Y(n_954)
);

OA21x2_ASAP7_75t_L g955 ( 
.A1(n_877),
.A2(n_902),
.B(n_881),
.Y(n_955)
);

NOR2x1_ASAP7_75t_L g956 ( 
.A(n_900),
.B(n_819),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_921),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_924),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_955),
.B(n_877),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_955),
.B(n_877),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_937),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_SL g962 ( 
.A1(n_954),
.A2(n_910),
.B1(n_895),
.B2(n_879),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_930),
.B(n_884),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_943),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_947),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_948),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_941),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_940),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_940),
.B(n_878),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_936),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_939),
.B(n_884),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_930),
.B(n_884),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_936),
.B(n_889),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_920),
.B(n_888),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_919),
.B(n_888),
.Y(n_975)
);

INVx5_ASAP7_75t_L g976 ( 
.A(n_949),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_918),
.A2(n_910),
.B1(n_879),
.B2(n_900),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_922),
.B(n_893),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_934),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_927),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_925),
.B(n_893),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_945),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_945),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_971),
.B(n_893),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_958),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_980),
.B(n_916),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_SL g987 ( 
.A1(n_982),
.A2(n_933),
.B1(n_926),
.B2(n_942),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_958),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_971),
.B(n_887),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_959),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_971),
.B(n_887),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_958),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_958),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_961),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_980),
.B(n_925),
.Y(n_995)
);

AOI221xp5_ASAP7_75t_L g996 ( 
.A1(n_962),
.A2(n_954),
.B1(n_917),
.B2(n_926),
.C(n_931),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_959),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_961),
.Y(n_998)
);

OAI33xp33_ASAP7_75t_L g999 ( 
.A1(n_973),
.A2(n_983),
.A3(n_982),
.B1(n_969),
.B2(n_957),
.B3(n_964),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_974),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_979),
.B(n_970),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_980),
.B(n_959),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_980),
.B(n_887),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_SL g1004 ( 
.A1(n_976),
.A2(n_928),
.B1(n_951),
.B2(n_910),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_986),
.B(n_983),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_1000),
.B(n_976),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_995),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_985),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_985),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_988),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_986),
.B(n_970),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_988),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_990),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_992),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_987),
.B(n_979),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_992),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1008),
.Y(n_1017)
);

NAND2x2_ASAP7_75t_L g1018 ( 
.A(n_1015),
.B(n_1000),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1008),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1006),
.B(n_1000),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_1006),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_1013),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_1011),
.B(n_1005),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1009),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1017),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1021),
.B(n_1007),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1019),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1020),
.B(n_989),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_1023),
.B(n_1013),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_1026),
.B(n_819),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_SL g1031 ( 
.A1(n_1028),
.A2(n_1018),
.B1(n_987),
.B2(n_1020),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1028),
.Y(n_1032)
);

AOI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_1025),
.A2(n_1021),
.B1(n_996),
.B2(n_999),
.C(n_1024),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1029),
.B(n_1023),
.Y(n_1034)
);

AOI221xp5_ASAP7_75t_SL g1035 ( 
.A1(n_1027),
.A2(n_996),
.B1(n_1018),
.B2(n_991),
.C(n_989),
.Y(n_1035)
);

OAI32xp33_ASAP7_75t_L g1036 ( 
.A1(n_1029),
.A2(n_1022),
.A3(n_969),
.B1(n_968),
.B2(n_1001),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1025),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1025),
.B(n_984),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1025),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1028),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1025),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_1030),
.B(n_956),
.C(n_935),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_1032),
.B(n_1022),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_1031),
.B(n_1004),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1030),
.B(n_1002),
.Y(n_1045)
);

AOI221xp5_ASAP7_75t_L g1046 ( 
.A1(n_1035),
.A2(n_999),
.B1(n_1022),
.B2(n_962),
.C(n_1004),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_1034),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1037),
.Y(n_1048)
);

AOI211xp5_ASAP7_75t_L g1049 ( 
.A1(n_1033),
.A2(n_952),
.B(n_931),
.C(n_946),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1032),
.B(n_989),
.Y(n_1050)
);

OAI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_1040),
.A2(n_976),
.B1(n_977),
.B2(n_969),
.Y(n_1051)
);

OA211x2_ASAP7_75t_L g1052 ( 
.A1(n_1038),
.A2(n_923),
.B(n_973),
.C(n_951),
.Y(n_1052)
);

AOI22x1_ASAP7_75t_SL g1053 ( 
.A1(n_1041),
.A2(n_1016),
.B1(n_1009),
.B2(n_1012),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1040),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1034),
.A2(n_1039),
.B(n_1036),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_1032),
.B(n_1016),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1031),
.A2(n_976),
.B1(n_977),
.B2(n_991),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_1030),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1044),
.A2(n_915),
.B(n_1010),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1047),
.B(n_991),
.Y(n_1060)
);

NOR4xp25_ASAP7_75t_L g1061 ( 
.A(n_1058),
.B(n_1014),
.C(n_953),
.D(n_1001),
.Y(n_1061)
);

AOI222xp33_ASAP7_75t_L g1062 ( 
.A1(n_1055),
.A2(n_1046),
.B1(n_1057),
.B2(n_1048),
.C1(n_1045),
.C2(n_1054),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1043),
.Y(n_1063)
);

OAI31xp33_ASAP7_75t_L g1064 ( 
.A1(n_1051),
.A2(n_984),
.A3(n_968),
.B(n_946),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1049),
.A2(n_950),
.B1(n_968),
.B2(n_928),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_1053),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_1042),
.B(n_984),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1049),
.B(n_990),
.Y(n_1068)
);

NAND3x1_ASAP7_75t_L g1069 ( 
.A(n_1050),
.B(n_1002),
.C(n_995),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1056),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1056),
.Y(n_1071)
);

XNOR2xp5_ASAP7_75t_L g1072 ( 
.A(n_1052),
.B(n_932),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1047),
.B(n_990),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_SL g1074 ( 
.A1(n_1044),
.A2(n_997),
.B(n_965),
.C(n_993),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1054),
.Y(n_1075)
);

OAI21xp33_ASAP7_75t_SL g1076 ( 
.A1(n_1044),
.A2(n_1002),
.B(n_997),
.Y(n_1076)
);

NAND5xp2_ASAP7_75t_L g1077 ( 
.A(n_1058),
.B(n_1003),
.C(n_967),
.D(n_912),
.E(n_972),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1070),
.Y(n_1078)
);

NOR3xp33_ASAP7_75t_L g1079 ( 
.A(n_1063),
.B(n_1066),
.C(n_1075),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_1061),
.B(n_976),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1068),
.B(n_997),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_SL g1082 ( 
.A(n_1064),
.B(n_976),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_1062),
.B(n_968),
.C(n_976),
.Y(n_1083)
);

AOI211xp5_ASAP7_75t_L g1084 ( 
.A1(n_1076),
.A2(n_975),
.B(n_974),
.C(n_9),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1071),
.Y(n_1085)
);

NOR3x1_ASAP7_75t_L g1086 ( 
.A(n_1060),
.B(n_965),
.C(n_966),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_1072),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1073),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1067),
.B(n_976),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1065),
.B(n_836),
.Y(n_1090)
);

NAND5xp2_ASAP7_75t_L g1091 ( 
.A(n_1065),
.B(n_1003),
.C(n_6),
.D(n_9),
.E(n_10),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1067),
.B(n_976),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_L g1093 ( 
.A(n_1059),
.B(n_907),
.C(n_900),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1074),
.B(n_979),
.Y(n_1094)
);

AOI221xp5_ASAP7_75t_L g1095 ( 
.A1(n_1083),
.A2(n_1077),
.B1(n_1069),
.B2(n_998),
.C(n_994),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1079),
.B(n_1003),
.Y(n_1096)
);

OAI211xp5_ASAP7_75t_SL g1097 ( 
.A1(n_1087),
.A2(n_5),
.B(n_6),
.C(n_11),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1078),
.Y(n_1098)
);

AOI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_1091),
.A2(n_998),
.B1(n_994),
.B2(n_993),
.C(n_967),
.Y(n_1099)
);

AOI221xp5_ASAP7_75t_SL g1100 ( 
.A1(n_1091),
.A2(n_966),
.B1(n_979),
.B2(n_957),
.C(n_964),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1082),
.A2(n_975),
.B1(n_974),
.B2(n_963),
.Y(n_1101)
);

NOR3x1_ASAP7_75t_L g1102 ( 
.A(n_1085),
.B(n_965),
.C(n_966),
.Y(n_1102)
);

AOI221x1_ASAP7_75t_L g1103 ( 
.A1(n_1090),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_1103)
);

AND5x1_ASAP7_75t_L g1104 ( 
.A(n_1084),
.B(n_12),
.C(n_15),
.D(n_16),
.E(n_17),
.Y(n_1104)
);

AOI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1093),
.A2(n_974),
.B1(n_975),
.B2(n_944),
.C(n_963),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1080),
.A2(n_975),
.B1(n_974),
.B2(n_963),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1088),
.A2(n_975),
.B(n_960),
.C(n_900),
.Y(n_1107)
);

OAI211xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1089),
.A2(n_16),
.B(n_19),
.C(n_20),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1086),
.B(n_978),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1081),
.Y(n_1110)
);

AOI221x1_ASAP7_75t_L g1111 ( 
.A1(n_1094),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.C(n_22),
.Y(n_1111)
);

AOI211xp5_ASAP7_75t_L g1112 ( 
.A1(n_1092),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1079),
.B(n_978),
.Y(n_1113)
);

OAI221xp5_ASAP7_75t_L g1114 ( 
.A1(n_1083),
.A2(n_949),
.B1(n_836),
.B2(n_828),
.C(n_879),
.Y(n_1114)
);

AOI221x1_ASAP7_75t_L g1115 ( 
.A1(n_1079),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.C(n_28),
.Y(n_1115)
);

AOI211xp5_ASAP7_75t_L g1116 ( 
.A1(n_1079),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1078),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1078),
.Y(n_1118)
);

AND4x1_ASAP7_75t_L g1119 ( 
.A(n_1116),
.B(n_29),
.C(n_30),
.D(n_31),
.Y(n_1119)
);

AOI221xp5_ASAP7_75t_L g1120 ( 
.A1(n_1116),
.A2(n_1097),
.B1(n_1117),
.B2(n_1098),
.C(n_1118),
.Y(n_1120)
);

OAI211xp5_ASAP7_75t_SL g1121 ( 
.A1(n_1110),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_1121)
);

AOI222xp33_ASAP7_75t_L g1122 ( 
.A1(n_1108),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.C1(n_38),
.C2(n_39),
.Y(n_1122)
);

AOI221xp5_ASAP7_75t_L g1123 ( 
.A1(n_1100),
.A2(n_963),
.B1(n_944),
.B2(n_40),
.C(n_41),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1115),
.B(n_978),
.Y(n_1124)
);

AOI221xp5_ASAP7_75t_L g1125 ( 
.A1(n_1096),
.A2(n_963),
.B1(n_36),
.B2(n_41),
.C(n_42),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1113),
.A2(n_949),
.B1(n_879),
.B2(n_828),
.Y(n_1126)
);

XOR2xp5_ASAP7_75t_L g1127 ( 
.A(n_1101),
.B(n_32),
.Y(n_1127)
);

OAI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1104),
.A2(n_879),
.B1(n_900),
.B2(n_907),
.C(n_878),
.Y(n_1128)
);

AOI311xp33_ASAP7_75t_L g1129 ( 
.A1(n_1114),
.A2(n_42),
.A3(n_43),
.B(n_44),
.C(n_45),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_1109),
.Y(n_1130)
);

AOI21xp33_ASAP7_75t_L g1131 ( 
.A1(n_1112),
.A2(n_43),
.B(n_44),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1095),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.C(n_50),
.Y(n_1132)
);

AOI211xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1106),
.A2(n_46),
.B(n_50),
.C(n_51),
.Y(n_1133)
);

AO22x1_ASAP7_75t_L g1134 ( 
.A1(n_1102),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1134)
);

OAI211xp5_ASAP7_75t_SL g1135 ( 
.A1(n_1105),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1099),
.B(n_981),
.Y(n_1136)
);

OAI311xp33_ASAP7_75t_L g1137 ( 
.A1(n_1107),
.A2(n_56),
.A3(n_58),
.B1(n_59),
.C1(n_907),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1103),
.B(n_932),
.Y(n_1138)
);

OAI322xp33_ASAP7_75t_L g1139 ( 
.A1(n_1111),
.A2(n_59),
.A3(n_878),
.B1(n_961),
.B2(n_960),
.C1(n_912),
.C2(n_981),
.Y(n_1139)
);

AOI221xp5_ASAP7_75t_L g1140 ( 
.A1(n_1116),
.A2(n_972),
.B1(n_981),
.B2(n_960),
.C(n_961),
.Y(n_1140)
);

AOI211xp5_ASAP7_75t_L g1141 ( 
.A1(n_1097),
.A2(n_972),
.B(n_938),
.C(n_907),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1113),
.Y(n_1142)
);

NAND3x1_ASAP7_75t_L g1143 ( 
.A(n_1119),
.B(n_907),
.C(n_897),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1130),
.Y(n_1144)
);

AO22x2_ASAP7_75t_L g1145 ( 
.A1(n_1142),
.A2(n_1127),
.B1(n_1138),
.B2(n_1124),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1134),
.Y(n_1146)
);

XNOR2xp5_ASAP7_75t_L g1147 ( 
.A(n_1120),
.B(n_1125),
.Y(n_1147)
);

NOR2x1_ASAP7_75t_L g1148 ( 
.A(n_1121),
.B(n_391),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1136),
.B(n_938),
.Y(n_1149)
);

OAI322xp33_ASAP7_75t_L g1150 ( 
.A1(n_1126),
.A2(n_1137),
.A3(n_1132),
.B1(n_1129),
.B2(n_1123),
.C1(n_1128),
.C2(n_1133),
.Y(n_1150)
);

NAND4xp75_ASAP7_75t_L g1151 ( 
.A(n_1131),
.B(n_929),
.C(n_897),
.D(n_885),
.Y(n_1151)
);

NAND4xp75_ASAP7_75t_L g1152 ( 
.A(n_1140),
.B(n_929),
.C(n_899),
.D(n_894),
.Y(n_1152)
);

NOR2x1_ASAP7_75t_L g1153 ( 
.A(n_1139),
.B(n_391),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_1122),
.B(n_62),
.Y(n_1154)
);

NOR3xp33_ASAP7_75t_L g1155 ( 
.A(n_1135),
.B(n_899),
.C(n_391),
.Y(n_1155)
);

XOR2x1_ASAP7_75t_L g1156 ( 
.A(n_1122),
.B(n_64),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1141),
.A2(n_899),
.B(n_911),
.Y(n_1157)
);

XOR2x1_ASAP7_75t_L g1158 ( 
.A(n_1142),
.B(n_65),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1130),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1130),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1135),
.A2(n_879),
.B1(n_887),
.B2(n_911),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1130),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1130),
.B(n_911),
.Y(n_1163)
);

XNOR2x1_ASAP7_75t_L g1164 ( 
.A(n_1142),
.B(n_72),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1145),
.A2(n_915),
.B(n_911),
.Y(n_1165)
);

AOI222xp33_ASAP7_75t_L g1166 ( 
.A1(n_1154),
.A2(n_915),
.B1(n_883),
.B2(n_882),
.C1(n_887),
.C2(n_85),
.Y(n_1166)
);

AOI322xp5_ASAP7_75t_L g1167 ( 
.A1(n_1146),
.A2(n_883),
.A3(n_882),
.B1(n_887),
.B2(n_891),
.C1(n_886),
.C2(n_89),
.Y(n_1167)
);

AOI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1150),
.A2(n_887),
.B1(n_883),
.B2(n_882),
.C(n_891),
.Y(n_1168)
);

NOR3xp33_ASAP7_75t_L g1169 ( 
.A(n_1144),
.B(n_1159),
.C(n_1160),
.Y(n_1169)
);

OAI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1162),
.A2(n_887),
.B1(n_883),
.B2(n_882),
.Y(n_1170)
);

AOI221xp5_ASAP7_75t_L g1171 ( 
.A1(n_1145),
.A2(n_891),
.B1(n_886),
.B2(n_82),
.C(n_84),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1147),
.B(n_76),
.C(n_77),
.Y(n_1172)
);

NOR2x1_ASAP7_75t_L g1173 ( 
.A(n_1164),
.B(n_391),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1148),
.B(n_400),
.C(n_396),
.Y(n_1174)
);

NOR3xp33_ASAP7_75t_L g1175 ( 
.A(n_1153),
.B(n_391),
.C(n_396),
.Y(n_1175)
);

AND3x4_ASAP7_75t_L g1176 ( 
.A(n_1155),
.B(n_891),
.C(n_886),
.Y(n_1176)
);

OAI221xp5_ASAP7_75t_L g1177 ( 
.A1(n_1161),
.A2(n_886),
.B1(n_903),
.B2(n_96),
.C(n_97),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_SL g1178 ( 
.A(n_1156),
.B(n_87),
.C(n_90),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1158),
.B(n_99),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1179),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1173),
.Y(n_1181)
);

XNOR2xp5_ASAP7_75t_L g1182 ( 
.A(n_1178),
.B(n_1143),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1169),
.B(n_1163),
.Y(n_1183)
);

OAI22x1_ASAP7_75t_L g1184 ( 
.A1(n_1176),
.A2(n_1149),
.B1(n_1151),
.B2(n_1152),
.Y(n_1184)
);

OA22x2_ASAP7_75t_L g1185 ( 
.A1(n_1172),
.A2(n_1157),
.B1(n_103),
.B2(n_106),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1171),
.A2(n_903),
.B(n_896),
.Y(n_1186)
);

OAI22x1_ASAP7_75t_L g1187 ( 
.A1(n_1174),
.A2(n_903),
.B1(n_108),
.B2(n_110),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1177),
.A2(n_903),
.B1(n_400),
.B2(n_506),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1175),
.Y(n_1189)
);

OAI211xp5_ASAP7_75t_L g1190 ( 
.A1(n_1167),
.A2(n_100),
.B(n_112),
.C(n_114),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1165),
.B(n_115),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1168),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1170),
.Y(n_1193)
);

OAI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1166),
.A2(n_903),
.B1(n_122),
.B2(n_125),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1183),
.A2(n_118),
.B1(n_127),
.B2(n_132),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1180),
.A2(n_903),
.B1(n_896),
.B2(n_400),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1192),
.A2(n_896),
.B1(n_400),
.B2(n_509),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1182),
.Y(n_1198)
);

OAI22x1_ASAP7_75t_L g1199 ( 
.A1(n_1193),
.A2(n_135),
.B1(n_136),
.B2(n_140),
.Y(n_1199)
);

AO22x2_ASAP7_75t_L g1200 ( 
.A1(n_1181),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_1200)
);

AO22x2_ASAP7_75t_L g1201 ( 
.A1(n_1189),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1185),
.A2(n_1190),
.B1(n_1191),
.B2(n_1184),
.Y(n_1202)
);

OAI22x1_ASAP7_75t_L g1203 ( 
.A1(n_1187),
.A2(n_156),
.B1(n_157),
.B2(n_160),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1194),
.A2(n_896),
.B1(n_400),
.B2(n_482),
.Y(n_1204)
);

XNOR2xp5_ASAP7_75t_L g1205 ( 
.A(n_1202),
.B(n_1188),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1201),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1198),
.A2(n_1186),
.B(n_811),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1199),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1204),
.A2(n_512),
.B1(n_509),
.B2(n_507),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1200),
.B(n_163),
.Y(n_1210)
);

AOI22x1_ASAP7_75t_L g1211 ( 
.A1(n_1206),
.A2(n_1203),
.B1(n_1195),
.B2(n_1197),
.Y(n_1211)
);

NAND2x1p5_ASAP7_75t_L g1212 ( 
.A(n_1208),
.B(n_1196),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1210),
.B(n_169),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1205),
.A2(n_482),
.B1(n_512),
.B2(n_509),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1212),
.A2(n_1207),
.B1(n_1209),
.B2(n_175),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1215),
.B(n_1213),
.Y(n_1216)
);

AO22x2_ASAP7_75t_L g1217 ( 
.A1(n_1216),
.A2(n_1214),
.B1(n_1211),
.B2(n_176),
.Y(n_1217)
);

XNOR2xp5_ASAP7_75t_L g1218 ( 
.A(n_1217),
.B(n_171),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1218),
.A2(n_485),
.B1(n_507),
.B2(n_506),
.Y(n_1219)
);

AOI211xp5_ASAP7_75t_L g1220 ( 
.A1(n_1219),
.A2(n_172),
.B(n_177),
.C(n_178),
.Y(n_1220)
);


endmodule