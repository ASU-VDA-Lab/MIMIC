module fake_jpeg_4197_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_14),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_24),
.Y(n_73)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_30),
.B1(n_22),
.B2(n_15),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_30),
.B1(n_15),
.B2(n_22),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_23),
.C(n_16),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_64),
.B1(n_30),
.B2(n_22),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_25),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_30),
.B1(n_22),
.B2(n_15),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_43),
.B1(n_52),
.B2(n_65),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_81),
.B1(n_48),
.B2(n_57),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_76),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_80),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_38),
.B1(n_29),
.B2(n_24),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_41),
.B1(n_23),
.B2(n_25),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_48),
.B1(n_57),
.B2(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_49),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_98),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_58),
.CI(n_44),
.CON(n_93),
.SN(n_93)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_88),
.Y(n_133)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_111),
.Y(n_124)
);

HB1xp67_ASAP7_75t_SL g97 ( 
.A(n_66),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_103),
.B(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_86),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_55),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_42),
.C(n_53),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_26),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_61),
.B(n_54),
.C(n_48),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_116),
.B1(n_72),
.B2(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_115),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_29),
.B(n_16),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_41),
.B1(n_33),
.B2(n_29),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_37),
.B(n_31),
.C(n_28),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_63),
.B1(n_16),
.B2(n_18),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_122),
.B(n_130),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_90),
.B1(n_84),
.B2(n_82),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_125),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_101),
.B1(n_94),
.B2(n_140),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_72),
.B1(n_88),
.B2(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_78),
.Y(n_129)
);

OR2x2_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_14),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_91),
.B(n_47),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_47),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_91),
.A2(n_37),
.B(n_31),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_117),
.C(n_122),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_114),
.B1(n_93),
.B2(n_104),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_105),
.B1(n_108),
.B2(n_99),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_93),
.A2(n_37),
.B(n_31),
.C(n_28),
.D(n_26),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_116),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_98),
.B(n_0),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_87),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_103),
.C(n_95),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_154),
.C(n_133),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_157),
.B(n_26),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_102),
.Y(n_151)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_102),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_155),
.A2(n_121),
.B(n_130),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_168),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_108),
.Y(n_162)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_143),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_101),
.B1(n_112),
.B2(n_115),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_19),
.B1(n_18),
.B2(n_28),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_124),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_28),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_152),
.B(n_156),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_158),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_185),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_119),
.C(n_126),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_182),
.C(n_187),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_136),
.B1(n_128),
.B2(n_138),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_179),
.B1(n_144),
.B2(n_165),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_87),
.Y(n_178)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_143),
.B1(n_121),
.B2(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_186),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_189),
.B(n_193),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_141),
.C(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_192),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_121),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_28),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_158),
.A2(n_19),
.B1(n_18),
.B2(n_26),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_196),
.B1(n_149),
.B2(n_147),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_20),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_148),
.A2(n_28),
.B(n_20),
.C(n_19),
.D(n_18),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_160),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_204),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_202),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_163),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_217),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_169),
.C(n_163),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.C(n_211),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_151),
.C(n_153),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_193),
.B1(n_183),
.B2(n_175),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_153),
.C(n_144),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_145),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_214),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_145),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_177),
.B(n_186),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_182),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_20),
.C(n_14),
.Y(n_236)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_193),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_218),
.B(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_238),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_194),
.B1(n_155),
.B2(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_225),
.A2(n_226),
.B1(n_205),
.B2(n_224),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_149),
.B1(n_184),
.B2(n_160),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_202),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_235),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_20),
.B(n_2),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_239),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_20),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_20),
.C(n_2),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_206),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_222),
.B1(n_221),
.B2(n_227),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_201),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_256),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_207),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_208),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_259),
.C(n_198),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_225),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_258),
.B(n_228),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_268),
.C(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_266),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_241),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_264),
.B(n_3),
.Y(n_287)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_236),
.B(n_234),
.C(n_240),
.D(n_13),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_1),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_13),
.B(n_12),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_246),
.A2(n_244),
.B(n_251),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_252),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_12),
.B(n_10),
.C(n_9),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_273),
.A2(n_274),
.B(n_1),
.Y(n_276)
);

OAI321xp33_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_12),
.A3(n_9),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_274)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_259),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_286),
.C(n_269),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_281),
.B(n_284),
.Y(n_288)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_273),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_268),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_2),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_287),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_280),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_295),
.B(n_296),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_4),
.B(n_5),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_4),
.B(n_5),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_4),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_282),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_304),
.B(n_290),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_279),
.B1(n_7),
.B2(n_8),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_6),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_299),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_301),
.B(n_298),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_312),
.C(n_306),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_292),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.C(n_311),
.Y(n_315)
);

AO21x2_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_308),
.B(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_8),
.Y(n_317)
);


endmodule