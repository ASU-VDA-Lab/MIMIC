module fake_jpeg_28205_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_SL g10 ( 
.A(n_7),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_18),
.B(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_9),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_13),
.C(n_8),
.Y(n_33)
);

NOR2xp67_ASAP7_75t_R g31 ( 
.A(n_30),
.B(n_9),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_17),
.B1(n_26),
.B2(n_11),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_11),
.B1(n_3),
.B2(n_2),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_19),
.C(n_25),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_19),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_15),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_8),
.B(n_13),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_13),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_36),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_40),
.C(n_39),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_37),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_50),
.C(n_42),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_44),
.B1(n_4),
.B2(n_5),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_43),
.B(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_4),
.B1(n_6),
.B2(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_54),
.Y(n_58)
);


endmodule