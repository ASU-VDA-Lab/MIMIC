module fake_jpeg_30225_n_96 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_37),
.B1(n_28),
.B2(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_51),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_35),
.B1(n_36),
.B2(n_34),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_28),
.B(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_1),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_52),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_27),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_70),
.B1(n_53),
.B2(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_3),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_57),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_68),
.B(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_81),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_80),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_57),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

AOI21x1_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_87),
.B(n_85),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_76),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_74),
.B(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_72),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_4),
.C(n_12),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_4),
.B(n_8),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_93),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_16),
.B(n_20),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_21),
.Y(n_96)
);


endmodule