module fake_netlist_6_2216_n_1719 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_190, n_262, n_187, n_60, n_361, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1719);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1719;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_1697;
wire n_979;
wire n_905;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_1664;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_527;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1617;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_576;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1632;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_277),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_16),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_224),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_341),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_310),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_364),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_61),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_164),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_70),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_371),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_122),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_311),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_140),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_301),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_69),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_56),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_15),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_114),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_158),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_177),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_270),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_355),
.Y(n_398)
);

BUFx10_ASAP7_75t_L g399 ( 
.A(n_176),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_285),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_119),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_204),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_186),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_375),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_278),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_127),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_324),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_232),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_209),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_351),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_154),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_93),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_257),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_256),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_4),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_124),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_77),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_316),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_141),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_296),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_288),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_42),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_88),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_68),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_243),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_208),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_147),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_212),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_98),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_136),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_346),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_269),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_35),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_170),
.Y(n_437)
);

INVx4_ASAP7_75t_R g438 ( 
.A(n_321),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_193),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_132),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_242),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_357),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_263),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_290),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_54),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_326),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_56),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_91),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_262),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_94),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_354),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_62),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_61),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_78),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_29),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_292),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_138),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_342),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_57),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_19),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_139),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_312),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_18),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_96),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_205),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_331),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_104),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_356),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_72),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_82),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_240),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_210),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_25),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_272),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_151),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_309),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_336),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_226),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_15),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_343),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_89),
.Y(n_482)
);

CKINVDCx14_ASAP7_75t_R g483 ( 
.A(n_228),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_298),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_246),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_9),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_332),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_115),
.Y(n_488)
);

BUFx10_ASAP7_75t_L g489 ( 
.A(n_137),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_366),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_362),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_175),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_130),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_198),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_329),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_16),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_152),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_289),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_111),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_23),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_215),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_118),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_161),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_293),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_17),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_216),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_83),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_123),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_249),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_237),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_282),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_245),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_35),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_370),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_303),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_184),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_274),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_317),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_109),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_268),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_340),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_199),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_50),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_338),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_172),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_159),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_267),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_238),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_229),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_43),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_3),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_128),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_352),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_13),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_248),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_291),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_368),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_144),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_211),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_353),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_218),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_102),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_100),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_81),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_253),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_280),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_302),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_227),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_148),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_234),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_173),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_284),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_259),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_275),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_206),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_363),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_146),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_182),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_347),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_180),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_108),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_192),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_160),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_143),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_112),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_273),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_156),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_79),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_306),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_325),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_369),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_34),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_244),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_133),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_217),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_276),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_121),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_135),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_344),
.Y(n_579)
);

BUFx5_ASAP7_75t_L g580 ( 
.A(n_335),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_169),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_116),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_300),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_233),
.Y(n_584)
);

BUFx8_ASAP7_75t_SL g585 ( 
.A(n_70),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_223),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_54),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_266),
.Y(n_588)
);

HB1xp67_ASAP7_75t_SL g589 ( 
.A(n_62),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_2),
.Y(n_590)
);

INVx4_ASAP7_75t_R g591 ( 
.A(n_44),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_190),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_213),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_166),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_348),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_304),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_327),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_131),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_307),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_333),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_251),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_203),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_196),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_281),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_110),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_197),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_287),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_157),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_92),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_207),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_167),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_31),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_505),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_585),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_580),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_585),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_460),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_474),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_546),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_376),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_379),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_384),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_474),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_400),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_388),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_514),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_397),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_387),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_393),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_420),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_389),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_395),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_427),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_396),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_393),
.Y(n_636)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_478),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_393),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_466),
.B(n_0),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_L g640 ( 
.A(n_572),
.B(n_0),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_440),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_393),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_398),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_392),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_599),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_377),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_436),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_R g648 ( 
.A(n_483),
.B(n_80),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_445),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_589),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_400),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_453),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_466),
.B(n_1),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_402),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_404),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_382),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_405),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_412),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_414),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_414),
.Y(n_660)
);

CKINVDCx16_ASAP7_75t_R g661 ( 
.A(n_555),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_413),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_462),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_454),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_415),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_462),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_542),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_418),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_382),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_461),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_383),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_580),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_470),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_486),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_515),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_391),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_452),
.B(n_1),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_416),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_513),
.Y(n_679)
);

CKINVDCx16_ASAP7_75t_R g680 ( 
.A(n_483),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_580),
.Y(n_681)
);

INVxp67_ASAP7_75t_SL g682 ( 
.A(n_515),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_531),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_534),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_587),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_520),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_590),
.Y(n_687)
);

INVxp67_ASAP7_75t_SL g688 ( 
.A(n_520),
.Y(n_688)
);

INVxp33_ASAP7_75t_SL g689 ( 
.A(n_424),
.Y(n_689)
);

INVxp33_ASAP7_75t_L g690 ( 
.A(n_385),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_612),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_538),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_426),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_538),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_419),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_407),
.B(n_2),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_378),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_380),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_428),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_464),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_R g701 ( 
.A(n_431),
.B(n_433),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_604),
.B(n_421),
.Y(n_702)
);

CKINVDCx16_ASAP7_75t_R g703 ( 
.A(n_447),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_447),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_381),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_480),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_386),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_441),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_394),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_421),
.B(n_3),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_401),
.Y(n_711)
);

INVxp33_ASAP7_75t_SL g712 ( 
.A(n_496),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_500),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_442),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_R g715 ( 
.A(n_443),
.B(n_4),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_530),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_403),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_406),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_447),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_408),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_410),
.Y(n_721)
);

INVxp33_ASAP7_75t_SL g722 ( 
.A(n_523),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_444),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_411),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_417),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_446),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_580),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_580),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_422),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_580),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_448),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_423),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_425),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_449),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_450),
.B(n_5),
.Y(n_735)
);

CKINVDCx16_ASAP7_75t_R g736 ( 
.A(n_399),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_450),
.B(n_5),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_429),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_451),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_455),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_430),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_432),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_457),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_459),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_434),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_399),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_465),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_467),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_435),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_468),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_473),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_475),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_479),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_493),
.B(n_6),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_437),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_481),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_456),
.Y(n_757)
);

CKINVDCx16_ASAP7_75t_R g758 ( 
.A(n_399),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_439),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_385),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_485),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_487),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_490),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_580),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_524),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_491),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_492),
.Y(n_767)
);

INVxp33_ASAP7_75t_SL g768 ( 
.A(n_494),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_493),
.B(n_6),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_502),
.B(n_7),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_489),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_489),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_458),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_626),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_630),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_636),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_621),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_765),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_638),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_628),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_765),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_642),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_722),
.A2(n_409),
.B1(n_521),
.B2(n_390),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_R g784 ( 
.A(n_700),
.B(n_7),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_615),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_656),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_746),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_656),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_746),
.B(n_502),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_622),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_680),
.B(n_489),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_615),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_760),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_644),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_647),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_697),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_623),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_639),
.B(n_525),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_698),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_619),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_686),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_629),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_646),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_632),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_705),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_686),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_707),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_672),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_631),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_672),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_633),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_635),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_643),
.B(n_508),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_654),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_655),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_657),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_658),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_681),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_709),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_704),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_711),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_650),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_717),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_662),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_649),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_652),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_640),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_665),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_664),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_718),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_627),
.B(n_525),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_670),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_669),
.B(n_508),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_720),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_721),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_673),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_668),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_757),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_R g839 ( 
.A(n_695),
.B(n_495),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_724),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_613),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_725),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_674),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_699),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_634),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_653),
.B(n_525),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_616),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_708),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_714),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_726),
.B(n_545),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_681),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_727),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_729),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_692),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_671),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_732),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_679),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_733),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_738),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_694),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_741),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_667),
.B(n_543),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_742),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_745),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_683),
.Y(n_865)
);

CKINVDCx16_ASAP7_75t_R g866 ( 
.A(n_736),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_749),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_684),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_641),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_755),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_731),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_759),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_773),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_685),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_624),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_739),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_687),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_691),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_743),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_727),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_675),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_822),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_796),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_799),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_805),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_786),
.B(n_682),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_786),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_807),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_880),
.Y(n_889)
);

INVx4_ASAP7_75t_L g890 ( 
.A(n_788),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_819),
.Y(n_891)
);

BUFx10_ASAP7_75t_L g892 ( 
.A(n_777),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_880),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_788),
.B(n_688),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_798),
.B(n_768),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_778),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_798),
.B(n_689),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_790),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_801),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_801),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_820),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_785),
.B(n_792),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_806),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_822),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_846),
.B(n_712),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_821),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_783),
.A2(n_846),
.B1(n_620),
.B2(n_772),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_778),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_791),
.B(n_637),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_813),
.B(n_744),
.Y(n_910)
);

OAI21xp33_ASAP7_75t_L g911 ( 
.A1(n_833),
.A2(n_735),
.B(n_710),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_787),
.B(n_661),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_823),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_850),
.B(n_747),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_806),
.B(n_769),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_839),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_778),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_839),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_830),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_778),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_834),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_833),
.A2(n_702),
.B1(n_770),
.B2(n_754),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_793),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_797),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_876),
.B(n_558),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_794),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_881),
.A2(n_737),
.B1(n_696),
.B2(n_677),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_781),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_831),
.B(n_758),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_785),
.B(n_728),
.Y(n_930)
);

NAND3xp33_ASAP7_75t_L g931 ( 
.A(n_854),
.B(n_553),
.C(n_545),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_835),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_840),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_789),
.B(n_463),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_842),
.Y(n_935)
);

INVx4_ASAP7_75t_SL g936 ( 
.A(n_789),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_827),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_781),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_802),
.B(n_748),
.Y(n_939)
);

INVx4_ASAP7_75t_SL g940 ( 
.A(n_862),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_792),
.B(n_808),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_804),
.B(n_751),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_853),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_811),
.B(n_752),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_781),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_856),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_781),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_858),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_808),
.B(n_728),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_859),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_779),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_861),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_800),
.B(n_753),
.Y(n_953)
);

AO21x2_ASAP7_75t_L g954 ( 
.A1(n_810),
.A2(n_648),
.B(n_701),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_782),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_803),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_793),
.B(n_761),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_838),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_863),
.Y(n_959)
);

AND2x2_ASAP7_75t_SL g960 ( 
.A(n_866),
.B(n_703),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_864),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_838),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_810),
.B(n_818),
.Y(n_963)
);

AND2x6_ASAP7_75t_L g964 ( 
.A(n_875),
.B(n_553),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_812),
.B(n_762),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_854),
.A2(n_690),
.B1(n_564),
.B2(n_607),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_794),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_818),
.B(n_730),
.Y(n_968)
);

INVx8_ASAP7_75t_L g969 ( 
.A(n_814),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_827),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_794),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_775),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_851),
.B(n_730),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_815),
.B(n_766),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_867),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_816),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_870),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_800),
.B(n_767),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_860),
.B(n_841),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_851),
.B(n_764),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_843),
.B(n_597),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_872),
.Y(n_982)
);

INVxp67_ASAP7_75t_SL g983 ( 
.A(n_860),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_883),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_895),
.B(n_817),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_911),
.A2(n_584),
.B1(n_607),
.B2(n_564),
.Y(n_986)
);

OAI221xp5_ASAP7_75t_L g987 ( 
.A1(n_922),
.A2(n_784),
.B1(n_841),
.B2(n_847),
.C(n_873),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_902),
.B(n_852),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_902),
.B(n_852),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_910),
.B(n_824),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_941),
.B(n_847),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_898),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_897),
.B(n_905),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_941),
.B(n_764),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_884),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_885),
.Y(n_996)
);

INVx8_ASAP7_75t_L g997 ( 
.A(n_969),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_953),
.B(n_828),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_901),
.B(n_803),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_887),
.B(n_837),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_907),
.B(n_855),
.C(n_617),
.Y(n_1001)
);

OAI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_907),
.A2(n_914),
.B1(n_923),
.B2(n_978),
.Y(n_1002)
);

AND2x6_ASAP7_75t_SL g1003 ( 
.A(n_939),
.B(n_469),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_889),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_927),
.A2(n_772),
.B1(n_771),
.B2(n_690),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_903),
.A2(n_776),
.B(n_825),
.Y(n_1006)
);

NOR2xp67_ASAP7_75t_L g1007 ( 
.A(n_942),
.B(n_844),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_888),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_911),
.A2(n_584),
.B(n_471),
.C(n_476),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_887),
.B(n_848),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_899),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_889),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_891),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_958),
.B(n_614),
.Y(n_1014)
);

BUFx8_ASAP7_75t_L g1015 ( 
.A(n_962),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_900),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_934),
.A2(n_472),
.B1(n_482),
.B2(n_477),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_890),
.B(n_886),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_890),
.B(n_849),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_906),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_886),
.B(n_871),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_893),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_957),
.B(n_879),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_936),
.B(n_836),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_963),
.B(n_843),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_969),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_967),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_893),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_937),
.B(n_723),
.Y(n_1029)
);

INVx8_ASAP7_75t_L g1030 ( 
.A(n_969),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_958),
.B(n_645),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_894),
.B(n_734),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_913),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_894),
.B(n_740),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_963),
.B(n_865),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_882),
.B(n_865),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_930),
.B(n_868),
.Y(n_1037)
);

AND2x2_ASAP7_75t_SL g1038 ( 
.A(n_960),
.B(n_916),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_L g1039 ( 
.A(n_964),
.B(n_498),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_904),
.B(n_877),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_970),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_930),
.B(n_794),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_934),
.A2(n_484),
.B1(n_497),
.B2(n_488),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_940),
.B(n_750),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_915),
.B(n_756),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_915),
.B(n_763),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_919),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_956),
.B(n_771),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_967),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_964),
.A2(n_517),
.B1(n_526),
.B2(n_511),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_918),
.B(n_533),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_940),
.B(n_671),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_954),
.B(n_795),
.Y(n_1053)
);

AND2x6_ASAP7_75t_SL g1054 ( 
.A(n_944),
.B(n_539),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_951),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_954),
.B(n_795),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_979),
.B(n_676),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_955),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_979),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_972),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_924),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_921),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_936),
.B(n_676),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_983),
.B(n_678),
.Y(n_1064)
);

NAND2x1_ASAP7_75t_L g1065 ( 
.A(n_896),
.B(n_938),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_932),
.B(n_795),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_948),
.B(n_878),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_933),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_929),
.A2(n_693),
.B1(n_706),
.B2(n_678),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_964),
.A2(n_540),
.B1(n_551),
.B2(n_541),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_974),
.B(n_774),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_965),
.B(n_693),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_935),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_943),
.A2(n_567),
.B(n_575),
.C(n_568),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_981),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_946),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_950),
.B(n_961),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_952),
.B(n_795),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_925),
.B(n_780),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_975),
.B(n_826),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_977),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_959),
.B(n_706),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_909),
.B(n_713),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_892),
.B(n_713),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_982),
.B(n_716),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_SL g1086 ( 
.A(n_976),
.B(n_543),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_908),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_908),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_892),
.B(n_716),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_967),
.B(n_826),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_912),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1076),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1016),
.B(n_931),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_R g1094 ( 
.A(n_1061),
.B(n_809),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_993),
.B(n_651),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_1041),
.B(n_931),
.Y(n_1096)
);

OR2x6_ASAP7_75t_L g1097 ( 
.A(n_997),
.B(n_1030),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1055),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1011),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_SL g1100 ( 
.A(n_1086),
.B(n_625),
.C(n_659),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1002),
.B(n_971),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_986),
.A2(n_964),
.B1(n_577),
.B2(n_579),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_999),
.B(n_660),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_984),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1058),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_995),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_996),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_1011),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1008),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1025),
.B(n_949),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_990),
.A2(n_998),
.B(n_1009),
.C(n_1025),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1013),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_992),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1035),
.B(n_949),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_R g1115 ( 
.A(n_997),
.B(n_845),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1036),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1020),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1033),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1087),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1011),
.B(n_869),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1035),
.B(n_968),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1047),
.Y(n_1122)
);

INVxp33_ASAP7_75t_SL g1123 ( 
.A(n_1031),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1062),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1059),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1068),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1088),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1073),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1037),
.B(n_968),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1081),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1077),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_987),
.A2(n_625),
.B1(n_666),
.B2(n_663),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_997),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1040),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_R g1135 ( 
.A(n_1030),
.B(n_618),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1037),
.B(n_973),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1015),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1026),
.Y(n_1138)
);

NAND2x1_ASAP7_75t_L g1139 ( 
.A(n_1027),
.B(n_896),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1060),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1004),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_991),
.B(n_973),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1041),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_991),
.B(n_980),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1007),
.B(n_971),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1012),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1022),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1018),
.B(n_971),
.Y(n_1148)
);

BUFx12f_ASAP7_75t_L g1149 ( 
.A(n_1015),
.Y(n_1149)
);

XNOR2xp5_ASAP7_75t_L g1150 ( 
.A(n_1038),
.B(n_618),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_SL g1151 ( 
.A(n_1005),
.B(n_784),
.C(n_715),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1028),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1024),
.B(n_917),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1042),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_994),
.B(n_980),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1024),
.B(n_920),
.Y(n_1156)
);

BUFx4f_ASAP7_75t_L g1157 ( 
.A(n_1030),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1066),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_1082),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1000),
.B(n_938),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1086),
.A2(n_719),
.B1(n_578),
.B2(n_594),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1010),
.B(n_966),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_1048),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1080),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_994),
.B(n_908),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_988),
.B(n_928),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1042),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1065),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_1027),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_985),
.B(n_719),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1067),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_988),
.B(n_928),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_989),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_1079),
.B(n_588),
.Y(n_1174)
);

NOR3xp33_ASAP7_75t_SL g1175 ( 
.A(n_1005),
.B(n_1091),
.C(n_1057),
.Y(n_1175)
);

XOR2xp5_ASAP7_75t_L g1176 ( 
.A(n_1069),
.B(n_499),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1049),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1049),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1064),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1067),
.B(n_826),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_R g1181 ( 
.A(n_1072),
.B(n_501),
.Y(n_1181)
);

O2A1O1Ixp5_ASAP7_75t_L g1182 ( 
.A1(n_1111),
.A2(n_1053),
.B(n_1056),
.C(n_1090),
.Y(n_1182)
);

NOR2x1_ASAP7_75t_SL g1183 ( 
.A(n_1097),
.B(n_1019),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1143),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1155),
.A2(n_989),
.B(n_1021),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1173),
.A2(n_1051),
.B1(n_1043),
.B2(n_1017),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1131),
.B(n_1032),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1159),
.B(n_1084),
.Y(n_1189)
);

OAI22x1_ASAP7_75t_L g1190 ( 
.A1(n_1176),
.A2(n_1083),
.B1(n_1023),
.B2(n_1085),
.Y(n_1190)
);

O2A1O1Ixp5_ASAP7_75t_L g1191 ( 
.A1(n_1101),
.A2(n_1074),
.B(n_1006),
.C(n_1078),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1165),
.A2(n_1078),
.B(n_1034),
.Y(n_1192)
);

AOI21xp33_ASAP7_75t_L g1193 ( 
.A1(n_1162),
.A2(n_1046),
.B(n_1045),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1165),
.A2(n_1051),
.B(n_1050),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1166),
.A2(n_1070),
.B(n_598),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1155),
.A2(n_1039),
.B(n_947),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_SL g1197 ( 
.A1(n_1160),
.A2(n_601),
.B(n_595),
.Y(n_1197)
);

OA22x2_ASAP7_75t_L g1198 ( 
.A1(n_1132),
.A2(n_1079),
.B1(n_1071),
.B2(n_1052),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1107),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1177),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1166),
.A2(n_1172),
.B(n_1148),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1142),
.A2(n_1029),
.B1(n_1075),
.B2(n_1079),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1144),
.B(n_1044),
.Y(n_1203)
);

BUFx8_ASAP7_75t_L g1204 ( 
.A(n_1149),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1167),
.B(n_1089),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1154),
.B(n_1014),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1110),
.A2(n_947),
.B(n_926),
.Y(n_1207)
);

NOR4xp25_ASAP7_75t_L g1208 ( 
.A(n_1161),
.B(n_603),
.C(n_611),
.D(n_610),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1129),
.B(n_1063),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1123),
.B(n_1071),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1104),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1129),
.B(n_1001),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1172),
.A2(n_945),
.B(n_928),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1110),
.A2(n_926),
.B(n_945),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1114),
.A2(n_945),
.B(n_926),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1114),
.A2(n_591),
.A3(n_1054),
.B(n_1003),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1136),
.A2(n_1071),
.B1(n_524),
.B2(n_503),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1136),
.B(n_826),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1138),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1094),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1121),
.B(n_829),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1121),
.B(n_829),
.Y(n_1222)
);

O2A1O1Ixp5_ASAP7_75t_L g1223 ( 
.A1(n_1145),
.A2(n_438),
.B(n_547),
.C(n_543),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1158),
.A2(n_506),
.B(n_504),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1164),
.B(n_829),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1139),
.A2(n_85),
.B(n_84),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1177),
.A2(n_524),
.B(n_509),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1178),
.A2(n_524),
.B(n_510),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_SL g1229 ( 
.A1(n_1093),
.A2(n_569),
.B(n_547),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1133),
.B(n_829),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_SL g1231 ( 
.A1(n_1133),
.A2(n_1169),
.B(n_1117),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1106),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1112),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1168),
.A2(n_87),
.B(n_86),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1168),
.A2(n_95),
.B(n_90),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1119),
.A2(n_99),
.B(n_97),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1118),
.B(n_832),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1119),
.A2(n_103),
.B(n_101),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1175),
.A2(n_512),
.B(n_516),
.C(n_507),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1178),
.A2(n_519),
.B(n_518),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1099),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1115),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1109),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1122),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1151),
.A2(n_527),
.B1(n_528),
.B2(n_522),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1127),
.A2(n_106),
.B(n_105),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1180),
.A2(n_532),
.B(n_529),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1179),
.B(n_832),
.Y(n_1248)
);

NAND2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1157),
.B(n_1169),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1157),
.B(n_832),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1128),
.B(n_832),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1124),
.B(n_857),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1127),
.A2(n_113),
.B(n_107),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1132),
.B(n_857),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1102),
.A2(n_536),
.B(n_535),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1185),
.A2(n_1180),
.B(n_1130),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1217),
.A2(n_1095),
.B1(n_1100),
.B2(n_1170),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1188),
.B(n_1126),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1196),
.A2(n_1182),
.B(n_1218),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1211),
.Y(n_1260)
);

CKINVDCx8_ASAP7_75t_R g1261 ( 
.A(n_1220),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1206),
.A2(n_1096),
.B1(n_1163),
.B2(n_1134),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1213),
.A2(n_1146),
.B(n_1141),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1190),
.A2(n_1150),
.B1(n_1174),
.B2(n_1137),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1215),
.A2(n_1146),
.B(n_1152),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1201),
.A2(n_1140),
.B(n_1147),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1232),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1203),
.B(n_1103),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1233),
.Y(n_1269)
);

NOR2xp67_ASAP7_75t_L g1270 ( 
.A(n_1187),
.B(n_1205),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1198),
.A2(n_1181),
.B1(n_1135),
.B2(n_1174),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1212),
.B(n_1092),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1217),
.A2(n_1098),
.A3(n_1105),
.B(n_1125),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1244),
.Y(n_1274)
);

AOI21xp33_ASAP7_75t_L g1275 ( 
.A1(n_1209),
.A2(n_1093),
.B(n_1174),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1193),
.B(n_1116),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1184),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1219),
.B(n_1097),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1248),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1199),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1242),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1193),
.A2(n_1153),
.B(n_1156),
.C(n_1171),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1243),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1204),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_SL g1285 ( 
.A1(n_1239),
.A2(n_1171),
.B(n_569),
.C(n_547),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1204),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1194),
.A2(n_1097),
.B(n_1153),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1191),
.A2(n_1156),
.B(n_544),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1192),
.A2(n_1120),
.B(n_1171),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1202),
.A2(n_1120),
.B1(n_1108),
.B2(n_1099),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1252),
.Y(n_1291)
);

AOI22x1_ASAP7_75t_L g1292 ( 
.A1(n_1197),
.A2(n_1099),
.B1(n_1108),
.B2(n_537),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1200),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1189),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1237),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1200),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1241),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1202),
.B(n_1108),
.C(n_874),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_SL g1299 ( 
.A1(n_1183),
.A2(n_120),
.B(n_117),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1236),
.A2(n_126),
.B(n_125),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1251),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1241),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1225),
.Y(n_1303)
);

AND2x4_ASAP7_75t_SL g1304 ( 
.A(n_1241),
.B(n_1113),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1221),
.A2(n_549),
.B(n_548),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1210),
.B(n_569),
.Y(n_1306)
);

CKINVDCx8_ASAP7_75t_R g1307 ( 
.A(n_1230),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1195),
.A2(n_552),
.B(n_550),
.Y(n_1308)
);

INVx8_ASAP7_75t_L g1309 ( 
.A(n_1230),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1238),
.A2(n_134),
.B(n_129),
.Y(n_1310)
);

INVxp67_ASAP7_75t_SL g1311 ( 
.A(n_1222),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1225),
.Y(n_1312)
);

BUFx12f_ASAP7_75t_L g1313 ( 
.A(n_1249),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1254),
.Y(n_1314)
);

OAI221xp5_ASAP7_75t_L g1315 ( 
.A1(n_1208),
.A2(n_878),
.B1(n_874),
.B2(n_857),
.C(n_609),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1231),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1216),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1216),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_SL g1319 ( 
.A1(n_1224),
.A2(n_214),
.B(n_271),
.C(n_265),
.Y(n_1319)
);

NOR2xp67_ASAP7_75t_L g1320 ( 
.A(n_1245),
.B(n_142),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1245),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1216),
.B(n_857),
.Y(n_1322)
);

INVx5_ASAP7_75t_L g1323 ( 
.A(n_1250),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1234),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1207),
.A2(n_556),
.B(n_554),
.Y(n_1325)
);

NAND2x1p5_ASAP7_75t_L g1326 ( 
.A(n_1226),
.B(n_874),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1224),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1208),
.A2(n_559),
.B(n_557),
.Y(n_1328)
);

AOI21xp33_ASAP7_75t_L g1329 ( 
.A1(n_1257),
.A2(n_1186),
.B(n_1223),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1327),
.A2(n_1186),
.B1(n_1255),
.B2(n_1247),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1287),
.A2(n_1253),
.B(n_1246),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1260),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1280),
.Y(n_1333)
);

BUFx2_ASAP7_75t_SL g1334 ( 
.A(n_1261),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1268),
.B(n_1240),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1258),
.B(n_1214),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1321),
.A2(n_1255),
.B1(n_1228),
.B2(n_1227),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1281),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1267),
.Y(n_1339)
);

CKINVDCx6p67_ASAP7_75t_R g1340 ( 
.A(n_1297),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1259),
.A2(n_1235),
.B(n_1229),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1294),
.B(n_874),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1258),
.B(n_560),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1264),
.A2(n_1275),
.B1(n_1271),
.B2(n_1276),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1275),
.A2(n_878),
.B1(n_608),
.B2(n_606),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1269),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1274),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1304),
.Y(n_1348)
);

NAND2xp33_ASAP7_75t_R g1349 ( 
.A(n_1278),
.B(n_561),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1277),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1283),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1279),
.B(n_562),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1309),
.Y(n_1353)
);

OAI211xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1271),
.A2(n_878),
.B(n_605),
.C(n_602),
.Y(n_1354)
);

NOR2xp67_ASAP7_75t_SL g1355 ( 
.A(n_1307),
.B(n_563),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1306),
.A2(n_600),
.B1(n_596),
.B2(n_593),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1270),
.B(n_565),
.Y(n_1357)
);

OAI211xp5_ASAP7_75t_L g1358 ( 
.A1(n_1328),
.A2(n_592),
.B(n_586),
.C(n_583),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1328),
.A2(n_582),
.B1(n_581),
.B2(n_576),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1256),
.A2(n_149),
.B(n_145),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1290),
.A2(n_574),
.B1(n_573),
.B2(n_571),
.Y(n_1361)
);

NOR3xp33_ASAP7_75t_SL g1362 ( 
.A(n_1262),
.B(n_570),
.C(n_566),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1272),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1272),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1256),
.A2(n_153),
.B(n_150),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1303),
.B(n_8),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1309),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1300),
.A2(n_162),
.B(n_155),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1314),
.B(n_8),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1278),
.B(n_163),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1293),
.Y(n_1371)
);

NAND2x1_ASAP7_75t_L g1372 ( 
.A(n_1316),
.B(n_165),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1296),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1312),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1289),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1311),
.B(n_10),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1318),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1259),
.A2(n_185),
.B(n_373),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1309),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1302),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1266),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1302),
.Y(n_1382)
);

AOI21xp33_ASAP7_75t_L g1383 ( 
.A1(n_1315),
.A2(n_12),
.B(n_14),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1266),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1289),
.B(n_168),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1311),
.B(n_14),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1315),
.A2(n_1298),
.B1(n_1282),
.B2(n_1301),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1273),
.Y(n_1388)
);

BUFx4f_ASAP7_75t_L g1389 ( 
.A(n_1313),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1273),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1273),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1295),
.B(n_17),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1317),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1291),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1322),
.Y(n_1395)
);

NOR2x1_ASAP7_75t_SL g1396 ( 
.A(n_1323),
.B(n_1298),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1320),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1284),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1344),
.B(n_1305),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1382),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1389),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1333),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1350),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1330),
.A2(n_1292),
.B1(n_1299),
.B2(n_1305),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1359),
.A2(n_1323),
.B1(n_1286),
.B2(n_1326),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1389),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1379),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1358),
.A2(n_1325),
.B1(n_1323),
.B2(n_1288),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1380),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1369),
.B(n_1325),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1339),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1346),
.Y(n_1412)
);

NAND3xp33_ASAP7_75t_L g1413 ( 
.A(n_1383),
.B(n_1319),
.C(n_1285),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1351),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1379),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1347),
.Y(n_1416)
);

AOI222xp33_ASAP7_75t_L g1417 ( 
.A1(n_1377),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.C1(n_24),
.C2(n_25),
.Y(n_1417)
);

AOI21xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1349),
.A2(n_24),
.B(n_26),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1363),
.B(n_1323),
.Y(n_1419)
);

AOI211xp5_ASAP7_75t_L g1420 ( 
.A1(n_1383),
.A2(n_1329),
.B(n_1335),
.C(n_1354),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1397),
.A2(n_1288),
.B1(n_1308),
.B2(n_1324),
.Y(n_1421)
);

AOI222xp33_ASAP7_75t_L g1422 ( 
.A1(n_1393),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.C1(n_29),
.C2(n_30),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1348),
.Y(n_1423)
);

AOI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1387),
.A2(n_1310),
.B(n_1308),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1329),
.A2(n_1324),
.B1(n_1265),
.B2(n_1263),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1353),
.B(n_1324),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1365),
.A2(n_1326),
.B(n_201),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1387),
.A2(n_200),
.B(n_372),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1365),
.A2(n_1337),
.B1(n_1376),
.B2(n_1386),
.C(n_1378),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1362),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1332),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1341),
.A2(n_202),
.B(n_367),
.Y(n_1432)
);

AOI222xp33_ASAP7_75t_L g1433 ( 
.A1(n_1343),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.C1(n_34),
.C2(n_36),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1374),
.Y(n_1434)
);

OAI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1375),
.A2(n_1376),
.B1(n_1386),
.B2(n_1364),
.Y(n_1435)
);

AOI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1392),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.C(n_37),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1357),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_1437)
);

AOI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1392),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.C(n_41),
.Y(n_1438)
);

OAI211xp5_ASAP7_75t_L g1439 ( 
.A1(n_1356),
.A2(n_1343),
.B(n_1366),
.C(n_1378),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1345),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_1440)
);

AOI222xp33_ASAP7_75t_L g1441 ( 
.A1(n_1352),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.C1(n_46),
.C2(n_47),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1394),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1370),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_1443)
);

OR2x2_ASAP7_75t_SL g1444 ( 
.A(n_1342),
.B(n_48),
.Y(n_1444)
);

AOI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1341),
.A2(n_235),
.B(n_365),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1361),
.B(n_1366),
.C(n_1336),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1340),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1370),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1334),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1385),
.B(n_171),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1336),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1373),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1353),
.B(n_174),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1371),
.B(n_1367),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1367),
.B(n_178),
.Y(n_1455)
);

CKINVDCx16_ASAP7_75t_R g1456 ( 
.A(n_1338),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1388),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1395),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1385),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1372),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1390),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1361),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_1462)
);

OAI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1398),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.C(n_63),
.Y(n_1463)
);

OAI22x1_ASAP7_75t_L g1464 ( 
.A1(n_1391),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1381),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1384),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1355),
.B(n_179),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1360),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1400),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1409),
.B(n_1331),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1403),
.B(n_1396),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1411),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1412),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1426),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1416),
.B(n_1368),
.Y(n_1475)
);

NAND2xp33_ASAP7_75t_R g1476 ( 
.A(n_1450),
.B(n_67),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1457),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1423),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1459),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1461),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1434),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1465),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1410),
.B(n_68),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1431),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1442),
.B(n_69),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1414),
.B(n_71),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1402),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1426),
.B(n_261),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1429),
.B(n_71),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1452),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1424),
.A2(n_72),
.B(n_73),
.Y(n_1491)
);

AO31x2_ASAP7_75t_L g1492 ( 
.A1(n_1427),
.A2(n_73),
.A3(n_74),
.B(n_75),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1454),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1429),
.B(n_74),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1419),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1446),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1446),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1407),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1407),
.B(n_283),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1399),
.B(n_75),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1435),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1444),
.B(n_1413),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1435),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1415),
.Y(n_1504)
);

INVx5_ASAP7_75t_L g1505 ( 
.A(n_1450),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1420),
.B(n_76),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1464),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1451),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1439),
.B(n_76),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1413),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1445),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1425),
.B(n_181),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1456),
.B(n_183),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1415),
.B(n_187),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1420),
.B(n_188),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1460),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1460),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1428),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1466),
.Y(n_1519)
);

AO21x2_ASAP7_75t_L g1520 ( 
.A1(n_1432),
.A2(n_189),
.B(n_191),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1450),
.B(n_194),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1458),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1433),
.B(n_195),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1473),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1509),
.A2(n_1463),
.B1(n_1418),
.B2(n_1447),
.C(n_1436),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1473),
.B(n_1408),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1472),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1484),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_L g1529 ( 
.A(n_1510),
.B(n_1405),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1479),
.Y(n_1530)
);

AOI222xp33_ASAP7_75t_L g1531 ( 
.A1(n_1523),
.A2(n_1438),
.B1(n_1462),
.B2(n_1440),
.C1(n_1430),
.C2(n_1437),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1481),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1470),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1477),
.B(n_1421),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1502),
.A2(n_1443),
.B1(n_1448),
.B2(n_1468),
.Y(n_1535)
);

NAND2xp33_ASAP7_75t_R g1536 ( 
.A(n_1502),
.B(n_1509),
.Y(n_1536)
);

NOR3xp33_ASAP7_75t_L g1537 ( 
.A(n_1496),
.B(n_1467),
.C(n_1449),
.Y(n_1537)
);

INVxp67_ASAP7_75t_SL g1538 ( 
.A(n_1497),
.Y(n_1538)
);

OAI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1476),
.A2(n_1441),
.B1(n_1417),
.B2(n_1422),
.C(n_1404),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1476),
.A2(n_1460),
.B1(n_1455),
.B2(n_1453),
.Y(n_1540)
);

OAI33xp33_ASAP7_75t_L g1541 ( 
.A1(n_1501),
.A2(n_1406),
.A3(n_1401),
.B1(n_1455),
.B2(n_1453),
.B3(n_225),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1515),
.A2(n_1406),
.B1(n_1401),
.B2(n_221),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1469),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1489),
.B(n_1406),
.C(n_1401),
.Y(n_1544)
);

OR2x6_ASAP7_75t_L g1545 ( 
.A(n_1518),
.B(n_219),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1480),
.B(n_220),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1516),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1495),
.B(n_222),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1474),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1505),
.A2(n_230),
.B1(n_231),
.B2(n_236),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1516),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1482),
.Y(n_1552)
);

AOI33xp33_ASAP7_75t_L g1553 ( 
.A1(n_1506),
.A2(n_374),
.A3(n_241),
.B1(n_247),
.B2(n_250),
.B3(n_252),
.Y(n_1553)
);

OAI211xp5_ASAP7_75t_L g1554 ( 
.A1(n_1506),
.A2(n_1489),
.B(n_1494),
.C(n_1503),
.Y(n_1554)
);

NOR4xp25_ASAP7_75t_SL g1555 ( 
.A(n_1507),
.B(n_239),
.C(n_254),
.D(n_255),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1487),
.Y(n_1556)
);

AOI211xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1494),
.A2(n_258),
.B(n_260),
.C(n_264),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1527),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1527),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1533),
.B(n_1493),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1524),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1543),
.B(n_1528),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1538),
.B(n_1471),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1552),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1552),
.Y(n_1565)
);

NAND2x1p5_ASAP7_75t_L g1566 ( 
.A(n_1530),
.B(n_1505),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1556),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1532),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1556),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1530),
.B(n_1474),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1549),
.B(n_1474),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1549),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1549),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1536),
.A2(n_1505),
.B1(n_1515),
.B2(n_1508),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1544),
.B(n_1505),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1526),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1526),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1534),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1534),
.B(n_1483),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1547),
.B(n_1505),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1547),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1551),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1554),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_L g1584 ( 
.A(n_1536),
.B(n_1557),
.C(n_1525),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1551),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1570),
.Y(n_1586)
);

AND2x4_ASAP7_75t_SL g1587 ( 
.A(n_1574),
.B(n_1540),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1578),
.B(n_1483),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1576),
.B(n_1537),
.Y(n_1589)
);

NAND2x1_ASAP7_75t_SL g1590 ( 
.A(n_1583),
.B(n_1529),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1577),
.B(n_1504),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1562),
.B(n_1492),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1569),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1563),
.B(n_1492),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1583),
.B(n_1500),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_L g1596 ( 
.A(n_1584),
.B(n_1553),
.C(n_1539),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1579),
.B(n_1492),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1579),
.B(n_1500),
.Y(n_1598)
);

NAND2x1p5_ASAP7_75t_L g1599 ( 
.A(n_1575),
.B(n_1498),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1575),
.A2(n_1535),
.B1(n_1531),
.B2(n_1541),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1569),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1561),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1568),
.B(n_1490),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1475),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1581),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1559),
.B(n_1491),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1571),
.B(n_1475),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1602),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1589),
.B(n_1571),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1603),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1593),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1587),
.B(n_1585),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1600),
.B(n_1565),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1601),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1596),
.A2(n_1545),
.B(n_1555),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1586),
.B(n_1585),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1600),
.B(n_1564),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1596),
.B(n_1478),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1605),
.B(n_1580),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1597),
.B(n_1567),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1588),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1598),
.Y(n_1622)
);

NAND4xp25_ASAP7_75t_L g1623 ( 
.A(n_1595),
.B(n_1553),
.C(n_1542),
.D(n_1513),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1594),
.A2(n_1519),
.B1(n_1545),
.B2(n_1522),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1607),
.B(n_1582),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1591),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1592),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1604),
.B(n_1567),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1618),
.B(n_1599),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1612),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1615),
.A2(n_1545),
.B1(n_1566),
.B2(n_1580),
.Y(n_1631)
);

OAI21xp33_ASAP7_75t_L g1632 ( 
.A1(n_1615),
.A2(n_1606),
.B(n_1545),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1611),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1613),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1611),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1618),
.B(n_1606),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1617),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1621),
.B(n_1558),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1609),
.B(n_1616),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1634),
.B(n_1622),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1633),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1637),
.B(n_1626),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_SL g1644 ( 
.A(n_1630),
.B(n_1623),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1638),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1639),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1634),
.B(n_1610),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1632),
.B(n_1629),
.Y(n_1648)
);

XNOR2x2_ASAP7_75t_L g1649 ( 
.A(n_1643),
.B(n_1631),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1642),
.B(n_1636),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1646),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1644),
.A2(n_1624),
.B(n_1614),
.Y(n_1652)
);

AOI322xp5_ASAP7_75t_L g1653 ( 
.A1(n_1648),
.A2(n_1624),
.A3(n_1627),
.B1(n_1619),
.B2(n_1608),
.C1(n_1628),
.C2(n_1625),
.Y(n_1653)
);

NAND2xp33_ASAP7_75t_SL g1654 ( 
.A(n_1640),
.B(n_1647),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_L g1655 ( 
.A(n_1641),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1645),
.B(n_1620),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_L g1657 ( 
.A(n_1654),
.B(n_1548),
.C(n_1521),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1651),
.B(n_1573),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1652),
.B(n_1521),
.Y(n_1659)
);

NOR3xp33_ASAP7_75t_L g1660 ( 
.A(n_1650),
.B(n_1550),
.C(n_1486),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1656),
.B(n_1566),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1649),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1653),
.A2(n_1580),
.B(n_1499),
.Y(n_1663)
);

NAND2xp33_ASAP7_75t_L g1664 ( 
.A(n_1655),
.B(n_1573),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_SL g1665 ( 
.A(n_1654),
.B(n_1512),
.C(n_1485),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1662),
.A2(n_1491),
.B1(n_1520),
.B2(n_1488),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_SL g1667 ( 
.A(n_1657),
.B(n_1663),
.C(n_1661),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1664),
.A2(n_1491),
.B(n_1485),
.Y(n_1668)
);

AOI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1659),
.A2(n_1658),
.B(n_1665),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1660),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1664),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1662),
.B(n_1572),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1672),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1670),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1671),
.B(n_1572),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1668),
.B(n_1558),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1667),
.B(n_1486),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1669),
.A2(n_1546),
.B1(n_1520),
.B2(n_1512),
.C(n_1488),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1666),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1671),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1667),
.A2(n_1517),
.B1(n_1516),
.B2(n_1499),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1680),
.B(n_1492),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1673),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1677),
.A2(n_1520),
.B(n_1546),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_R g1685 ( 
.A(n_1674),
.B(n_279),
.Y(n_1685)
);

NAND3x1_ASAP7_75t_L g1686 ( 
.A(n_1679),
.B(n_1517),
.C(n_1514),
.Y(n_1686)
);

NAND4xp75_ASAP7_75t_L g1687 ( 
.A(n_1681),
.B(n_1498),
.C(n_1511),
.D(n_1499),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1675),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1676),
.Y(n_1689)
);

AOI211x1_ASAP7_75t_L g1690 ( 
.A1(n_1683),
.A2(n_1678),
.B(n_1517),
.C(n_1514),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1688),
.B(n_1514),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1685),
.Y(n_1692)
);

XOR2xp5_ASAP7_75t_L g1693 ( 
.A(n_1689),
.B(n_1488),
.Y(n_1693)
);

A2O1A1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1684),
.A2(n_1511),
.B(n_294),
.C(n_295),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1682),
.Y(n_1695)
);

NAND4xp25_ASAP7_75t_L g1696 ( 
.A(n_1686),
.B(n_286),
.C(n_297),
.D(n_299),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1693),
.Y(n_1697)
);

NAND2xp33_ASAP7_75t_L g1698 ( 
.A(n_1692),
.B(n_1687),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1691),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1695),
.B(n_1694),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1690),
.B(n_305),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1696),
.Y(n_1702)
);

NAND2x1_ASAP7_75t_L g1703 ( 
.A(n_1701),
.B(n_308),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_1702),
.Y(n_1704)
);

AOI22x1_ASAP7_75t_L g1705 ( 
.A1(n_1697),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_R g1706 ( 
.A(n_1698),
.B(n_1699),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1703),
.B(n_1700),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1706),
.A2(n_1700),
.B1(n_319),
.B2(n_320),
.Y(n_1708)
);

INVxp67_ASAP7_75t_SL g1709 ( 
.A(n_1705),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1707),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1709),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1708),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_1710),
.Y(n_1713)
);

OAI21xp33_ASAP7_75t_L g1714 ( 
.A1(n_1711),
.A2(n_1704),
.B(n_322),
.Y(n_1714)
);

OAI21xp33_ASAP7_75t_L g1715 ( 
.A1(n_1712),
.A2(n_318),
.B(n_328),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1713),
.A2(n_330),
.B(n_337),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1716),
.Y(n_1717)
);

OAI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1717),
.A2(n_1714),
.B1(n_1715),
.B2(n_358),
.C(n_360),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1718),
.A2(n_345),
.B(n_349),
.C(n_361),
.Y(n_1719)
);


endmodule