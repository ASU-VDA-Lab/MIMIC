module real_jpeg_4806_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_1),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_1),
.A2(n_43),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_43),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_43),
.B1(n_100),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_2),
.A2(n_21),
.B1(n_190),
.B2(n_193),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_5),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_5),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_5),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_6),
.A2(n_115),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_6),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_6),
.A2(n_137),
.B1(n_171),
.B2(n_175),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_6),
.A2(n_137),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_6),
.A2(n_137),
.B1(n_291),
.B2(n_293),
.Y(n_290)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_7),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_7),
.Y(n_134)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_8),
.Y(n_101)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_9),
.Y(n_139)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_10),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_10),
.A2(n_52),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_10),
.A2(n_52),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_10),
.B(n_132),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_10),
.A2(n_257),
.B(n_258),
.C(n_264),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_10),
.B(n_282),
.C(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_10),
.B(n_84),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_10),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_10),
.B(n_67),
.Y(n_323)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_224),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_222),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_197),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_16),
.B(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_142),
.C(n_176),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_17),
.B(n_176),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_82),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_18),
.B(n_112),
.C(n_140),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_19),
.B(n_46),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B(n_36),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_20),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_24),
.Y(n_293)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_29),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_31),
.B(n_40),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_31),
.A2(n_181),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_31),
.B(n_181),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_31),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_36),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_36),
.B(n_289),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_37),
.Y(n_148)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_39),
.Y(n_308)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_45),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_75),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_47),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_56),
.Y(n_47)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_48),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_52),
.B(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_52),
.A2(n_115),
.B(n_158),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_52),
.A2(n_259),
.B(n_261),
.Y(n_258)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_56),
.B(n_76),
.Y(n_196)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_56),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_56),
.B(n_270),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_67),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_62),
.Y(n_282)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_66),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_66),
.Y(n_195)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_66),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_66),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_67),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_67),
.B(n_270),
.Y(n_285)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_73),
.Y(n_182)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_74),
.Y(n_292)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_74),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_75),
.A2(n_189),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_75),
.B(n_269),
.Y(n_295)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_112),
.B1(n_140),
.B2(n_141),
.Y(n_82)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_94),
.B(n_107),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_84),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_84),
.B(n_170),
.Y(n_246)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_85),
.B(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_92),
.Y(n_260)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_94),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_94),
.B(n_107),
.Y(n_212)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_95),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_104),
.Y(n_96)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_110),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_102),
.Y(n_257)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_107),
.Y(n_168)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_135),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_132),
.Y(n_144)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_119),
.B(n_205),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_132),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_127),
.B2(n_130),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_132),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_135),
.B(n_240),
.Y(n_239)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_142),
.B(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.C(n_165),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_143),
.B(n_165),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_146),
.B(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_147),
.B(n_150),
.Y(n_237)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

AOI32xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_154),
.A3(n_155),
.B1(n_157),
.B2(n_161),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_162),
.Y(n_264)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_169),
.B(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_187),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_187),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_186),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_178),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_186),
.B(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B(n_196),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_188),
.A2(n_219),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_188),
.B(n_249),
.Y(n_268)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_196),
.B(n_285),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_197),
.Y(n_361)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_213),
.CI(n_221),
.CON(n_197),
.SN(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_212),
.B(n_246),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_214),
.A2(n_220),
.B1(n_256),
.B2(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_344),
.B(n_357),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_274),
.B(n_343),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_251),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_227),
.B(n_251),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_238),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_236),
.B2(n_237),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_230),
.B(n_236),
.C(n_238),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.C(n_234),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_234),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_235),
.B(n_305),
.Y(n_320)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_239),
.B(n_242),
.C(n_248),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_265),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_252),
.B(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_255),
.A2(n_265),
.B1(n_266),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_255),
.Y(n_340)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_281),
.Y(n_280)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_337),
.B(n_342),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_327),
.B(n_336),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_299),
.B(n_326),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_286),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_286),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_284),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_280),
.B1(n_284),
.B2(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_294),
.Y(n_286)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_306),
.Y(n_305)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_297),
.C(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_309),
.B(n_325),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_303),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_321),
.B(n_324),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_320),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_330),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_333),
.C(n_334),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_341),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_341),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_353),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_346),
.B(n_347),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_350),
.C(n_351),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_353),
.A2(n_358),
.B(n_359),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_354),
.B(n_356),
.Y(n_359)
);


endmodule