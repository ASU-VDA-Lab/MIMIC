module fake_aes_11474_n_35 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_6), .B(n_8), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
NAND2x1_ASAP7_75t_L g18 ( .A(n_12), .B(n_0), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_14), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_16), .B(n_0), .Y(n_21) );
BUFx12f_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_17), .B1(n_13), .B2(n_1), .Y(n_24) );
BUFx3_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
OAI31xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_20), .A3(n_18), .B(n_2), .Y(n_26) );
INVx2_ASAP7_75t_SL g27 ( .A(n_25), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_23), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_26), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_22), .B1(n_27), .B2(n_17), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_30), .B(n_31), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_30), .B(n_22), .Y(n_33) );
AND2x4_ASAP7_75t_L g34 ( .A(n_32), .B(n_27), .Y(n_34) );
AOI222xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_33), .B1(n_5), .B2(n_7), .C1(n_9), .C2(n_3), .Y(n_35) );
endmodule