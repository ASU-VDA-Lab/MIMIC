module fake_jpeg_31591_n_479 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_479);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_479;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_51),
.Y(n_119)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_53),
.B(n_55),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_54),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_0),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_67),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_16),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_22),
.B(n_1),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_72),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_29),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_75),
.B(n_80),
.Y(n_124)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_38),
.Y(n_79)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_82),
.Y(n_105)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_94),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_90),
.Y(n_147)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_32),
.B(n_3),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_32),
.C(n_43),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_32),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_47),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_123),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_44),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_27),
.B1(n_42),
.B2(n_41),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_103),
.A2(n_109),
.B1(n_115),
.B2(n_130),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_24),
.B1(n_19),
.B2(n_40),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_24),
.B1(n_19),
.B2(n_40),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_44),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_33),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_27),
.B1(n_42),
.B2(n_41),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_63),
.B(n_43),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_20),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_22),
.B1(n_36),
.B2(n_35),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_68),
.B1(n_81),
.B2(n_107),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_52),
.A2(n_34),
.B1(n_33),
.B2(n_20),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g196 ( 
.A1(n_138),
.A2(n_139),
.B1(n_143),
.B2(n_148),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_74),
.A2(n_34),
.B1(n_36),
.B2(n_35),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_24),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_60),
.A2(n_31),
.B1(n_30),
.B2(n_47),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_62),
.A2(n_31),
.B1(n_30),
.B2(n_24),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_91),
.B(n_51),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_154),
.B(n_198),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_102),
.A2(n_83),
.B1(n_50),
.B2(n_54),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_155),
.A2(n_158),
.B1(n_202),
.B2(n_101),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_161),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_100),
.B(n_64),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_157),
.B(n_185),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_93),
.B1(n_73),
.B2(n_56),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_159),
.A2(n_160),
.B1(n_175),
.B2(n_183),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_77),
.B1(n_82),
.B2(n_69),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_162),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_165),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_95),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_121),
.B(n_90),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_172),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_95),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_87),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_70),
.B1(n_20),
.B2(n_65),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_114),
.B(n_3),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_186),
.Y(n_214)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_181),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_87),
.B1(n_65),
.B2(n_45),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_108),
.B(n_132),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_4),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_192),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_133),
.B(n_4),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_147),
.B(n_4),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_199),
.Y(n_226)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_194),
.Y(n_233)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_130),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_197),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_123),
.A2(n_5),
.B(n_6),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_128),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_150),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_119),
.Y(n_232)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_201),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_140),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_98),
.C(n_123),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_206),
.B(n_230),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_215),
.A2(n_151),
.B(n_137),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_148),
.B1(n_106),
.B2(n_146),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_216),
.A2(n_219),
.B1(n_220),
.B2(n_215),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_110),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_219),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_154),
.B(n_139),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_153),
.B(n_143),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_220),
.B(n_223),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_153),
.B(n_150),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_168),
.B(n_101),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_174),
.B(n_106),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_187),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_119),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_196),
.A2(n_146),
.B1(n_113),
.B2(n_126),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_236),
.A2(n_118),
.B1(n_189),
.B2(n_194),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_171),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_244),
.B(n_247),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_200),
.B1(n_182),
.B2(n_196),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_245),
.A2(n_125),
.B1(n_105),
.B2(n_218),
.Y(n_315)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_195),
.Y(n_247)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_249),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_174),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_227),
.C(n_225),
.Y(n_313)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_196),
.B1(n_199),
.B2(n_198),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_254),
.Y(n_299)
);

AO21x2_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_187),
.B(n_122),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_255),
.A2(n_272),
.B(n_204),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_203),
.A2(n_197),
.B1(n_181),
.B2(n_180),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_256),
.A2(n_267),
.B(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_257),
.B(n_261),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_270),
.B1(n_257),
.B2(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_205),
.B(n_191),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_162),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_262),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_217),
.B(n_131),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_274),
.Y(n_281)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_188),
.B(n_184),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_265),
.A2(n_269),
.B(n_204),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_203),
.A2(n_179),
.B1(n_173),
.B2(n_178),
.Y(n_267)
);

BUFx8_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_268),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g269 ( 
.A1(n_231),
.A2(n_152),
.B(n_169),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_213),
.A2(n_113),
.B1(n_126),
.B2(n_122),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_190),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_271),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_206),
.A2(n_201),
.B(n_105),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_213),
.B(n_176),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_279),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_230),
.B1(n_237),
.B2(n_229),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_238),
.A2(n_165),
.B1(n_166),
.B2(n_163),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_228),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_282),
.A2(n_284),
.B1(n_297),
.B2(n_269),
.Y(n_323)
);

OAI32xp33_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_223),
.A3(n_207),
.B1(n_240),
.B2(n_210),
.Y(n_283)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_253),
.A2(n_207),
.B1(n_230),
.B2(n_237),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_286),
.A2(n_277),
.B1(n_255),
.B2(n_250),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_287),
.A2(n_255),
.B(n_269),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_228),
.B(n_243),
.C(n_239),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_289),
.B(n_302),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_248),
.B(n_233),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_305),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_248),
.A2(n_233),
.B1(n_235),
.B2(n_229),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_265),
.A2(n_272),
.B(n_279),
.C(n_263),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_268),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_235),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_309),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_251),
.B(n_225),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_273),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_311),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_270),
.C(n_276),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_241),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_315),
.A2(n_238),
.B1(n_250),
.B2(n_255),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_316),
.B(n_330),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_273),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_319),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_257),
.Y(n_319)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_298),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_325),
.C(n_327),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_323),
.A2(n_346),
.B1(n_294),
.B2(n_312),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_254),
.C(n_246),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_326),
.A2(n_338),
.B(n_340),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_264),
.C(n_259),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_304),
.A2(n_252),
.B1(n_275),
.B2(n_218),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_328),
.A2(n_336),
.B1(n_305),
.B2(n_294),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_288),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_331),
.B(n_345),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_241),
.C(n_234),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_333),
.C(n_344),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_295),
.C(n_285),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_268),
.Y(n_334)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_286),
.A2(n_296),
.B1(n_291),
.B2(n_307),
.Y(n_335)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_296),
.A2(n_234),
.B1(n_211),
.B2(n_268),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_287),
.A2(n_211),
.B(n_164),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_298),
.A2(n_6),
.B(n_9),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_341),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_291),
.A2(n_125),
.B1(n_187),
.B2(n_14),
.Y(n_343)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_343),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_285),
.B(n_11),
.C(n_12),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_293),
.B(n_11),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_297),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_346)
);

OA22x2_ASAP7_75t_L g350 ( 
.A1(n_342),
.A2(n_309),
.B1(n_289),
.B2(n_303),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_350),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_351),
.A2(n_366),
.B1(n_367),
.B2(n_321),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_316),
.B(n_314),
.C(n_281),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_358),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_299),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_357),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_355),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_300),
.C(n_288),
.Y(n_358)
);

INVx13_ASAP7_75t_L g360 ( 
.A(n_318),
.Y(n_360)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_360),
.Y(n_378)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_324),
.Y(n_362)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_362),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_373),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_323),
.A2(n_312),
.B1(n_292),
.B2(n_299),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_368),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_333),
.B(n_306),
.Y(n_369)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_369),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_319),
.B(n_292),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_330),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_327),
.B(n_300),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_371),
.B(n_370),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_334),
.B(n_308),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_329),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_326),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_380),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_362),
.Y(n_377)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_357),
.B(n_329),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_385),
.C(n_395),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_361),
.Y(n_384)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_337),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_387),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_388),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_SL g389 ( 
.A(n_350),
.B(n_338),
.C(n_340),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_389),
.A2(n_363),
.B(n_350),
.Y(n_404)
);

FAx1_ASAP7_75t_SL g400 ( 
.A(n_390),
.B(n_364),
.CI(n_353),
.CON(n_400),
.SN(n_400)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_391),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_392),
.A2(n_348),
.B1(n_347),
.B2(n_372),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_344),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_393),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_308),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_394),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_322),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_332),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_352),
.C(n_358),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_399),
.A2(n_366),
.B1(n_385),
.B2(n_350),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_410),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_415),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_376),
.A2(n_348),
.B1(n_356),
.B2(n_290),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_402),
.A2(n_383),
.B1(n_378),
.B2(n_301),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

BUFx12_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_404),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_379),
.A2(n_346),
.B1(n_336),
.B2(n_352),
.Y(n_413)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_413),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_397),
.A2(n_363),
.B(n_386),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_417),
.B(n_380),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_406),
.A2(n_397),
.B(n_392),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_418),
.B(n_411),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_421),
.B(n_423),
.Y(n_436)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_422),
.Y(n_434)
);

BUFx24_ASAP7_75t_SL g423 ( 
.A(n_409),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_430),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_395),
.C(n_398),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_425),
.B(n_432),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_412),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_431),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_429),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_408),
.A2(n_375),
.B1(n_396),
.B2(n_371),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_415),
.A2(n_390),
.B1(n_364),
.B2(n_301),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_403),
.C(n_409),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_433),
.B(n_444),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_417),
.Y(n_435)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_435),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_416),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_407),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_445),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_SL g440 ( 
.A(n_427),
.B(n_400),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_440),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_400),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_403),
.C(n_411),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_381),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_428),
.C(n_418),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_453),
.Y(n_461)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_405),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_414),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_360),
.Y(n_463)
);

AOI21x1_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_421),
.B(n_414),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_456),
.A2(n_458),
.B(n_434),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_457),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_443),
.A2(n_408),
.B(n_401),
.Y(n_458)
);

NOR2x1_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_443),
.Y(n_459)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_459),
.Y(n_468)
);

AOI21xp33_ASAP7_75t_L g460 ( 
.A1(n_451),
.A2(n_442),
.B(n_436),
.Y(n_460)
);

A2O1A1Ixp33_ASAP7_75t_SL g469 ( 
.A1(n_460),
.A2(n_447),
.B(n_455),
.C(n_449),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_450),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_463),
.B(n_466),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_448),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_459),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_469),
.A2(n_471),
.B(n_455),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_465),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_470),
.B(n_464),
.C(n_447),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_472),
.B(n_473),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_474),
.B(n_468),
.C(n_469),
.Y(n_476)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_476),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_477),
.A2(n_475),
.B(n_311),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_12),
.Y(n_479)
);


endmodule