module real_aes_1349_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_0), .B(n_503), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_1), .A2(n_505), .B(n_506), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_2), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_3), .B(n_181), .Y(n_539) );
INVx1_ASAP7_75t_L g136 ( .A(n_4), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_5), .B(n_145), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_6), .B(n_181), .Y(n_527) );
INVx1_ASAP7_75t_L g191 ( .A(n_7), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_8), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_9), .Y(n_207) );
NAND2xp33_ASAP7_75t_L g560 ( .A(n_10), .B(n_178), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_11), .A2(n_493), .B1(n_820), .B2(n_821), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_11), .Y(n_820) );
INVx2_ASAP7_75t_L g144 ( .A(n_12), .Y(n_144) );
AOI221x1_ASAP7_75t_L g584 ( .A1(n_13), .A2(n_27), .B1(n_503), .B2(n_505), .C(n_585), .Y(n_584) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_14), .B(n_108), .C(n_110), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_14), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_15), .B(n_503), .Y(n_556) );
INVx1_ASAP7_75t_L g179 ( .A(n_16), .Y(n_179) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_17), .A2(n_167), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_18), .B(n_221), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_19), .A2(n_100), .B1(n_111), .B2(n_822), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_20), .B(n_181), .Y(n_516) );
AO21x1_ASAP7_75t_L g534 ( .A1(n_21), .A2(n_503), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g105 ( .A(n_22), .Y(n_105) );
AOI221xp5_ASAP7_75t_L g113 ( .A1(n_23), .A2(n_114), .B1(n_794), .B2(n_795), .C(n_799), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g794 ( .A(n_23), .Y(n_794) );
INVx1_ASAP7_75t_L g176 ( .A(n_24), .Y(n_176) );
INVx1_ASAP7_75t_SL g251 ( .A(n_25), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_26), .B(n_156), .Y(n_155) );
AOI33xp33_ASAP7_75t_L g228 ( .A1(n_28), .A2(n_55), .A3(n_133), .B1(n_151), .B2(n_229), .B3(n_230), .Y(n_228) );
NAND2x1_ASAP7_75t_L g577 ( .A(n_29), .B(n_181), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_30), .Y(n_800) );
NAND2x1_ASAP7_75t_L g526 ( .A(n_31), .B(n_178), .Y(n_526) );
INVx1_ASAP7_75t_L g200 ( .A(n_32), .Y(n_200) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_33), .A2(n_86), .B(n_144), .Y(n_143) );
OR2x2_ASAP7_75t_L g146 ( .A(n_33), .B(n_86), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_34), .B(n_189), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_35), .B(n_178), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_36), .B(n_181), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_37), .B(n_178), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_38), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_39), .A2(n_505), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g139 ( .A(n_40), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g150 ( .A(n_40), .Y(n_150) );
AND2x2_ASAP7_75t_L g165 ( .A(n_40), .B(n_136), .Y(n_165) );
INVxp67_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
OR2x6_ASAP7_75t_L g120 ( .A(n_41), .B(n_104), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_42), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_43), .B(n_503), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_44), .B(n_189), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_45), .A2(n_130), .B1(n_142), .B2(n_145), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_46), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_47), .B(n_156), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_48), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_49), .B(n_178), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_50), .B(n_167), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_51), .B(n_156), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_52), .A2(n_505), .B(n_525), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_53), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_54), .B(n_178), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_56), .B(n_156), .Y(n_219) );
INVx1_ASAP7_75t_L g134 ( .A(n_57), .Y(n_134) );
INVx1_ASAP7_75t_L g158 ( .A(n_57), .Y(n_158) );
AND2x2_ASAP7_75t_L g220 ( .A(n_58), .B(n_221), .Y(n_220) );
AOI221xp5_ASAP7_75t_L g188 ( .A1(n_59), .A2(n_75), .B1(n_148), .B2(n_189), .C(n_190), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_60), .B(n_189), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_61), .B(n_181), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_62), .B(n_142), .Y(n_209) );
AOI21xp5_ASAP7_75t_SL g239 ( .A1(n_63), .A2(n_148), .B(n_240), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_64), .A2(n_505), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g172 ( .A(n_65), .Y(n_172) );
AO21x1_ASAP7_75t_L g536 ( .A1(n_66), .A2(n_505), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_67), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g218 ( .A(n_68), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_69), .B(n_503), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_70), .A2(n_148), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g550 ( .A(n_71), .B(n_222), .Y(n_550) );
INVx1_ASAP7_75t_L g140 ( .A(n_72), .Y(n_140) );
INVx1_ASAP7_75t_L g160 ( .A(n_72), .Y(n_160) );
AND2x2_ASAP7_75t_L g529 ( .A(n_73), .B(n_196), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_74), .B(n_189), .Y(n_231) );
AND2x2_ASAP7_75t_L g253 ( .A(n_76), .B(n_196), .Y(n_253) );
INVx1_ASAP7_75t_L g173 ( .A(n_77), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_78), .A2(n_148), .B(n_250), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_79), .A2(n_148), .B(n_154), .C(n_166), .Y(n_147) );
INVx1_ASAP7_75t_L g106 ( .A(n_80), .Y(n_106) );
AND2x2_ASAP7_75t_L g500 ( .A(n_81), .B(n_196), .Y(n_500) );
AND2x2_ASAP7_75t_SL g237 ( .A(n_82), .B(n_196), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_83), .B(n_503), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_84), .A2(n_148), .B1(n_226), .B2(n_227), .Y(n_225) );
AND2x2_ASAP7_75t_L g535 ( .A(n_85), .B(n_145), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_87), .B(n_178), .Y(n_517) );
AND2x2_ASAP7_75t_L g580 ( .A(n_88), .B(n_196), .Y(n_580) );
INVx1_ASAP7_75t_L g241 ( .A(n_89), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_90), .B(n_181), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_91), .A2(n_505), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_92), .B(n_178), .Y(n_586) );
AND2x2_ASAP7_75t_L g232 ( .A(n_93), .B(n_196), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_94), .B(n_181), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_95), .A2(n_198), .B(n_199), .C(n_201), .Y(n_197) );
BUFx2_ASAP7_75t_SL g816 ( .A(n_96), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_97), .A2(n_505), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_98), .B(n_156), .Y(n_242) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_SL g825 ( .A(n_102), .Y(n_825) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_107), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_812), .B(n_817), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g112 ( .A(n_113), .B(n_804), .Y(n_112) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_121), .B1(n_493), .B2(n_792), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_116), .A2(n_121), .B1(n_493), .B2(n_797), .Y(n_796) );
CKINVDCx11_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
OR2x6_ASAP7_75t_SL g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AND2x6_ASAP7_75t_SL g793 ( .A(n_118), .B(n_120), .Y(n_793) );
OR2x2_ASAP7_75t_L g803 ( .A(n_118), .B(n_120), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_118), .B(n_119), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_427), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_350), .Y(n_122) );
NAND3xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_297), .C(n_330), .Y(n_123) );
AOI211xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_254), .B(n_263), .C(n_287), .Y(n_124) );
OAI21xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_183), .B(n_233), .Y(n_125) );
OR2x2_ASAP7_75t_L g307 ( .A(n_126), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g462 ( .A(n_126), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_127), .A2(n_353), .B1(n_357), .B2(n_359), .Y(n_352) );
AND2x2_ASAP7_75t_L g389 ( .A(n_127), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_168), .Y(n_127) );
INVx1_ASAP7_75t_L g286 ( .A(n_128), .Y(n_286) );
AND2x4_ASAP7_75t_L g303 ( .A(n_128), .B(n_284), .Y(n_303) );
INVx2_ASAP7_75t_L g325 ( .A(n_128), .Y(n_325) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_128), .Y(n_408) );
AND2x2_ASAP7_75t_L g479 ( .A(n_128), .B(n_236), .Y(n_479) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_147), .Y(n_128) );
NOR3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_137), .C(n_141), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g189 ( .A(n_132), .B(n_138), .Y(n_189) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
OR2x6_ASAP7_75t_L g163 ( .A(n_133), .B(n_152), .Y(n_163) );
INVxp33_ASAP7_75t_L g229 ( .A(n_133), .Y(n_229) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g153 ( .A(n_134), .B(n_136), .Y(n_153) );
AND2x4_ASAP7_75t_L g181 ( .A(n_134), .B(n_159), .Y(n_181) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x6_ASAP7_75t_L g505 ( .A(n_139), .B(n_153), .Y(n_505) );
INVx2_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
AND2x6_ASAP7_75t_L g178 ( .A(n_140), .B(n_157), .Y(n_178) );
INVx4_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_142), .B(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx4f_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
AND2x4_ASAP7_75t_L g145 ( .A(n_144), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_144), .B(n_146), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_145), .B(n_164), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_145), .A2(n_239), .B(n_243), .Y(n_238) );
INVx1_ASAP7_75t_SL g512 ( .A(n_145), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_145), .B(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_145), .A2(n_556), .B(n_557), .Y(n_555) );
INVxp67_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NOR2x1p5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx1_ASAP7_75t_L g230 ( .A(n_151), .Y(n_230) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_161), .B(n_164), .Y(n_154) );
INVx1_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
AND2x4_ASAP7_75t_L g503 ( .A(n_156), .B(n_165), .Y(n_503) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_163), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_163), .A2(n_164), .B(n_191), .C(n_192), .Y(n_190) );
INVxp67_ASAP7_75t_L g198 ( .A(n_163), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_163), .A2(n_164), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_163), .A2(n_164), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g250 ( .A1(n_163), .A2(n_164), .B(n_251), .C(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g226 ( .A(n_164), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_164), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_164), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_164), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_164), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_164), .A2(n_547), .B(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_164), .A2(n_559), .B(n_560), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_164), .A2(n_577), .B(n_578), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_164), .A2(n_586), .B(n_587), .Y(n_585) );
INVx5_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_166), .A2(n_224), .B(n_232), .Y(n_223) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_166), .A2(n_224), .B(n_232), .Y(n_268) );
INVx2_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_167), .A2(n_188), .B(n_193), .Y(n_187) );
AND2x2_ASAP7_75t_L g244 ( .A(n_168), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g273 ( .A(n_168), .Y(n_273) );
INVx3_ASAP7_75t_L g284 ( .A(n_168), .Y(n_284) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_175), .B(n_182), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_174), .B(n_200), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B1(n_179), .B2(n_180), .Y(n_175) );
INVxp67_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVxp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_183), .A2(n_474), .B1(n_476), .B2(n_478), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_183), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_211), .Y(n_184) );
INVx3_ASAP7_75t_L g257 ( .A(n_185), .Y(n_257) );
AND2x2_ASAP7_75t_L g265 ( .A(n_185), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_185), .Y(n_295) );
NAND2x1_ASAP7_75t_SL g489 ( .A(n_185), .B(n_256), .Y(n_489) );
AND2x4_ASAP7_75t_L g185 ( .A(n_186), .B(n_194), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g262 ( .A(n_187), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_187), .B(n_268), .Y(n_280) );
AND2x2_ASAP7_75t_L g293 ( .A(n_187), .B(n_194), .Y(n_293) );
AND2x4_ASAP7_75t_L g300 ( .A(n_187), .B(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_187), .Y(n_349) );
INVxp67_ASAP7_75t_L g356 ( .A(n_187), .Y(n_356) );
INVx1_ASAP7_75t_L g361 ( .A(n_187), .Y(n_361) );
INVx1_ASAP7_75t_L g210 ( .A(n_189), .Y(n_210) );
INVx1_ASAP7_75t_L g260 ( .A(n_194), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_194), .B(n_270), .Y(n_279) );
INVx2_ASAP7_75t_L g347 ( .A(n_194), .Y(n_347) );
INVx1_ASAP7_75t_L g386 ( .A(n_194), .Y(n_386) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_204), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B1(n_202), .B2(n_203), .Y(n_195) );
INVx3_ASAP7_75t_L g203 ( .A(n_196), .Y(n_203) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_203), .A2(n_214), .B(n_220), .Y(n_213) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_203), .A2(n_214), .B(n_220), .Y(n_270) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_203), .A2(n_544), .B(n_550), .Y(n_543) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_203), .A2(n_544), .B(n_550), .Y(n_565) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_203), .A2(n_574), .B(n_580), .Y(n_573) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_203), .A2(n_574), .B(n_580), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_208), .B1(n_209), .B2(n_210), .Y(n_204) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g316 ( .A(n_211), .B(n_293), .Y(n_316) );
AND2x2_ASAP7_75t_L g384 ( .A(n_211), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g398 ( .A(n_211), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_211), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_223), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_213), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g354 ( .A(n_213), .B(n_347), .Y(n_354) );
AND2x2_ASAP7_75t_L g445 ( .A(n_213), .B(n_267), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_221), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_221), .A2(n_502), .B(n_504), .Y(n_501) );
OA21x2_ASAP7_75t_L g583 ( .A1(n_221), .A2(n_584), .B(n_588), .Y(n_583) );
OA21x2_ASAP7_75t_L g628 ( .A1(n_221), .A2(n_584), .B(n_588), .Y(n_628) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
INVx2_ASAP7_75t_L g301 ( .A(n_223), .Y(n_301) );
AND2x2_ASAP7_75t_L g346 ( .A(n_223), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_225), .B(n_231), .Y(n_224) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_244), .Y(n_234) );
AND2x2_ASAP7_75t_L g388 ( .A(n_235), .B(n_389), .Y(n_388) );
OR2x6_ASAP7_75t_L g447 ( .A(n_235), .B(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx4_ASAP7_75t_L g277 ( .A(n_236), .Y(n_277) );
AND2x4_ASAP7_75t_L g285 ( .A(n_236), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g320 ( .A(n_236), .B(n_245), .Y(n_320) );
INVx2_ASAP7_75t_L g369 ( .A(n_236), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_236), .B(n_343), .Y(n_418) );
AND2x2_ASAP7_75t_L g455 ( .A(n_236), .B(n_273), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_236), .B(n_338), .Y(n_463) );
OR2x6_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_L g296 ( .A(n_244), .B(n_285), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_244), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_244), .B(n_323), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_244), .B(n_336), .Y(n_457) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_245), .Y(n_275) );
AND2x2_ASAP7_75t_L g283 ( .A(n_245), .B(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_245), .Y(n_306) );
INVx2_ASAP7_75t_L g309 ( .A(n_245), .Y(n_309) );
INVx1_ASAP7_75t_L g342 ( .A(n_245), .Y(n_342) );
INVx1_ASAP7_75t_L g390 ( .A(n_245), .Y(n_390) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_253), .Y(n_245) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_246), .A2(n_523), .B(n_529), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
NAND2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_256), .B(n_259), .Y(n_332) );
OR2x2_ASAP7_75t_L g404 ( .A(n_256), .B(n_405), .Y(n_404) );
AND4x1_ASAP7_75t_SL g450 ( .A(n_256), .B(n_432), .C(n_451), .D(n_452), .Y(n_450) );
OR2x2_ASAP7_75t_L g474 ( .A(n_257), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g311 ( .A(n_260), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_260), .B(n_269), .Y(n_461) );
AND2x2_ASAP7_75t_L g486 ( .A(n_261), .B(n_346), .Y(n_486) );
OAI32xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_271), .A3(n_276), .B1(n_278), .B2(n_281), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g359 ( .A(n_266), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g459 ( .A(n_266), .B(n_413), .Y(n_459) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
AND2x2_ASAP7_75t_L g355 ( .A(n_267), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g441 ( .A(n_267), .Y(n_441) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_268), .B(n_270), .Y(n_475) );
INVx3_ASAP7_75t_L g292 ( .A(n_269), .Y(n_292) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_269), .B(n_397), .Y(n_470) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_270), .Y(n_329) );
AND2x2_ASAP7_75t_L g348 ( .A(n_270), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g482 ( .A(n_272), .Y(n_482) );
NAND2x1_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g322 ( .A(n_273), .Y(n_322) );
NOR2x1_ASAP7_75t_L g423 ( .A(n_273), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_276), .B(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g314 ( .A(n_277), .B(n_282), .Y(n_314) );
AND2x4_ASAP7_75t_L g336 ( .A(n_277), .B(n_286), .Y(n_336) );
AND2x4_ASAP7_75t_SL g407 ( .A(n_277), .B(n_408), .Y(n_407) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_277), .B(n_358), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_278), .A2(n_401), .B1(n_404), .B2(n_406), .Y(n_400) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_SL g420 ( .A(n_279), .Y(n_420) );
INVx2_ASAP7_75t_L g312 ( .A(n_280), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_283), .B(n_289), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_283), .A2(n_419), .B1(n_422), .B2(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g343 ( .A(n_284), .Y(n_343) );
AND2x2_ASAP7_75t_L g366 ( .A(n_284), .B(n_325), .Y(n_366) );
INVx2_ASAP7_75t_L g289 ( .A(n_285), .Y(n_289) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_290), .B(n_294), .Y(n_287) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_291), .A2(n_363), .B1(n_367), .B2(n_368), .Y(n_362) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_292), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_292), .B(n_360), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_292), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NOR3xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_313), .C(n_317), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B1(n_307), .B2(n_310), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g327 ( .A(n_300), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g367 ( .A(n_300), .B(n_354), .Y(n_367) );
AND2x2_ASAP7_75t_L g419 ( .A(n_300), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g436 ( .A(n_300), .B(n_386), .Y(n_436) );
AND2x2_ASAP7_75t_L g491 ( .A(n_300), .B(n_385), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx4_ASAP7_75t_L g358 ( .A(n_303), .Y(n_358) );
AND2x2_ASAP7_75t_L g368 ( .A(n_303), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g373 ( .A(n_306), .Y(n_373) );
AND2x2_ASAP7_75t_L g382 ( .A(n_306), .B(n_366), .Y(n_382) );
INVx1_ASAP7_75t_L g417 ( .A(n_308), .Y(n_417) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g338 ( .A(n_309), .Y(n_338) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_311), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_312), .B(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_326), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_319), .B(n_358), .Y(n_467) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AOI21xp33_ASAP7_75t_SL g330 ( .A1(n_322), .A2(n_331), .B(n_333), .Y(n_330) );
AND2x2_ASAP7_75t_L g477 ( .A(n_322), .B(n_336), .Y(n_477) );
AND2x4_ASAP7_75t_L g340 ( .A(n_323), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g374 ( .A(n_323), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_323), .B(n_390), .Y(n_456) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI21xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_339), .B(n_344), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_336), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_336), .B(n_341), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_337), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g399 ( .A(n_337), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_337), .Y(n_403) );
AND2x2_ASAP7_75t_L g487 ( .A(n_337), .B(n_455), .Y(n_487) );
AND2x2_ASAP7_75t_L g490 ( .A(n_337), .B(n_407), .Y(n_490) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_342), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g469 ( .A(n_346), .Y(n_469) );
AND2x2_ASAP7_75t_L g360 ( .A(n_347), .B(n_361), .Y(n_360) );
NAND4xp75_ASAP7_75t_L g350 ( .A(n_351), .B(n_370), .C(n_391), .D(n_409), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_362), .Y(n_351) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_354), .B(n_441), .Y(n_440) );
NAND2x1p5_ASAP7_75t_L g426 ( .A(n_355), .B(n_420), .Y(n_426) );
NAND2xp5_ASAP7_75t_R g442 ( .A(n_358), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g492 ( .A(n_358), .Y(n_492) );
INVx2_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
BUFx3_ASAP7_75t_L g397 ( .A(n_361), .Y(n_397) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g448 ( .A(n_366), .Y(n_448) );
AND2x2_ASAP7_75t_L g402 ( .A(n_368), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g424 ( .A(n_369), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .B(n_377), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_373), .B(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_374), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_376), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_381), .B1(n_383), .B2(n_387), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_385), .A2(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g413 ( .A(n_385), .Y(n_413) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g444 ( .A(n_386), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g452 ( .A(n_386), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_387), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g422 ( .A(n_390), .B(n_423), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_398), .B(n_400), .Y(n_391) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g439 ( .A(n_396), .B(n_440), .Y(n_439) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
INVx2_ASAP7_75t_SL g443 ( .A(n_407), .Y(n_443) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_421), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_414), .B1(n_416), .B2(n_419), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g472 ( .A(n_416), .Y(n_472) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_464), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_437), .C(n_449), .Y(n_428) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_434), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_442), .B1(n_444), .B2(n_446), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .C(n_460), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .B(n_458), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_483), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_473), .C(n_480), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_471), .B2(n_472), .Y(n_466) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_474), .B(n_479), .C(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI222xp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_487), .B1(n_488), .B2(n_490), .C1(n_491), .C2(n_492), .Y(n_483) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g821 ( .A(n_493), .Y(n_821) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_677), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_632), .C(n_661), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_496), .B(n_605), .Y(n_495) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_530), .B1(n_551), .B2(n_562), .C(n_566), .Y(n_496) );
INVx3_ASAP7_75t_SL g722 ( .A(n_497), .Y(n_722) );
AND2x2_ASAP7_75t_SL g497 ( .A(n_498), .B(n_509), .Y(n_497) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_498), .B(n_521), .Y(n_568) );
INVx4_ASAP7_75t_L g603 ( .A(n_498), .Y(n_603) );
AND2x2_ASAP7_75t_L g625 ( .A(n_498), .B(n_522), .Y(n_625) );
AND2x2_ASAP7_75t_L g631 ( .A(n_498), .B(n_570), .Y(n_631) );
INVx5_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g600 ( .A(n_499), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_499), .B(n_521), .Y(n_676) );
AND2x2_ASAP7_75t_L g681 ( .A(n_499), .B(n_522), .Y(n_681) );
AND2x2_ASAP7_75t_L g693 ( .A(n_499), .B(n_554), .Y(n_693) );
NOR2x1_ASAP7_75t_SL g732 ( .A(n_499), .B(n_570), .Y(n_732) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g561 ( .A(n_509), .Y(n_561) );
AND2x2_ASAP7_75t_L g665 ( .A(n_509), .B(n_614), .Y(n_665) );
AND2x2_ASAP7_75t_L g762 ( .A(n_509), .B(n_693), .Y(n_762) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g594 ( .A(n_511), .Y(n_594) );
INVx2_ASAP7_75t_L g616 ( .A(n_511), .Y(n_616) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_512), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .Y(n_513) );
AND2x2_ASAP7_75t_L g591 ( .A(n_521), .B(n_553), .Y(n_591) );
INVx2_ASAP7_75t_L g595 ( .A(n_521), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_521), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g694 ( .A(n_521), .B(n_659), .Y(n_694) );
OR2x2_ASAP7_75t_L g741 ( .A(n_521), .B(n_554), .Y(n_741) );
INVx4_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_522), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_528), .Y(n_523) );
AND2x2_ASAP7_75t_L g738 ( .A(n_530), .B(n_619), .Y(n_738) );
AND2x2_ASAP7_75t_L g788 ( .A(n_530), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g664 ( .A(n_531), .B(n_608), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_542), .Y(n_531) );
AND2x2_ASAP7_75t_L g597 ( .A(n_532), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g627 ( .A(n_532), .B(n_628), .Y(n_627) );
AND2x4_ASAP7_75t_L g648 ( .A(n_532), .B(n_628), .Y(n_648) );
AND2x4_ASAP7_75t_L g683 ( .A(n_532), .B(n_671), .Y(n_683) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g564 ( .A(n_533), .Y(n_564) );
OAI21x1_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_536), .B(n_540), .Y(n_533) );
INVx1_ASAP7_75t_L g541 ( .A(n_535), .Y(n_541) );
AND2x2_ASAP7_75t_L g610 ( .A(n_542), .B(n_563), .Y(n_610) );
AND2x2_ASAP7_75t_L g696 ( .A(n_542), .B(n_628), .Y(n_696) );
AND2x2_ASAP7_75t_L g707 ( .A(n_542), .B(n_572), .Y(n_707) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g571 ( .A(n_543), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g638 ( .A(n_543), .B(n_573), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_545), .B(n_549), .Y(n_544) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_561), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_553), .B(n_603), .Y(n_660) );
AND2x2_ASAP7_75t_L g704 ( .A(n_553), .B(n_570), .Y(n_704) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_554), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g614 ( .A(n_554), .Y(n_614) );
BUFx3_ASAP7_75t_L g623 ( .A(n_554), .Y(n_623) );
AND2x2_ASAP7_75t_L g646 ( .A(n_554), .B(n_616), .Y(n_646) );
OAI322xp33_ASAP7_75t_L g566 ( .A1(n_561), .A2(n_567), .A3(n_571), .B1(n_581), .B2(n_589), .C1(n_596), .C2(n_601), .Y(n_566) );
INVx1_ASAP7_75t_L g727 ( .A(n_561), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_562), .B(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_L g640 ( .A(n_562), .B(n_582), .Y(n_640) );
INVx2_ASAP7_75t_L g685 ( .A(n_562), .Y(n_685) );
AND2x2_ASAP7_75t_L g701 ( .A(n_562), .B(n_643), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_562), .B(n_719), .Y(n_749) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_563), .B(n_628), .Y(n_652) );
OR2x2_ASAP7_75t_L g673 ( .A(n_563), .B(n_590), .Y(n_673) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g645 ( .A(n_564), .Y(n_645) );
INVx2_ASAP7_75t_L g590 ( .A(n_565), .Y(n_590) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_565), .Y(n_592) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx2_ASAP7_75t_L g635 ( .A(n_568), .Y(n_635) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_569), .Y(n_655) );
INVx1_ASAP7_75t_L g753 ( .A(n_569), .Y(n_753) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_569), .Y(n_768) );
NAND2x1_ASAP7_75t_L g778 ( .A(n_571), .B(n_582), .Y(n_778) );
INVx1_ASAP7_75t_L g785 ( .A(n_571), .Y(n_785) );
BUFx2_ASAP7_75t_L g619 ( .A(n_572), .Y(n_619) );
AND2x2_ASAP7_75t_L g695 ( .A(n_572), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx3_ASAP7_75t_L g604 ( .A(n_573), .Y(n_604) );
INVxp67_ASAP7_75t_L g608 ( .A(n_573), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_579), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_581), .B(n_597), .C(n_599), .Y(n_596) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_SL g617 ( .A(n_582), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_582), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g769 ( .A(n_582), .B(n_718), .Y(n_769) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g671 ( .A(n_583), .Y(n_671) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_583), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_592), .B2(n_593), .Y(n_589) );
AND2x4_ASAP7_75t_SL g718 ( .A(n_590), .B(n_598), .Y(n_718) );
AND2x2_ASAP7_75t_L g731 ( .A(n_591), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_592), .Y(n_733) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx2_ASAP7_75t_L g690 ( .A(n_594), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_594), .B(n_603), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_595), .B(n_613), .Y(n_612) );
AND3x2_ASAP7_75t_L g630 ( .A(n_595), .B(n_623), .C(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g654 ( .A(n_595), .Y(n_654) );
AND2x2_ASAP7_75t_L g767 ( .A(n_595), .B(n_768), .Y(n_767) );
BUFx2_ASAP7_75t_L g643 ( .A(n_598), .Y(n_643) );
INVx1_ASAP7_75t_L g721 ( .A(n_598), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_599), .B(n_622), .Y(n_760) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_600), .B(n_704), .Y(n_709) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AND2x2_ASAP7_75t_L g700 ( .A(n_603), .B(n_646), .Y(n_700) );
INVx1_ASAP7_75t_SL g651 ( .A(n_604), .Y(n_651) );
AND2x2_ASAP7_75t_L g759 ( .A(n_604), .B(n_671), .Y(n_759) );
AND2x2_ASAP7_75t_L g780 ( .A(n_604), .B(n_652), .Y(n_780) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_611), .B1(n_617), .B2(n_620), .C(n_626), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g772 ( .A(n_608), .Y(n_772) );
AOI21xp33_ASAP7_75t_SL g626 ( .A1(n_609), .A2(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g618 ( .A(n_610), .B(n_619), .Y(n_618) );
AOI222xp33_ASAP7_75t_L g641 ( .A1(n_610), .A2(n_642), .B1(n_644), .B2(n_649), .C1(n_653), .C2(n_656), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_610), .B(n_759), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_611), .A2(n_640), .B1(n_663), .B2(n_665), .Y(n_662) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g647 ( .A(n_614), .Y(n_647) );
AND2x2_ASAP7_75t_L g766 ( .A(n_614), .B(n_732), .Y(n_766) );
OAI32xp33_ASAP7_75t_L g770 ( .A1(n_614), .A2(n_639), .A3(n_691), .B1(n_699), .B2(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g775 ( .A(n_614), .B(n_625), .Y(n_775) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g659 ( .A(n_616), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_617), .A2(n_667), .B(n_674), .Y(n_666) );
INVx1_ASAP7_75t_L g730 ( .A(n_619), .Y(n_730) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g634 ( .A(n_622), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g642 ( .A(n_625), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g715 ( .A(n_625), .B(n_646), .Y(n_715) );
INVx1_ASAP7_75t_SL g786 ( .A(n_627), .Y(n_786) );
AND2x2_ASAP7_75t_L g720 ( .A(n_628), .B(n_721), .Y(n_720) );
OAI222xp33_ASAP7_75t_L g773 ( .A1(n_629), .A2(n_682), .B1(n_761), .B2(n_774), .C1(n_776), .C2(n_778), .Y(n_773) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g746 ( .A(n_631), .B(n_747), .Y(n_746) );
OAI21xp33_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_636), .B(n_641), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_635), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g714 ( .A(n_637), .Y(n_714) );
INVx1_ASAP7_75t_L g682 ( .A(n_638), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_638), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g736 ( .A(n_643), .Y(n_736) );
AO22x1_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_644) );
OAI322xp33_ASAP7_75t_L g756 ( .A1(n_645), .A2(n_706), .A3(n_709), .B1(n_757), .B2(n_758), .C1(n_760), .C2(n_761), .Y(n_756) );
AND2x2_ASAP7_75t_SL g680 ( .A(n_646), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g675 ( .A(n_647), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_648), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g777 ( .A(n_648), .B(n_707), .Y(n_777) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g757 ( .A(n_651), .Y(n_757) );
INVx1_ASAP7_75t_SL g686 ( .A(n_652), .Y(n_686) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
OR2x2_ASAP7_75t_L g688 ( .A(n_660), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g726 ( .A(n_660), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_666), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_672), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g699 ( .A(n_670), .B(n_685), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_670), .B(n_707), .Y(n_706) );
BUFx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g729 ( .A(n_673), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NOR2x1_ASAP7_75t_L g677 ( .A(n_678), .B(n_742), .Y(n_677) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_697), .C(n_710), .D(n_723), .Y(n_678) );
AOI322xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_682), .A3(n_683), .B1(n_684), .B2(n_687), .C1(n_692), .C2(n_695), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g779 ( .A1(n_680), .A2(n_780), .B(n_781), .C(n_784), .Y(n_779) );
AND2x2_ASAP7_75t_L g791 ( .A(n_681), .B(n_768), .Y(n_791) );
INVx1_ASAP7_75t_L g713 ( .A(n_683), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_683), .B(n_718), .Y(n_755) );
NAND2xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_691), .B(n_704), .Y(n_771) );
AND2x4_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B1(n_701), .B2(n_702), .C1(n_705), .C2(n_708), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_700), .A2(n_711), .B1(n_714), .B2(n_715), .C(n_716), .Y(n_710) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI21xp33_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_719), .B(n_722), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_728), .B1(n_731), .B2(n_733), .C(n_734), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g783 ( .A(n_732), .Y(n_783) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B(n_739), .Y(n_734) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx2_ASAP7_75t_L g747 ( .A(n_741), .Y(n_747) );
OR2x2_ASAP7_75t_L g782 ( .A(n_741), .B(n_783), .Y(n_782) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_763), .C(n_779), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_756), .Y(n_743) );
OAI21xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B(n_750), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_754), .Y(n_750) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_769), .B1(n_770), .B2(n_772), .C(n_773), .Y(n_763) );
INVxp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NOR2x1_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_778), .B(n_782), .Y(n_781) );
O2A1O1Ixp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .B(n_787), .C(n_790), .Y(n_784) );
INVxp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
CKINVDCx11_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_793), .Y(n_798) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx3_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
INVx2_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
INVx3_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVxp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_805), .A2(n_810), .B(n_819), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
BUFx3_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_SL g812 ( .A(n_813), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_814), .B(n_818), .Y(n_817) );
CKINVDCx11_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
CKINVDCx8_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx3_ASAP7_75t_SL g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
endmodule