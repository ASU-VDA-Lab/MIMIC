module fake_jpeg_16111_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx11_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_7),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_29),
.B1(n_25),
.B2(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_51),
.B1(n_58),
.B2(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_28),
.B1(n_29),
.B2(n_19),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_50),
.B1(n_59),
.B2(n_38),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_31),
.B1(n_20),
.B2(n_19),
.Y(n_46)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_32),
.B1(n_27),
.B2(n_2),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_43),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_29),
.B1(n_24),
.B2(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_22),
.B1(n_26),
.B2(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_22),
.B1(n_26),
.B2(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_23),
.B1(n_31),
.B2(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_20),
.B1(n_23),
.B2(n_32),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_50),
.B1(n_46),
.B2(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_30),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_76),
.B1(n_55),
.B2(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_62),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_47),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_30),
.B1(n_32),
.B2(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_30),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_86),
.B(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_27),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_66),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_99),
.Y(n_118)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_109),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_63),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_100),
.C(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_81),
.B1(n_77),
.B2(n_68),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_49),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_64),
.C(n_48),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_46),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_108),
.B(n_111),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_66),
.C(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_57),
.Y(n_123)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_78),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_76),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_77),
.B1(n_83),
.B2(n_67),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_81),
.B(n_85),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_123),
.B(n_108),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_69),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_111),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_67),
.B(n_83),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_93),
.B(n_104),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_79),
.B1(n_87),
.B2(n_88),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_79),
.B1(n_65),
.B2(n_57),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_130),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_75),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_0),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_3),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_65),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_136),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_143),
.B(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_90),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_100),
.B(n_112),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_110),
.B1(n_105),
.B2(n_98),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_155),
.B1(n_114),
.B2(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_154),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_153),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_152),
.C(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_109),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_98),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_92),
.A3(n_102),
.B1(n_56),
.B2(n_57),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_156),
.B(n_131),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_164),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_160),
.B(n_169),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_177),
.B1(n_139),
.B2(n_143),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_132),
.C(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_130),
.C(n_129),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_170),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_137),
.C(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_119),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_146),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_157),
.B1(n_139),
.B2(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_184),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_144),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_167),
.Y(n_199)
);

INVxp33_ASAP7_75t_SL g186 ( 
.A(n_163),
.Y(n_186)
);

AO221x1_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_160),
.B1(n_178),
.B2(n_169),
.C(n_177),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_127),
.B1(n_145),
.B2(n_142),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_149),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_194),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_119),
.B1(n_115),
.B2(n_127),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_127),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_170),
.CI(n_166),
.CON(n_196),
.SN(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_159),
.C(n_164),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_204),
.C(n_205),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_185),
.Y(n_213)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_206),
.B(n_190),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_168),
.C(n_176),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_176),
.C(n_161),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_127),
.B(n_173),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_192),
.B1(n_194),
.B2(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_197),
.B(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_216),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_4),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_209),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_174),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_202),
.B1(n_6),
.B2(n_8),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_173),
.B(n_155),
.C(n_113),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_206),
.B(n_201),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_56),
.C(n_5),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_4),
.C(n_6),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_224),
.A2(n_225),
.B(n_215),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_SL g225 ( 
.A(n_210),
.B(n_196),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_202),
.A3(n_203),
.B1(n_207),
.B2(n_196),
.C1(n_200),
.C2(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_227),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.C(n_217),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_4),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_224),
.A2(n_215),
.B(n_220),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_228),
.B(n_221),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_222),
.B(n_217),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_236),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_213),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_241),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_9),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_235),
.B1(n_230),
.B2(n_11),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

AO221x1_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_245),
.B1(n_10),
.B2(n_14),
.C(n_239),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_9),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_244),
.B(n_10),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_247),
.Y(n_250)
);


endmodule