module fake_jpeg_4765_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_1),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_2),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_49),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_26),
.B1(n_15),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_50),
.B1(n_16),
.B2(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_26),
.B1(n_15),
.B2(n_24),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_21),
.C(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_20),
.B1(n_15),
.B2(n_23),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_23),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_26),
.B1(n_15),
.B2(n_24),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_28),
.B1(n_23),
.B2(n_16),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_53),
.C(n_45),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_74),
.B1(n_75),
.B2(n_22),
.Y(n_80)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_73),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_28),
.C(n_5),
.Y(n_82)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_51),
.B1(n_59),
.B2(n_57),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_36),
.B1(n_32),
.B2(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_51),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_46),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_89),
.B(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_85),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_25),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_18),
.Y(n_107)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_93),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_78),
.B1(n_77),
.B2(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_58),
.B1(n_41),
.B2(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_94),
.B1(n_66),
.B2(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_41),
.B(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_25),
.Y(n_109)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_36),
.B1(n_43),
.B2(n_32),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_28),
.B(n_27),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_106),
.B(n_86),
.Y(n_123)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_109),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_79),
.C(n_77),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_111),
.C(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_65),
.C(n_63),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_92),
.B(n_87),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_123),
.B(n_18),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_120),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_88),
.B(n_86),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_27),
.B(n_18),
.Y(n_141)
);

INVxp33_ASAP7_75t_SL g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_130),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_125),
.C(n_37),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_80),
.C(n_94),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_84),
.B(n_90),
.C(n_33),
.D(n_31),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_27),
.B(n_18),
.C(n_35),
.D(n_31),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_109),
.A3(n_96),
.B1(n_97),
.B2(n_104),
.C1(n_107),
.C2(n_14),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_43),
.B1(n_55),
.B2(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_134),
.B(n_141),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_63),
.B(n_33),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_93),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_37),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_144),
.C(n_145),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_134),
.CI(n_132),
.CON(n_157),
.SN(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_146),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_37),
.C(n_35),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_124),
.B1(n_114),
.B2(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_117),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_150),
.C(n_27),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_124),
.C(n_120),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_124),
.B1(n_119),
.B2(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_160),
.B(n_27),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_3),
.C(n_5),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_55),
.Y(n_159)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_135),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_169),
.C(n_172),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_153),
.A2(n_140),
.B(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

AOI321xp33_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_35),
.A3(n_27),
.B1(n_55),
.B2(n_14),
.C(n_12),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_171),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_155),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_3),
.B(n_5),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_168),
.B(n_6),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_152),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_175),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_178),
.B(n_157),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_147),
.C(n_149),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_162),
.C(n_168),
.Y(n_184)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_180),
.B1(n_17),
.B2(n_8),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.C(n_7),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_157),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_171),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_183),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_186),
.B(n_12),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_194),
.B(n_9),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_7),
.C(n_9),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_197),
.B(n_198),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_182),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_10),
.A3(n_11),
.B1(n_17),
.B2(n_185),
.C1(n_191),
.C2(n_187),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_10),
.B(n_11),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_17),
.Y(n_202)
);


endmodule