module fake_jpeg_12132_n_469 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_45),
.Y(n_139)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_52),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_8),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_54),
.B(n_72),
.Y(n_137)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_35),
.A2(n_7),
.B(n_14),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_86),
.Y(n_96)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_88),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_18),
.B1(n_17),
.B2(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_93),
.B(n_109),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_38),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_94),
.B(n_97),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_30),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_98),
.A2(n_80),
.B1(n_75),
.B2(n_57),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_102),
.A2(n_104),
.B1(n_129),
.B2(n_51),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_17),
.B1(n_23),
.B2(n_27),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_41),
.B1(n_40),
.B2(n_34),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_105),
.A2(n_142),
.B1(n_102),
.B2(n_104),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_30),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_45),
.B(n_41),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_139),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_17),
.B1(n_27),
.B2(n_42),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_47),
.B(n_34),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_138),
.B(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_49),
.B(n_34),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_53),
.A2(n_29),
.B1(n_40),
.B2(n_33),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_61),
.B(n_41),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_33),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_174),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_149),
.A2(n_162),
.B1(n_170),
.B2(n_183),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_29),
.B1(n_87),
.B2(n_86),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_151),
.A2(n_156),
.B1(n_166),
.B2(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_154),
.A2(n_98),
.B1(n_27),
.B2(n_129),
.Y(n_205)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_88),
.B1(n_68),
.B2(n_76),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_16),
.B1(n_32),
.B2(n_42),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_171),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_105),
.A2(n_74),
.B1(n_73),
.B2(n_69),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_42),
.B1(n_16),
.B2(n_32),
.Y(n_170)
);

AND2x4_ASAP7_75t_SL g171 ( 
.A(n_125),
.B(n_39),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_175),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_96),
.B(n_113),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_92),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_179),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_92),
.B(n_22),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_187),
.Y(n_199)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_112),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_181),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_188),
.C(n_189),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_116),
.A2(n_32),
.B1(n_16),
.B2(n_37),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_186),
.Y(n_201)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_22),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_114),
.B(n_37),
.C(n_22),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_108),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_216),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_205),
.A2(n_122),
.B1(n_130),
.B2(n_131),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_99),
.B(n_132),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_206),
.A2(n_211),
.B(n_178),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_99),
.B(n_134),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_148),
.B(n_108),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_156),
.A2(n_140),
.B1(n_107),
.B2(n_111),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_154),
.B1(n_159),
.B2(n_165),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_172),
.B(n_115),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_187),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_171),
.B(n_118),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_155),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_177),
.C(n_171),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_232),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_185),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_227),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_249),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_189),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_250),
.B(n_220),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_152),
.C(n_184),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_238),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_178),
.C(n_164),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_235),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_187),
.C(n_176),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_121),
.B1(n_107),
.B2(n_140),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_206),
.B1(n_186),
.B2(n_218),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_205),
.A2(n_204),
.B1(n_219),
.B2(n_216),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_240),
.A2(n_244),
.B1(n_253),
.B2(n_147),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_241),
.Y(n_276)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_190),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_245),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_211),
.A2(n_121),
.B1(n_110),
.B2(n_122),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_203),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_168),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_248),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_222),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_161),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

NAND2x1_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_118),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_251),
.A2(n_208),
.B1(n_217),
.B2(n_146),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_192),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_220),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_255),
.A2(n_275),
.B1(n_277),
.B2(n_225),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_230),
.A2(n_192),
.B1(n_200),
.B2(n_212),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_269),
.B1(n_274),
.B2(n_278),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_268),
.B(n_270),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_229),
.A2(n_221),
.B(n_212),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_210),
.B1(n_145),
.B2(n_202),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_231),
.A2(n_221),
.B(n_195),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_231),
.A2(n_245),
.B(n_240),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_266),
.B(n_270),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_226),
.A2(n_130),
.B1(n_210),
.B2(n_195),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_196),
.B1(n_214),
.B2(n_215),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_236),
.A2(n_213),
.B1(n_181),
.B2(n_173),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_228),
.A2(n_213),
.B1(n_175),
.B2(n_196),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_251),
.B1(n_237),
.B2(n_249),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_227),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_303),
.C(n_257),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_273),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_292),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_286),
.A2(n_288),
.B1(n_302),
.B2(n_306),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_287),
.A2(n_289),
.B1(n_258),
.B2(n_311),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_228),
.B1(n_243),
.B2(n_253),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_291),
.A2(n_301),
.B(n_265),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_278),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_299),
.Y(n_338)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_232),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_305),
.C(n_309),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_247),
.Y(n_298)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

INVx3_ASAP7_75t_SL g299 ( 
.A(n_259),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_263),
.B(n_248),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_300),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_250),
.B(n_224),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_259),
.A2(n_252),
.B1(n_235),
.B2(n_232),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_234),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_224),
.C(n_246),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_255),
.A2(n_238),
.B1(n_233),
.B2(n_250),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_260),
.A2(n_250),
.B1(n_225),
.B2(n_214),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_131),
.B1(n_100),
.B2(n_27),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_191),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_268),
.A2(n_242),
.B(n_215),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_277),
.A2(n_197),
.B1(n_179),
.B2(n_190),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_311),
.A2(n_269),
.B1(n_259),
.B2(n_264),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_197),
.C(n_220),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_275),
.C(n_160),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_271),
.B(n_37),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_313),
.B(n_305),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_300),
.B(n_276),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_314),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_316),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_317),
.A2(n_321),
.B1(n_285),
.B2(n_286),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_289),
.A2(n_299),
.B1(n_293),
.B2(n_288),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_320),
.A2(n_299),
.B1(n_310),
.B2(n_295),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_309),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_331),
.C(n_332),
.Y(n_351)
);

AOI22x1_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_262),
.B1(n_265),
.B2(n_261),
.Y(n_323)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_292),
.A2(n_262),
.B1(n_276),
.B2(n_271),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_324),
.A2(n_301),
.B1(n_308),
.B2(n_291),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_298),
.B(n_257),
.Y(n_325)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_325),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_330),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_158),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_318),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_SL g334 ( 
.A(n_312),
.B(n_100),
.Y(n_334)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_334),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_337),
.A2(n_284),
.B1(n_134),
.B2(n_33),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_294),
.Y(n_340)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_340),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_344),
.A2(n_353),
.B1(n_357),
.B2(n_321),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_364),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_336),
.A2(n_338),
.B(n_330),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_349),
.A2(n_354),
.B(n_366),
.Y(n_371)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_320),
.A2(n_290),
.B1(n_307),
.B2(n_304),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_336),
.A2(n_290),
.B(n_285),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_317),
.A2(n_284),
.B1(n_313),
.B2(n_40),
.Y(n_356)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_338),
.A2(n_31),
.B1(n_39),
.B2(n_2),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_359),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_335),
.A2(n_31),
.B1(n_39),
.B2(n_2),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_322),
.C(n_332),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_39),
.C(n_9),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_360),
.Y(n_370)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_339),
.Y(n_362)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_339),
.Y(n_363)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_323),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_367),
.Y(n_377)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_341),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_369),
.A2(n_373),
.B1(n_385),
.B2(n_356),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_376),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_352),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_353),
.A2(n_327),
.B1(n_324),
.B2(n_326),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_354),
.A2(n_323),
.B(n_327),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_374),
.A2(n_384),
.B(n_371),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_319),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_333),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_390),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_349),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_347),
.Y(n_394)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_367),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_380),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_331),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_383),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_345),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_329),
.B(n_340),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_344),
.A2(n_315),
.B1(n_328),
.B2(n_31),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_388),
.B(n_0),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_7),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_343),
.Y(n_391)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_391),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_395),
.Y(n_410)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_394),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_374),
.A2(n_348),
.B(n_342),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_352),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_396),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_397),
.A2(n_401),
.B1(n_387),
.B2(n_381),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_372),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_357),
.C(n_358),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_402),
.C(n_404),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_359),
.C(n_1),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_7),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_405),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_0),
.C(n_1),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_7),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_9),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_409),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_381),
.A2(n_9),
.B1(n_12),
.B2(n_3),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_369),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_4),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_412),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_390),
.Y(n_414)
);

AOI21x1_ASAP7_75t_L g433 ( 
.A1(n_414),
.A2(n_4),
.B(n_6),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_418),
.A2(n_422),
.B1(n_423),
.B2(n_6),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_400),
.A2(n_373),
.B1(n_387),
.B2(n_385),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_419),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_399),
.A2(n_375),
.B1(n_386),
.B2(n_389),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_407),
.A2(n_375),
.B1(n_388),
.B2(n_380),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_0),
.C(n_1),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_425),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_1),
.C(n_15),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_393),
.C(n_408),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_428),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_403),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_412),
.A2(n_407),
.B(n_396),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_429),
.A2(n_430),
.B(n_417),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_415),
.A2(n_404),
.B(n_402),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_410),
.B(n_3),
.Y(n_431)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_431),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_3),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_435),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_433),
.A2(n_420),
.B(n_425),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_434),
.B(n_416),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_421),
.B(n_4),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_419),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_437),
.B(n_423),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_439),
.Y(n_448)
);

FAx1_ASAP7_75t_SL g440 ( 
.A(n_426),
.B(n_422),
.CI(n_416),
.CON(n_440),
.SN(n_440)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_440),
.B(n_443),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_442),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_445),
.B(n_449),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_424),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_448),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_439),
.B(n_9),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_444),
.B(n_437),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_451),
.A2(n_457),
.B(n_15),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_438),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_458),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_440),
.A2(n_434),
.B(n_436),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_10),
.C(n_11),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_452),
.A2(n_450),
.B(n_446),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_459),
.B(n_460),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_457),
.A2(n_11),
.B(n_12),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_461),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_454),
.C(n_451),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_464),
.B(n_462),
.C(n_463),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_465),
.C(n_455),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_11),
.C(n_12),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_468),
.Y(n_469)
);


endmodule