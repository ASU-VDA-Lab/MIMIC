module fake_aes_1170_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
O2A1O1Ixp33_ASAP7_75t_SL g5 ( .A1(n_4), .A2(n_3), .B(n_1), .C(n_2), .Y(n_5) );
CKINVDCx6p67_ASAP7_75t_R g6 ( .A(n_3), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_7), .B(n_5), .Y(n_10) );
AOI211xp5_ASAP7_75t_SL g11 ( .A1(n_10), .A2(n_8), .B(n_9), .C(n_2), .Y(n_11) );
AOI21xp5_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_0), .B(n_1), .Y(n_12) );
OR2x2_ASAP7_75t_L g13 ( .A(n_12), .B(n_0), .Y(n_13) );
AND3x4_ASAP7_75t_L g14 ( .A(n_11), .B(n_0), .C(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
AOI22xp33_ASAP7_75t_SL g16 ( .A1(n_15), .A2(n_14), .B1(n_0), .B2(n_2), .Y(n_16) );
endmodule