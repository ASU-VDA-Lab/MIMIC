module fake_jpeg_28312_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_40),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_60),
.Y(n_62)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

CKINVDCx12_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_49),
.B1(n_54),
.B2(n_44),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_75),
.B1(n_22),
.B2(n_36),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_46),
.B1(n_54),
.B2(n_53),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_42),
.B1(n_20),
.B2(n_21),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_84),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_88),
.B1(n_86),
.B2(n_91),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_67),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_86),
.Y(n_96)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_87),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_2),
.Y(n_86)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_90),
.Y(n_102)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_5),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_97),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_18),
.B1(n_35),
.B2(n_34),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_6),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_102),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_92),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_7),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_93),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_108),
.B1(n_110),
.B2(n_107),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_110),
.B1(n_105),
.B2(n_109),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_115),
.B1(n_111),
.B2(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_120),
.B1(n_25),
.B2(n_10),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_83),
.B(n_26),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_23),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_16),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_27),
.A3(n_38),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_29),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_28),
.B1(n_79),
.B2(n_8),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_9),
.Y(n_129)
);


endmodule