module fake_jpeg_23290_n_228 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_29),
.B(n_2),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_21),
.C(n_31),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_19),
.B(n_33),
.C(n_20),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_50),
.A2(n_18),
.B(n_9),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_26),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_59),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_27),
.B1(n_24),
.B2(n_28),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_25),
.B1(n_18),
.B2(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_27),
.B1(n_35),
.B2(n_33),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_64),
.B1(n_67),
.B2(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_26),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_34),
.B1(n_29),
.B2(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_17),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_36),
.A2(n_34),
.B1(n_25),
.B2(n_5),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_3),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_80),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_34),
.B1(n_39),
.B2(n_43),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_25),
.B1(n_5),
.B2(n_6),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_86),
.B1(n_89),
.B2(n_91),
.Y(n_118)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_47),
.B1(n_46),
.B2(n_32),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_46),
.B1(n_47),
.B2(n_45),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_46),
.B1(n_32),
.B2(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_92),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_45),
.B1(n_44),
.B2(n_32),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_44),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_44),
.B1(n_32),
.B2(n_30),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_54),
.B1(n_71),
.B2(n_65),
.Y(n_121)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_51),
.A2(n_30),
.B1(n_18),
.B2(n_10),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_55),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_30),
.B1(n_18),
.B2(n_10),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_4),
.Y(n_123)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_109),
.Y(n_149)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_51),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_116),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_121),
.B1(n_94),
.B2(n_88),
.Y(n_144)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_77),
.B(n_73),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_49),
.C(n_65),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_125),
.Y(n_133)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_49),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_85),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_81),
.B(n_101),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_56),
.C(n_63),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_98),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_126),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_71),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_18),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_143),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_83),
.B(n_78),
.C(n_82),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_142),
.B(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_148),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_99),
.B1(n_103),
.B2(n_93),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_131),
.B1(n_130),
.B2(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_75),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_139),
.B(n_107),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_144),
.B1(n_146),
.B2(n_113),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_89),
.B(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_122),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_90),
.B1(n_96),
.B2(n_63),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_90),
.B(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_128),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_171),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_117),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_160),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_125),
.C(n_112),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_167),
.C(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_106),
.B1(n_146),
.B2(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_106),
.B1(n_123),
.B2(n_115),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_142),
.B1(n_141),
.B2(n_148),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_63),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_134),
.A2(n_119),
.B1(n_109),
.B2(n_4),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_138),
.A2(n_108),
.B(n_9),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_140),
.B(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_183),
.B1(n_171),
.B2(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_139),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_134),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_178),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_129),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_186),
.C(n_166),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_135),
.C(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_175),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_189),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_153),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_185),
.C(n_132),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_156),
.C(n_160),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_192),
.C(n_195),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_179),
.C(n_180),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_197),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_156),
.C(n_170),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_167),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_181),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_178),
.C(n_173),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_174),
.C(n_137),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_152),
.Y(n_207)
);

OA21x2_ASAP7_75t_SL g201 ( 
.A1(n_193),
.A2(n_172),
.B(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_207),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_205),
.C(n_184),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_194),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_161),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_202),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_15),
.C(n_16),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_11),
.B(n_12),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_215),
.B1(n_213),
.B2(n_14),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_209),
.A2(n_202),
.B1(n_200),
.B2(n_15),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_219),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_220),
.Y(n_223)
);

AOI211xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_212),
.B(n_210),
.C(n_16),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_216),
.C(n_9),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_223),
.B1(n_224),
.B2(n_222),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_226),
.Y(n_228)
);


endmodule