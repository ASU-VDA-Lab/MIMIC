module real_jpeg_26580_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_336, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_336;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx5_ASAP7_75t_L g114 ( 
.A(n_0),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_0),
.Y(n_119)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_0),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_1),
.A2(n_31),
.B1(n_33),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_1),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_1),
.A2(n_27),
.B1(n_35),
.B2(n_129),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_129),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_1),
.A2(n_65),
.B1(n_67),
.B2(n_129),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_2),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_2),
.B(n_30),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_2),
.B(n_33),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_2),
.A2(n_33),
.B(n_176),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_134),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_2),
.A2(n_62),
.B(n_65),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_2),
.B(n_90),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_2),
.A2(n_111),
.B1(n_114),
.B2(n_227),
.Y(n_230)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_4),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_4),
.A2(n_31),
.B1(n_33),
.B2(n_38),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_38),
.B1(n_65),
.B2(n_67),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_4),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_31),
.B1(n_33),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_7),
.A2(n_27),
.B1(n_35),
.B2(n_56),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_7),
.A2(n_56),
.B1(n_65),
.B2(n_67),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_8),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_131),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_8),
.A2(n_65),
.B1(n_67),
.B2(n_131),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_8),
.A2(n_27),
.B1(n_35),
.B2(n_131),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_31),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_9),
.A2(n_53),
.B1(n_65),
.B2(n_67),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_9),
.A2(n_27),
.B1(n_35),
.B2(n_53),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_10),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_10),
.A2(n_36),
.B1(n_65),
.B2(n_67),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_283)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_12),
.A2(n_27),
.B1(n_35),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_12),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_12),
.A2(n_31),
.B1(n_33),
.B2(n_136),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_136),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_12),
.A2(n_65),
.B1(n_67),
.B2(n_136),
.Y(n_227)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_15),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_97),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_95),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_82),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.C(n_76),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_20),
.A2(n_21),
.B1(n_72),
.B2(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_40),
.B1(n_41),
.B2(n_71),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_23),
.A2(n_39),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_23),
.A2(n_39),
.B1(n_142),
.B2(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_23),
.A2(n_267),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_24),
.B(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_24),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_24),
.A2(n_30),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_24),
.A2(n_87),
.B(n_287),
.Y(n_311)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_25),
.B(n_33),
.Y(n_148)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_27),
.B(n_134),
.CON(n_133),
.SN(n_133)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_29),
.A2(n_31),
.B1(n_133),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_30),
.B(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_31),
.A2(n_33),
.B1(n_50),
.B2(n_51),
.Y(n_58)
);

AOI32xp33_ASAP7_75t_L g175 ( 
.A1(n_31),
.A2(n_46),
.A3(n_49),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_34),
.A2(n_39),
.B(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_59),
.B2(n_70),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_43),
.B(n_59),
.C(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_54),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_44),
.A2(n_78),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_52),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_45),
.A2(n_57),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_45),
.A2(n_57),
.B1(n_128),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_45),
.A2(n_57),
.B1(n_159),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_45),
.A2(n_57),
.B1(n_80),
.B2(n_305),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_47),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g177 ( 
.A(n_47),
.B(n_50),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_47),
.A2(n_63),
.B(n_134),
.C(n_204),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_54),
.A2(n_90),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_59),
.A2(n_70),
.B1(n_77),
.B2(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_64),
.B(n_68),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_60),
.A2(n_68),
.B(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_60),
.A2(n_64),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_60),
.A2(n_184),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_60),
.A2(n_64),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_60),
.A2(n_64),
.B1(n_183),
.B2(n_202),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_60),
.A2(n_64),
.B1(n_106),
.B2(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_60),
.A2(n_124),
.B(n_260),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_106),
.B(n_107),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_64),
.B(n_134),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_65),
.Y(n_67)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_67),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_69),
.B(n_125),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_72),
.C(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_72),
.A2(n_319),
.B1(n_321),
.B2(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_72),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_76),
.B(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_77),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B(n_81),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_78),
.A2(n_81),
.B(n_91),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_315),
.A3(n_327),
.B1(n_333),
.B2(n_334),
.C(n_336),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_297),
.B(n_314),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_273),
.B(n_296),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_166),
.B(n_251),
.C(n_272),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_151),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_102),
.B(n_151),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_137),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_121),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_104),
.B(n_121),
.C(n_137),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_105),
.B(n_110),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_107),
.B(n_194),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_115),
.B(n_116),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_111),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_111),
.A2(n_219),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_111),
.A2(n_163),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_112),
.B(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_112),
.A2(n_117),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_112),
.A2(n_214),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_132),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_134),
.B(n_163),
.Y(n_232)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_146),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_139),
.B(n_144),
.C(n_146),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_149),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_157),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_152),
.A2(n_153),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_162),
.Y(n_189)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_164),
.B(n_213),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_250),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_243),
.B(n_249),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_195),
.B(n_242),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_185),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_170),
.B(n_185),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.C(n_181),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_171),
.A2(n_172),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_175),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_174),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_186),
.B(n_192),
.C(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_236),
.B(n_241),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_215),
.B(n_235),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_205),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_198),
.B(n_205),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_212),
.Y(n_220)
);

INVx11_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_223),
.B(n_234),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_217),
.B(n_221),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_229),
.B(n_233),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_252),
.B(n_253),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_270),
.B2(n_271),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_261),
.B2(n_262),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_262),
.C(n_271),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_265),
.C(n_269),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_275),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_295),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_288),
.B2(n_289),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_289),
.C(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_282),
.C(n_284),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_290),
.A2(n_291),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_293),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_291),
.A2(n_308),
.B(n_311),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_298),
.B(n_299),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_312),
.B2(n_313),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_307),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_307),
.C(n_313),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_317),
.C(n_323),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_306),
.A2(n_317),
.B1(n_318),
.B2(n_332),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_306),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_325),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_325),
.Y(n_334)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_324),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);


endmodule