module fake_jpeg_21806_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_8),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_29),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_31),
.B1(n_29),
.B2(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_14),
.Y(n_40)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_40),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_20),
.B1(n_21),
.B2(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_20),
.B1(n_21),
.B2(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_12),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_20),
.B1(n_14),
.B2(n_19),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_27),
.B1(n_36),
.B2(n_46),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_60),
.B1(n_47),
.B2(n_32),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_25),
.Y(n_54)
);

OR2x4_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_13),
.Y(n_69)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVxp33_ASAP7_75t_SL g67 ( 
.A(n_59),
.Y(n_67)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_36),
.B1(n_27),
.B2(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_31),
.B1(n_30),
.B2(n_36),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_37),
.B1(n_13),
.B2(n_18),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_23),
.B1(n_18),
.B2(n_35),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_18),
.B1(n_25),
.B2(n_16),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_38),
.B1(n_43),
.B2(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_63),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_49),
.C(n_50),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_70),
.C(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_52),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_22),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_74),
.B1(n_76),
.B2(n_60),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_60),
.B1(n_65),
.B2(n_69),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_32),
.B1(n_24),
.B2(n_3),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_81),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_86),
.B(n_66),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_56),
.B(n_60),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_84),
.B1(n_65),
.B2(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_68),
.C(n_74),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_92),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_93),
.B1(n_80),
.B2(n_84),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_77),
.B1(n_75),
.B2(n_70),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_77),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_84),
.B(n_24),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_90),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_94),
.A3(n_91),
.B1(n_6),
.B2(n_5),
.C1(n_8),
.C2(n_9),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_91),
.C(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_102),
.B(n_0),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.C(n_105),
.Y(n_106)
);

AOI31xp67_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_5),
.A3(n_1),
.B(n_3),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_101),
.C(n_99),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_106),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);


endmodule