module fake_aes_284_n_31 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_31);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_6), .Y(n_8) );
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_1), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_7), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
A2O1A1Ixp33_ASAP7_75t_L g14 ( .A1(n_10), .A2(n_0), .B(n_2), .C(n_3), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_12), .B(n_0), .Y(n_16) );
BUFx12f_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
INVx4_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_18), .B(n_13), .Y(n_19) );
NOR2x1p5_ASAP7_75t_L g20 ( .A(n_17), .B(n_12), .Y(n_20) );
BUFx8_ASAP7_75t_L g21 ( .A(n_15), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
OAI21xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_16), .B(n_14), .Y(n_24) );
OAI322xp33_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_9), .A3(n_16), .B1(n_18), .B2(n_14), .C1(n_20), .C2(n_21), .Y(n_25) );
AOI21xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_23), .B(n_0), .Y(n_26) );
A2O1A1Ixp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_3), .B(n_4), .C(n_5), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_27), .Y(n_28) );
NOR2x1_ASAP7_75t_L g29 ( .A(n_26), .B(n_7), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
AOI22xp33_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_5), .B1(n_29), .B2(n_28), .Y(n_31) );
endmodule