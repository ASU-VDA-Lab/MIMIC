module fake_jpeg_16212_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_70),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_2),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_62),
.Y(n_85)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_63),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_70),
.A2(n_59),
.B1(n_47),
.B2(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_87),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_52),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_48),
.B1(n_50),
.B2(n_60),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_48),
.B1(n_60),
.B2(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_54),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_56),
.B1(n_57),
.B2(n_51),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_90),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_46),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_51),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_100),
.C(n_5),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_54),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_3),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_105),
.B1(n_106),
.B2(n_96),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_80),
.B1(n_49),
.B2(n_78),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_116),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_23),
.B(n_42),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_97),
.B(n_104),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_114),
.A2(n_116),
.B1(n_113),
.B2(n_111),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_115),
.B1(n_103),
.B2(n_114),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_121),
.B(n_122),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_97),
.B(n_106),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_124),
.B(n_127),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_108),
.C(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_105),
.Y(n_134)
);

OAI21x1_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_88),
.B(n_120),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_129),
.B(n_9),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_110),
.B1(n_98),
.B2(n_108),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_133),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_25),
.B1(n_43),
.B2(n_41),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_21),
.B(n_39),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_136),
.C(n_133),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_137),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_138),
.B1(n_132),
.B2(n_28),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_139),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_131),
.B(n_22),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_17),
.B(n_38),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_16),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_27),
.Y(n_146)
);

AOI21x1_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_15),
.B(n_36),
.Y(n_147)
);

OAI321xp33_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_14),
.A3(n_34),
.B1(n_33),
.B2(n_32),
.C(n_30),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_40),
.B(n_29),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_13),
.B(n_10),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_150),
.B(n_9),
.Y(n_151)
);


endmodule