module fake_jpeg_14698_n_203 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_28),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_16),
.CON(n_39),
.SN(n_39)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_1),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_28),
.B(n_29),
.C(n_16),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_53),
.B(n_29),
.C(n_13),
.Y(n_58)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_48),
.B(n_49),
.Y(n_62)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_30),
.A2(n_20),
.B1(n_25),
.B2(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_22),
.B1(n_20),
.B2(n_14),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_27),
.A2(n_17),
.B1(n_13),
.B2(n_16),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_14),
.B1(n_25),
.B2(n_24),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_37),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_23),
.Y(n_86)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_60),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_30),
.B1(n_24),
.B2(n_22),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_40),
.B(n_25),
.Y(n_83)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_46),
.B1(n_54),
.B2(n_44),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_72),
.B1(n_81),
.B2(n_86),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_46),
.B1(n_44),
.B2(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_87),
.Y(n_90)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_83),
.B(n_86),
.Y(n_102)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_47),
.B1(n_33),
.B2(n_19),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_69),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_32),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_70),
.B(n_51),
.C(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_36),
.B1(n_66),
.B2(n_50),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_99),
.B1(n_101),
.B2(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_94),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_98),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_53),
.B(n_18),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_85),
.B1(n_82),
.B2(n_31),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_28),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_19),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_104),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_27),
.B1(n_40),
.B2(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_110),
.B(n_115),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_102),
.C(n_90),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_117),
.C(n_118),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_120),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_87),
.B1(n_51),
.B2(n_77),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_113),
.B1(n_114),
.B2(n_118),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_22),
.B(n_20),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_80),
.B(n_78),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_32),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_34),
.C(n_73),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_88),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_125),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_96),
.C(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_138),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_98),
.C(n_93),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_137),
.C(n_18),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_89),
.B1(n_97),
.B2(n_77),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_97),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_23),
.B(n_18),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_134),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_110),
.B1(n_120),
.B2(n_45),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_19),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_136),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_45),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_117),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_149),
.C(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_143),
.B(n_122),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_61),
.B1(n_73),
.B2(n_4),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_34),
.C(n_18),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_130),
.B(n_133),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_157),
.B(n_163),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_129),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_159),
.C(n_150),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_137),
.C(n_138),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_162),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_152),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_2),
.Y(n_174)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_171),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_175),
.C(n_176),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_140),
.B1(n_147),
.B2(n_141),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_141),
.B1(n_144),
.B2(n_151),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_3),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_26),
.C(n_21),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_161),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_179),
.A2(n_170),
.B1(n_173),
.B2(n_176),
.Y(n_186)
);

BUFx6f_ASAP7_75t_SL g180 ( 
.A(n_168),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_180),
.B(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_182),
.B(n_184),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_158),
.C(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_7),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_7),
.B(n_8),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_191),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_7),
.B(n_8),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_188),
.A3(n_194),
.B1(n_186),
.B2(n_193),
.C1(n_182),
.C2(n_21),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_198),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_26),
.Y(n_198)
);

AOI21x1_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_8),
.B(n_9),
.Y(n_199)
);

AOI321xp33_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_200),
.C(n_26),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_201),
.B(n_9),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_10),
.Y(n_203)
);


endmodule