module fake_jpeg_13342_n_437 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_437);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_437;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_25),
.B(n_10),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_55),
.B(n_50),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_56),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_62),
.Y(n_120)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx2_ASAP7_75t_SL g189 ( 
.A(n_60),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_18),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_65),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_66),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_67),
.Y(n_188)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_10),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_73),
.B(n_104),
.Y(n_143)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_97),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_27),
.B(n_7),
.C(n_16),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_45),
.C(n_44),
.Y(n_131)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_92),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_96),
.Y(n_135)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_98),
.B(n_100),
.Y(n_167)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_103),
.Y(n_121)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_23),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_108),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_105),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_106),
.B(n_107),
.Y(n_186)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

INVx11_ASAP7_75t_SL g109 ( 
.A(n_37),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_111),
.B(n_0),
.Y(n_142)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_29),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_113),
.Y(n_144)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_114),
.B(n_57),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_4),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_47),
.B1(n_48),
.B2(n_39),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_118),
.A2(n_125),
.B1(n_133),
.B2(n_134),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_124),
.B(n_142),
.C(n_147),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_81),
.A2(n_39),
.B1(n_48),
.B2(n_33),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_52),
.B1(n_45),
.B2(n_29),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_127),
.A2(n_132),
.B1(n_137),
.B2(n_145),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_53),
.B1(n_24),
.B2(n_30),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_128),
.A2(n_149),
.B1(n_157),
.B2(n_121),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_55),
.B(n_52),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_130),
.B(n_154),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_171),
.C(n_158),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_78),
.A2(n_44),
.B1(n_30),
.B2(n_24),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_67),
.A2(n_33),
.B1(n_21),
.B2(n_2),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_113),
.A2(n_21),
.B1(n_1),
.B2(n_3),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_84),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_94),
.A2(n_12),
.B1(n_16),
.B2(n_13),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_91),
.A2(n_11),
.B(n_13),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_101),
.B1(n_95),
.B2(n_114),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_61),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_152),
.A2(n_178),
.B1(n_180),
.B2(n_183),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_106),
.A2(n_17),
.B1(n_11),
.B2(n_13),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_66),
.A2(n_11),
.B1(n_76),
.B2(n_70),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_160),
.A2(n_176),
.B1(n_150),
.B2(n_181),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_71),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_163),
.B(n_169),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_91),
.B(n_57),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_110),
.B(n_108),
.C(n_66),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_110),
.A2(n_109),
.B1(n_75),
.B2(n_60),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_59),
.A2(n_46),
.B1(n_38),
.B2(n_41),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_59),
.A2(n_46),
.B1(n_38),
.B2(n_41),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_59),
.A2(n_58),
.B1(n_74),
.B2(n_87),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_185),
.B1(n_176),
.B2(n_188),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_59),
.A2(n_46),
.B1(n_38),
.B2(n_41),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_93),
.B(n_112),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_146),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_131),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_190),
.B(n_195),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_193),
.B(n_213),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_127),
.A2(n_137),
.B1(n_182),
.B2(n_167),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_194),
.A2(n_219),
.B1(n_226),
.B2(n_237),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_121),
.B1(n_151),
.B2(n_162),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_196),
.A2(n_202),
.B1(n_209),
.B2(n_214),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_197),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_199),
.B(n_200),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_120),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_159),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_201),
.B(n_242),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_144),
.B(n_141),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_203),
.B(n_205),
.Y(n_268)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_117),
.B(n_138),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_208),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_186),
.B1(n_175),
.B2(n_139),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_138),
.B(n_179),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_210),
.B(n_211),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_140),
.B(n_139),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_175),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_212),
.B(n_220),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_136),
.A2(n_171),
.B1(n_161),
.B2(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_158),
.A2(n_129),
.B(n_189),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_216),
.Y(n_281)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_136),
.Y(n_217)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_217),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_158),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_218),
.B(n_221),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_155),
.A2(n_161),
.B1(n_174),
.B2(n_166),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_119),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_148),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_116),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_153),
.A2(n_164),
.B1(n_170),
.B2(n_148),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_119),
.Y(n_225)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_166),
.A2(n_177),
.B1(n_165),
.B2(n_156),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_122),
.Y(n_228)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

BUFx12_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_150),
.B(n_122),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_153),
.A2(n_164),
.B1(n_170),
.B2(n_181),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_247),
.B(n_202),
.Y(n_255)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_177),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_123),
.Y(n_234)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_234),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_165),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_123),
.Y(n_236)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_236),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_168),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_126),
.B(n_143),
.C(n_131),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_244),
.C(n_191),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_168),
.B(n_143),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_245),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_143),
.B(n_131),
.C(n_159),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_184),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_251),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_127),
.A2(n_38),
.B1(n_46),
.B2(n_59),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_116),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_124),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_249),
.B(n_250),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_124),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_184),
.B(n_124),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_227),
.A2(n_213),
.B1(n_242),
.B2(n_241),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_254),
.A2(n_274),
.B1(n_284),
.B2(n_259),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_193),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_201),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_262),
.B(n_264),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_229),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_209),
.A2(n_193),
.B1(n_218),
.B2(n_207),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_266),
.A2(n_248),
.B1(n_240),
.B2(n_234),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_271),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g271 ( 
.A(n_190),
.B(n_244),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_227),
.A2(n_206),
.B1(n_224),
.B2(n_246),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_191),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_278),
.B(n_292),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_204),
.A2(n_243),
.B1(n_237),
.B2(n_193),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_238),
.B(n_192),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.C(n_216),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_225),
.B(n_239),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_214),
.C(n_230),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_295),
.C(n_300),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_253),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_235),
.B1(n_236),
.B2(n_221),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_296),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_233),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_303),
.Y(n_340)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_260),
.Y(n_299)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_273),
.C(n_265),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_223),
.B(n_228),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_302),
.A2(n_324),
.B(n_275),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_215),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_232),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_306),
.B(n_309),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_273),
.B(n_217),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_307),
.B(n_311),
.Y(n_337)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_310),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_198),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_312),
.A2(n_313),
.B1(n_288),
.B2(n_263),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_272),
.A2(n_208),
.B1(n_197),
.B2(n_229),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_271),
.C(n_258),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_267),
.C(n_268),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_222),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_272),
.B(n_256),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_323),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_318),
.A2(n_284),
.B1(n_270),
.B2(n_259),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_287),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_319),
.B(n_321),
.Y(n_339)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_261),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_283),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_322),
.B(n_325),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_256),
.B(n_258),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_274),
.A2(n_288),
.B1(n_279),
.B2(n_285),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_257),
.B(n_269),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_327),
.A2(n_338),
.B(n_343),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_290),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_344),
.C(n_293),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_331),
.A2(n_347),
.B1(n_348),
.B2(n_313),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_315),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_335),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_301),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_316),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_297),
.A2(n_279),
.B(n_276),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_297),
.A2(n_275),
.B(n_276),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_264),
.C(n_252),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_317),
.A2(n_280),
.B(n_285),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_345),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_318),
.A2(n_307),
.B1(n_303),
.B2(n_298),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_295),
.A2(n_286),
.B1(n_289),
.B2(n_263),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_349),
.B(n_370),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_359),
.C(n_368),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_294),
.Y(n_351)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_351),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_352),
.B(n_358),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_342),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_366),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_331),
.A2(n_347),
.B1(n_346),
.B2(n_327),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_356),
.Y(n_379)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_330),
.Y(n_355)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_330),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_338),
.A2(n_312),
.B1(n_302),
.B2(n_316),
.Y(n_357)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_357),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_330),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_304),
.C(n_323),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_360),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_345),
.A2(n_310),
.B1(n_308),
.B2(n_305),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_361),
.A2(n_363),
.B1(n_364),
.B2(n_333),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_335),
.A2(n_299),
.B1(n_319),
.B2(n_325),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_343),
.A2(n_311),
.B1(n_321),
.B2(n_322),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_320),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_315),
.C(n_280),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_328),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_329),
.B(n_289),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_357),
.A2(n_341),
.B(n_344),
.Y(n_373)
);

AND2x2_ASAP7_75t_SL g395 ( 
.A(n_373),
.B(n_385),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_378),
.C(n_368),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_334),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_367),
.A2(n_337),
.B(n_340),
.Y(n_381)
);

AO21x1_ASAP7_75t_L g397 ( 
.A1(n_381),
.A2(n_365),
.B(n_360),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_351),
.B(n_342),
.Y(n_382)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_382),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_326),
.Y(n_384)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_363),
.A2(n_348),
.B1(n_340),
.B2(n_339),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_386),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_390),
.B(n_397),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_356),
.Y(n_391)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_391),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_377),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_392),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_383),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_394),
.Y(n_404)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_380),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g396 ( 
.A(n_381),
.B(n_367),
.CI(n_366),
.CON(n_396),
.SN(n_396)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_396),
.B(n_373),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_369),
.C(n_365),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_401),
.C(n_375),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_387),
.A2(n_362),
.B1(n_355),
.B2(n_358),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_400),
.A2(n_379),
.B(n_371),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_354),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_401),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_400),
.A2(n_379),
.B(n_387),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_406),
.A2(n_371),
.B(n_385),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_399),
.B(n_372),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_410),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_409),
.B(n_390),
.C(n_398),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_394),
.Y(n_411)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_411),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_414),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_403),
.B(n_389),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_415),
.B(n_410),
.C(n_395),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_405),
.A2(n_388),
.B1(n_386),
.B2(n_376),
.Y(n_417)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_417),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_418),
.A2(n_419),
.B1(n_397),
.B2(n_409),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_378),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_420),
.B(n_422),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_421),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_395),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_404),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_416),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_427),
.B(n_429),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_412),
.C(n_395),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_425),
.C(n_422),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_430),
.Y(n_433)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g431 ( 
.A1(n_428),
.A2(n_383),
.B(n_388),
.C(n_391),
.D(n_421),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_431),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_434),
.A2(n_432),
.B(n_427),
.Y(n_435)
);

BUFx24_ASAP7_75t_SL g436 ( 
.A(n_435),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_433),
.C(n_408),
.Y(n_437)
);


endmodule