module fake_jpeg_10580_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_9),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_17),
.B1(n_20),
.B2(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_28),
.B1(n_20),
.B2(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_25),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_48),
.Y(n_52)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_15),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_27),
.B1(n_18),
.B2(n_33),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_34),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_21),
.C(n_23),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_12),
.C(n_15),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_59),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_30),
.B1(n_17),
.B2(n_20),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_65),
.B1(n_69),
.B2(n_73),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_30),
.B1(n_17),
.B2(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_68),
.Y(n_84)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_20),
.B1(n_28),
.B2(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_40),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_36),
.B(n_35),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_28),
.B1(n_35),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_28),
.B1(n_16),
.B2(n_29),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_26),
.B1(n_34),
.B2(n_32),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_47),
.B1(n_41),
.B2(n_31),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_90),
.B1(n_95),
.B2(n_111),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_79),
.B(n_86),
.C(n_27),
.Y(n_143)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_88),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_83),
.A2(n_111),
.B(n_82),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_34),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_106),
.B(n_77),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_47),
.B1(n_40),
.B2(n_39),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_91),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_26),
.B1(n_23),
.B2(n_32),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_93),
.A2(n_49),
.B1(n_16),
.B2(n_33),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_98),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_40),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_99),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_39),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_39),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_109),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_104),
.Y(n_132)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_107),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_23),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_19),
.B1(n_32),
.B2(n_21),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_24),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_33),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_114),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_33),
.B1(n_27),
.B2(n_18),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_60),
.B(n_57),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_116),
.B(n_137),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_71),
.B1(n_64),
.B2(n_57),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_83),
.B1(n_103),
.B2(n_107),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_16),
.B(n_29),
.C(n_49),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_106),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_80),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_136),
.B1(n_141),
.B2(n_144),
.Y(n_167)
);

AOI22x1_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_115),
.B1(n_90),
.B2(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_86),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_96),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_11),
.Y(n_174)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_79),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_78),
.A2(n_60),
.B1(n_27),
.B2(n_18),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_146),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_178),
.B1(n_156),
.B2(n_168),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_148),
.B(n_158),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_156),
.B1(n_176),
.B2(n_118),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_146),
.A2(n_95),
.B1(n_108),
.B2(n_80),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_163),
.B1(n_164),
.B2(n_172),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_131),
.B1(n_128),
.B2(n_135),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_151),
.A2(n_160),
.B1(n_168),
.B2(n_136),
.Y(n_185)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_157),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_162),
.B(n_164),
.Y(n_184)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_129),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_95),
.B1(n_81),
.B2(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_161),
.B(n_165),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_86),
.B1(n_115),
.B2(n_92),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_115),
.B(n_114),
.C(n_106),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_169),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_92),
.B1(n_101),
.B2(n_89),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

BUFx4f_ASAP7_75t_SL g170 ( 
.A(n_133),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_89),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_1),
.B(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_119),
.A2(n_85),
.B1(n_102),
.B2(n_91),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_179),
.Y(n_209)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_119),
.B(n_85),
.Y(n_180)
);

NOR2xp67_ASAP7_75t_R g197 ( 
.A(n_180),
.B(n_155),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_182),
.B(n_186),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_179),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_126),
.B1(n_142),
.B2(n_139),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_205),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_125),
.B1(n_116),
.B2(n_127),
.Y(n_192)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_180),
.A2(n_124),
.B1(n_141),
.B2(n_125),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_196),
.B(n_197),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_143),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_129),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_123),
.Y(n_202)
);

AO22x1_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_139),
.B1(n_123),
.B2(n_118),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_149),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_147),
.A2(n_127),
.B1(n_138),
.B2(n_137),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_166),
.A2(n_85),
.B1(n_140),
.B2(n_133),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_211),
.B(n_14),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_150),
.A2(n_133),
.B1(n_110),
.B2(n_121),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_212),
.B1(n_3),
.B2(n_4),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_175),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_170),
.C(n_169),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_181),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_214),
.B(n_215),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

AOI32xp33_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_175),
.A3(n_171),
.B1(n_165),
.B2(n_161),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_219),
.A2(n_224),
.B(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_226),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_153),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_229),
.C(n_230),
.Y(n_244)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_152),
.Y(n_227)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_193),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_170),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_169),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_234),
.C(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_207),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_193),
.A2(n_1),
.B(n_2),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_212),
.B1(n_195),
.B2(n_211),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_157),
.C(n_3),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_186),
.B(n_157),
.Y(n_236)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_1),
.C(n_3),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_239),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_260)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_185),
.B1(n_182),
.B2(n_188),
.Y(n_246)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_235),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_245),
.B(n_247),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_246),
.A2(n_248),
.B1(n_251),
.B2(n_254),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_204),
.B1(n_194),
.B2(n_208),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_260),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_203),
.B1(n_196),
.B2(n_184),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_216),
.A2(n_203),
.B1(n_184),
.B2(n_200),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_241),
.B1(n_221),
.B2(n_226),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_200),
.B1(n_189),
.B2(n_209),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_10),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_257),
.C(n_229),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_230),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_218),
.Y(n_264)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_220),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_228),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_220),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_239),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_269),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_276),
.C(n_277),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_281),
.B(n_267),
.Y(n_292)
);

OAI31xp33_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_240),
.A3(n_225),
.B(n_232),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_242),
.B(n_263),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_231),
.C(n_234),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_251),
.C(n_255),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_282),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_233),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_283),
.A2(n_222),
.B1(n_6),
.B2(n_7),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_250),
.B(n_262),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_286),
.A2(n_298),
.B(n_265),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_283),
.A2(n_248),
.B(n_253),
.C(n_250),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_292),
.B1(n_265),
.B2(n_279),
.Y(n_307)
);

AO22x1_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_242),
.B1(n_247),
.B2(n_260),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_252),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_294),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_261),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_271),
.C(n_276),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_237),
.B(n_14),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_280),
.Y(n_301)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_304),
.C(n_285),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_296),
.C(n_290),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_266),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_308),
.Y(n_320)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_268),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_287),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_270),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_312),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_313),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_316),
.C(n_320),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_295),
.B1(n_284),
.B2(n_288),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_321),
.B1(n_309),
.B2(n_301),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_289),
.C(n_287),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_291),
.B1(n_299),
.B2(n_269),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_323),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_303),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_325),
.B(n_327),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_302),
.C(n_308),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_313),
.B1(n_321),
.B2(n_297),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_298),
.B(n_306),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_319),
.B(n_318),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_328),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_334),
.B(n_330),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_325),
.B(n_320),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_4),
.B(n_7),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_7),
.B(n_9),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_9),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_9),
.Y(n_339)
);


endmodule