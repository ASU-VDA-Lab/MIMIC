module fake_jpeg_30242_n_220 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_31),
.B(n_26),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_19),
.Y(n_55)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.C(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_49),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_64),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_46),
.B1(n_44),
.B2(n_40),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_68),
.B1(n_73),
.B2(n_79),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_32),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_77),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_21),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_27),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_31),
.B1(n_25),
.B2(n_27),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_19),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_27),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_87),
.Y(n_131)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_81),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_94),
.Y(n_129)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_99),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_27),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_79),
.B(n_57),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_80),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_15),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_107),
.B(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_11),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_78),
.B1(n_70),
.B2(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_87),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_60),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_130),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_94),
.B(n_100),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_87),
.B(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_70),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_3),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_4),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_133),
.A2(n_122),
.B(n_123),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_110),
.B1(n_102),
.B2(n_106),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_149),
.B1(n_120),
.B2(n_117),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_91),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_150),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_89),
.C(n_92),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_142),
.C(n_137),
.Y(n_166)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_85),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_14),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_96),
.B1(n_111),
.B2(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_113),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_84),
.B(n_108),
.C(n_105),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_84),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_154),
.B(n_156),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_155),
.A2(n_126),
.B1(n_134),
.B2(n_117),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_6),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_171),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_169),
.B1(n_170),
.B2(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_144),
.C(n_143),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_128),
.B1(n_120),
.B2(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_115),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_152),
.B(n_138),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_174),
.A2(n_181),
.B(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_179),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_185),
.C(n_162),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_152),
.B(n_149),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_139),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_172),
.B1(n_165),
.B2(n_163),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_139),
.C(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_153),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_196),
.C(n_179),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_181),
.B(n_182),
.Y(n_200)
);

NAND4xp25_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_172),
.C(n_164),
.D(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_174),
.B(n_175),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_164),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_186),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_168),
.C(n_167),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_198),
.C(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_203),
.B(n_188),
.Y(n_205)
);

OAI322xp33_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_183),
.A3(n_159),
.B1(n_168),
.B2(n_151),
.C1(n_129),
.C2(n_115),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_196),
.B(n_170),
.Y(n_209)
);

AO21x1_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_159),
.B(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

NAND4xp25_ASAP7_75t_SL g206 ( 
.A(n_203),
.B(n_8),
.C(n_9),
.D(n_193),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_190),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_209),
.B(n_116),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_135),
.C(n_134),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_198),
.B1(n_192),
.B2(n_197),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_211),
.B(n_212),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_207),
.B(n_205),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_216),
.B(n_116),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_135),
.B(n_145),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

AOI21x1_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_218),
.B(n_116),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_145),
.Y(n_220)
);


endmodule