module fake_jpeg_22728_n_335 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_18),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_43),
.Y(n_53)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_19),
.B1(n_21),
.B2(n_30),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_21),
.B1(n_43),
.B2(n_25),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_24),
.B(n_34),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_33),
.B(n_24),
.C(n_34),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_19),
.B1(n_21),
.B2(n_20),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_67),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_19),
.B1(n_21),
.B2(n_20),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_30),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_11),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_65),
.A3(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_74),
.A2(n_61),
.B1(n_32),
.B2(n_39),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_43),
.B1(n_25),
.B2(n_20),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_92),
.B1(n_56),
.B2(n_61),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_81),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_88),
.Y(n_118)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_94),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_93),
.B(n_18),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_65),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_32),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_32),
.C(n_31),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_38),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_26),
.Y(n_99)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_115),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_111),
.B(n_42),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_39),
.Y(n_114)
);

NAND2x1_ASAP7_75t_SL g152 ( 
.A(n_114),
.B(n_42),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_116),
.B(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_127),
.B1(n_74),
.B2(n_90),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_94),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_68),
.B(n_65),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_83),
.B(n_95),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_77),
.B1(n_75),
.B2(n_87),
.Y(n_130)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_122),
.A2(n_60),
.B1(n_45),
.B2(n_89),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_70),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_101),
.B(n_116),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_45),
.B1(n_60),
.B2(n_64),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_134),
.B1(n_120),
.B2(n_106),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_152),
.B(n_154),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_139),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_142),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_143),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_83),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_150),
.C(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_148),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_84),
.C(n_80),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_101),
.B(n_126),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_73),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_86),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_125),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_114),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_0),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_158),
.A2(n_93),
.B(n_26),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_171),
.B1(n_191),
.B2(n_130),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_144),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_166),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_182),
.B(n_138),
.Y(n_208)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_173),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_143),
.B1(n_156),
.B2(n_131),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_156),
.A2(n_110),
.B1(n_125),
.B2(n_124),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_174),
.A2(n_183),
.B(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_147),
.B(n_145),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_138),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_132),
.A2(n_102),
.B(n_100),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_161),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_102),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_117),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_100),
.C(n_103),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_148),
.A2(n_103),
.B1(n_104),
.B2(n_128),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_42),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_205),
.B1(n_221),
.B2(n_170),
.Y(n_227)
);

BUFx12f_ASAP7_75t_SL g195 ( 
.A(n_168),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_195),
.A2(n_218),
.B1(n_152),
.B2(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_198),
.B(n_199),
.Y(n_230)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_203),
.Y(n_228)
);

BUFx12_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_136),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_22),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_140),
.B(n_141),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_153),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_215),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_187),
.Y(n_225)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_211),
.Y(n_236)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_219),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_154),
.Y(n_215)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_170),
.A2(n_154),
.B1(n_152),
.B2(n_136),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_172),
.C(n_192),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_226),
.C(n_243),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_229),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_173),
.C(n_169),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_234),
.B1(n_240),
.B2(n_218),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_174),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_232),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_233),
.B(n_211),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_160),
.B1(n_175),
.B2(n_181),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_181),
.B1(n_162),
.B2(n_179),
.Y(n_235)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_165),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_245),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_221),
.A2(n_162),
.B1(n_178),
.B2(n_190),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_242),
.A2(n_246),
.B(n_202),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_183),
.C(n_184),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_215),
.C(n_205),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_247),
.C(n_46),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_158),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_59),
.C(n_149),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_204),
.B(n_197),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_248),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_250),
.B(n_237),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_196),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_209),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_259),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_193),
.B1(n_213),
.B2(n_220),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_247),
.B1(n_243),
.B2(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_265),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_208),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_268),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_242),
.A2(n_149),
.B1(n_104),
.B2(n_81),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_222),
.B1(n_50),
.B2(n_58),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_122),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_266),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_86),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_76),
.C(n_58),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_225),
.B(n_46),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_246),
.B(n_244),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_283),
.B(n_268),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_273),
.B(n_0),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_263),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_229),
.B1(n_223),
.B2(n_245),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_253),
.B1(n_23),
.B2(n_35),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_223),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_285),
.C(n_249),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_259),
.A2(n_258),
.B(n_250),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_46),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_249),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_299),
.C(n_269),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_270),
.B1(n_285),
.B2(n_274),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_251),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_288),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_282),
.B(n_280),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_294),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_261),
.B(n_267),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_290),
.A2(n_278),
.B(n_284),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_295),
.B(n_296),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_297),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_256),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_253),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_12),
.Y(n_298)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_23),
.B(n_35),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_76),
.C(n_58),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_12),
.C(n_16),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_304),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_269),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_29),
.B(n_10),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_295),
.C(n_76),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_298),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_311),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_273),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_286),
.Y(n_313)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_311),
.B(n_307),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_319),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_292),
.C(n_300),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_314),
.A2(n_316),
.B(n_317),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_318),
.C(n_6),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_301),
.A2(n_50),
.B(n_23),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_1),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_50),
.C(n_29),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_318),
.B1(n_320),
.B2(n_13),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_310),
.A3(n_9),
.B1(n_11),
.B2(n_16),
.C1(n_5),
.C2(n_6),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_327),
.A3(n_329),
.B1(n_15),
.B2(n_2),
.C1(n_3),
.C2(n_4),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_8),
.B(n_15),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_326),
.B(n_5),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_328),
.B1(n_2),
.B2(n_3),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_5),
.A3(n_15),
.B1(n_14),
.B2(n_11),
.C1(n_16),
.C2(n_4),
.Y(n_329)
);

AOI321xp33_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_331),
.A3(n_332),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_3),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_4),
.Y(n_335)
);


endmodule