module fake_ibex_1421_n_3180 (n_151, n_85, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_568, n_52, n_448, n_99, n_466, n_269, n_156, n_570, n_126, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_558, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_267, n_245, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3180);

input n_151;
input n_85;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3180;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_3168;
wire n_884;
wire n_667;
wire n_2396;
wire n_3135;
wire n_850;
wire n_3175;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_2995;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2436;
wire n_1663;
wire n_2333;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1960;
wire n_1723;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_2373;
wire n_630;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_2723;
wire n_1616;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_3117;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2573;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_594;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_944;
wire n_3003;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2979;
wire n_2376;
wire n_2476;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3167;
wire n_997;
wire n_2308;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2875;
wire n_2684;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_2997;
wire n_1349;
wire n_961;
wire n_991;
wire n_634;
wire n_1331;
wire n_1223;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_2619;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_2862;
wire n_3100;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_604;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_595;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_839;
wire n_768;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2251;
wire n_722;
wire n_2012;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_2818;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3011;
wire n_818;
wire n_1167;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_1256;
wire n_2798;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3109;
wire n_1961;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_3104;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3035;
wire n_1029;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_632;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_635;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2303;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3114;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2324;
wire n_2738;
wire n_2246;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_2282;
wire n_970;
wire n_2673;
wire n_2676;
wire n_921;
wire n_2430;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;

BUFx3_ASAP7_75t_L g589 ( 
.A(n_548),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_571),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_539),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_172),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_374),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_429),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_291),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_64),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_360),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_455),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_343),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_475),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_183),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_181),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_152),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_266),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_374),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_573),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_131),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_579),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_400),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_74),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_116),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_441),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_223),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_428),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_351),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_65),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_373),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_343),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_387),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_280),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_52),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_460),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_268),
.Y(n_623)
);

BUFx5_ASAP7_75t_L g624 ( 
.A(n_26),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_576),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_163),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_14),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_547),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_263),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_155),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_585),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_48),
.Y(n_632)
);

NOR2xp67_ASAP7_75t_L g633 ( 
.A(n_159),
.B(n_115),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_540),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_141),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_423),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_331),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_248),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_57),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_527),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_106),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_391),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_485),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_575),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_234),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_96),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_554),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_221),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_284),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_57),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_347),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_415),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_157),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_276),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_577),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_131),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_562),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_299),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_534),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_192),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_201),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_97),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_314),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_544),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_532),
.Y(n_665)
);

NOR2xp67_ASAP7_75t_L g666 ( 
.A(n_436),
.B(n_331),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_502),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_10),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_446),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_263),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_369),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_317),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_299),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_284),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_253),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_264),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_493),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_553),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_157),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_552),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_46),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_542),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_351),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_254),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_317),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_470),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_153),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_42),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_235),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_565),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_191),
.Y(n_691)
);

CKINVDCx16_ASAP7_75t_R g692 ( 
.A(n_237),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_191),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_561),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_302),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_258),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_219),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_232),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_567),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_588),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_454),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_405),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_327),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_574),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_528),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_523),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_429),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_104),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_275),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_550),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_556),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_407),
.B(n_489),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_147),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_243),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_321),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_46),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_60),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_202),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_526),
.Y(n_719)
);

BUFx2_ASAP7_75t_SL g720 ( 
.A(n_525),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_583),
.B(n_560),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_207),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_111),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_337),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_484),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_543),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_180),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_185),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_270),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_298),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_380),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_521),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_129),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_430),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_68),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_529),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_16),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_545),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_6),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_486),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_460),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_119),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_372),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_308),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_125),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_304),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_101),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_533),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_500),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_329),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_490),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_524),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_458),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_572),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_110),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_266),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_430),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_109),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_584),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_242),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_563),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_120),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_494),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_146),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_488),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_221),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_438),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_52),
.Y(n_768)
);

CKINVDCx14_ASAP7_75t_R g769 ( 
.A(n_330),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_172),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_198),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_272),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_369),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_133),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_582),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_88),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_241),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_255),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_87),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_178),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_31),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_363),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_282),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_511),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_444),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_338),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_220),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_518),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_11),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_16),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_402),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_222),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_217),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_304),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_320),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_101),
.B(n_457),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_370),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_325),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_148),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_569),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_18),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_405),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_426),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_587),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_177),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_426),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_279),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_273),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_49),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_277),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_288),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_119),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_332),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_8),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_201),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_280),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_214),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_530),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_421),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_419),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_69),
.Y(n_821)
);

BUFx10_ASAP7_75t_L g822 ( 
.A(n_22),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_558),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_438),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_461),
.Y(n_825)
);

CKINVDCx16_ASAP7_75t_R g826 ( 
.A(n_488),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_233),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_440),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_224),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_385),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_246),
.Y(n_831)
);

BUFx5_ASAP7_75t_L g832 ( 
.A(n_102),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_79),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_564),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_20),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_321),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_506),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_380),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_36),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_258),
.Y(n_840)
);

BUFx10_ASAP7_75t_L g841 ( 
.A(n_536),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_35),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_89),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_77),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_134),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_586),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_452),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_295),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_463),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_238),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_169),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_195),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_238),
.Y(n_853)
);

CKINVDCx16_ASAP7_75t_R g854 ( 
.A(n_487),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_281),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_566),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_43),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_73),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_123),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_475),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_290),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_581),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_236),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_559),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_330),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_166),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_551),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_165),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_190),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_499),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_143),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_41),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_72),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_14),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_555),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_440),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_259),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_522),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_549),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_400),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_176),
.B(n_82),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_310),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_309),
.Y(n_883)
);

CKINVDCx16_ASAP7_75t_R g884 ( 
.A(n_102),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_409),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_466),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_557),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_181),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_231),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_149),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_10),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_160),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_261),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_546),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_94),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_62),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_399),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_328),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_312),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_421),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_11),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_97),
.Y(n_902)
);

BUFx8_ASAP7_75t_SL g903 ( 
.A(n_128),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_350),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_38),
.Y(n_905)
);

BUFx5_ASAP7_75t_L g906 ( 
.A(n_570),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_227),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_228),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_381),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_80),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_222),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_354),
.Y(n_912)
);

CKINVDCx16_ASAP7_75t_R g913 ( 
.A(n_486),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_456),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_146),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_189),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_313),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_260),
.B(n_470),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_568),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_305),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_95),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_541),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_39),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_13),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_39),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_164),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_27),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_504),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_88),
.Y(n_929)
);

OAI22x1_ASAP7_75t_R g930 ( 
.A1(n_595),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_657),
.Y(n_931)
);

BUFx12f_ASAP7_75t_L g932 ( 
.A(n_675),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_659),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_659),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_622),
.B(n_0),
.Y(n_935)
);

BUFx12f_ASAP7_75t_L g936 ( 
.A(n_675),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_661),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_661),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_723),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_675),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_723),
.Y(n_941)
);

INVx6_ASAP7_75t_L g942 ( 
.A(n_657),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_624),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_733),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_733),
.B(n_1),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_773),
.Y(n_946)
);

OAI22x1_ASAP7_75t_L g947 ( 
.A1(n_616),
.A2(n_619),
.B1(n_623),
.B2(n_618),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_659),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_819),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_769),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_808),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_594),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_736),
.B(n_2),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_592),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_736),
.B(n_867),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_907),
.B(n_867),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_636),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_613),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_830),
.B(n_4),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_659),
.Y(n_960)
);

OA21x2_ASAP7_75t_L g961 ( 
.A1(n_748),
.A2(n_505),
.B(n_503),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_670),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_636),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_908),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_688),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_648),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_641),
.B(n_7),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_624),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_648),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_641),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_624),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_688),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_903),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_604),
.B(n_8),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_649),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_740),
.B(n_9),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_648),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_596),
.B(n_9),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_674),
.Y(n_979)
);

XNOR2x2_ASAP7_75t_L g980 ( 
.A(n_881),
.B(n_12),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_649),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_688),
.Y(n_982)
);

AOI22x1_ASAP7_75t_SL g983 ( 
.A1(n_595),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_722),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_624),
.Y(n_985)
);

BUFx8_ASAP7_75t_L g986 ( 
.A(n_624),
.Y(n_986)
);

OA21x2_ASAP7_75t_L g987 ( 
.A1(n_748),
.A2(n_508),
.B(n_507),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_683),
.Y(n_988)
);

OA21x2_ASAP7_75t_L g989 ( 
.A1(n_775),
.A2(n_510),
.B(n_509),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_624),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_624),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_832),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_683),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_662),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_674),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_674),
.Y(n_996)
);

OA21x2_ASAP7_75t_L g997 ( 
.A1(n_775),
.A2(n_513),
.B(n_512),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_674),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_728),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_692),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_1000)
);

AND2x2_ASAP7_75t_SL g1001 ( 
.A(n_606),
.B(n_514),
.Y(n_1001)
);

BUFx8_ASAP7_75t_SL g1002 ( 
.A(n_903),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_790),
.B(n_19),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_845),
.Y(n_1004)
);

INVx6_ASAP7_75t_L g1005 ( 
.A(n_657),
.Y(n_1005)
);

INVx6_ASAP7_75t_L g1006 ( 
.A(n_841),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_832),
.Y(n_1007)
);

CKINVDCx16_ASAP7_75t_R g1008 ( 
.A(n_826),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_854),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_728),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_813),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_722),
.Y(n_1012)
);

AND2x2_ASAP7_75t_SL g1013 ( 
.A(n_608),
.B(n_631),
.Y(n_1013)
);

INVx5_ASAP7_75t_L g1014 ( 
.A(n_841),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_859),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_841),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_722),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_859),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_864),
.A2(n_516),
.B(n_515),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_893),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_893),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_845),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_832),
.Y(n_1023)
);

NOR2x1_ASAP7_75t_L g1024 ( 
.A(n_615),
.B(n_517),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_845),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_832),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_589),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_914),
.Y(n_1028)
);

INVx5_ASAP7_75t_L g1029 ( 
.A(n_589),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_832),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_655),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_929),
.B(n_597),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_590),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_665),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1014),
.B(n_616),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_967),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_968),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_971),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_967),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_937),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_950),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_985),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_938),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_939),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_941),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_1002),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_990),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_1013),
.B(n_928),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_1013),
.B(n_928),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_944),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1014),
.B(n_618),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_991),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_992),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_950),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_942),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1007),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_946),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_940),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_952),
.B(n_958),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_1008),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1023),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_986),
.B(n_906),
.Y(n_1062)
);

CKINVDCx6p67_ASAP7_75t_R g1063 ( 
.A(n_932),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_965),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_951),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_SL g1066 ( 
.A(n_1001),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1026),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_965),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_945),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_942),
.Y(n_1070)
);

CKINVDCx6p67_ASAP7_75t_R g1071 ( 
.A(n_936),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_945),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1014),
.B(n_1033),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_957),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1030),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_933),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_L g1077 ( 
.A(n_1024),
.B(n_906),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_933),
.Y(n_1078)
);

CKINVDCx11_ASAP7_75t_R g1079 ( 
.A(n_973),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_963),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_SL g1081 ( 
.A(n_1001),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_970),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_933),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_975),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_982),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_934),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_982),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_1005),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_981),
.Y(n_1089)
);

OAI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_994),
.A2(n_913),
.B1(n_884),
.B2(n_617),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_934),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_948),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_988),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_993),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1005),
.B(n_640),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_948),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_948),
.Y(n_1097)
);

BUFx10_ASAP7_75t_L g1098 ( 
.A(n_1005),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_1017),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_999),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_972),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1010),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1015),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_948),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1033),
.B(n_1034),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_960),
.Y(n_1106)
);

NOR2x1p5_ASAP7_75t_L g1107 ( 
.A(n_1017),
.B(n_623),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1006),
.B(n_647),
.Y(n_1108)
);

AND3x2_ASAP7_75t_L g1109 ( 
.A(n_952),
.B(n_889),
.C(n_796),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1018),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1020),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1021),
.Y(n_1112)
);

NOR2x1p5_ASAP7_75t_L g1113 ( 
.A(n_931),
.B(n_626),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_956),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_960),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1034),
.B(n_626),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_960),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_956),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1027),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1031),
.Y(n_1120)
);

CKINVDCx8_ASAP7_75t_R g1121 ( 
.A(n_1002),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_966),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_973),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1006),
.B(n_632),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_953),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_966),
.Y(n_1126)
);

AO22x2_ASAP7_75t_L g1127 ( 
.A1(n_983),
.A2(n_918),
.B1(n_621),
.B2(n_663),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_953),
.Y(n_1128)
);

AND2x2_ASAP7_75t_SL g1129 ( 
.A(n_935),
.B(n_615),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_962),
.B(n_822),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1028),
.A2(n_632),
.B1(n_642),
.B2(n_635),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1029),
.B(n_906),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_977),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1016),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_978),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_962),
.B(n_1011),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_977),
.Y(n_1137)
);

AND3x2_ASAP7_75t_L g1138 ( 
.A(n_1011),
.B(n_663),
.C(n_621),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_979),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_978),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_947),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_979),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_979),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_979),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1032),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1032),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_995),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_995),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_955),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1029),
.B(n_906),
.Y(n_1150)
);

INVx8_ASAP7_75t_L g1151 ( 
.A(n_1029),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_1029),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1028),
.B(n_635),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_949),
.B(n_822),
.Y(n_1154)
);

INVx8_ASAP7_75t_L g1155 ( 
.A(n_1006),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_961),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_955),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_995),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_969),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_959),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_949),
.B(n_1012),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_959),
.Y(n_1162)
);

AND3x2_ASAP7_75t_L g1163 ( 
.A(n_930),
.B(n_715),
.C(n_681),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_996),
.Y(n_1164)
);

INVx5_ASAP7_75t_L g1165 ( 
.A(n_996),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_974),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_996),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_984),
.B(n_642),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_996),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_998),
.Y(n_1170)
);

INVxp33_ASAP7_75t_SL g1171 ( 
.A(n_974),
.Y(n_1171)
);

NOR2x1p5_ASAP7_75t_L g1172 ( 
.A(n_980),
.B(n_643),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_976),
.B(n_643),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_998),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_969),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_998),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_987),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_954),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_976),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1003),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1003),
.B(n_645),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1004),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1004),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_987),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1022),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_969),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1009),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1022),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_954),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1000),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_989),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1022),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1022),
.B(n_906),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1025),
.B(n_719),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_SL g1195 ( 
.A(n_1025),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1025),
.B(n_726),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_964),
.B(n_732),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1019),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1019),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1000),
.B(n_761),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_997),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1014),
.B(n_693),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1013),
.B(n_804),
.Y(n_1203)
);

BUFx10_ASAP7_75t_L g1204 ( 
.A(n_942),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_943),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1114),
.B(n_1118),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1160),
.A2(n_667),
.B1(n_894),
.B2(n_591),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1069),
.B(n_625),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1072),
.B(n_625),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1145),
.B(n_628),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1041),
.Y(n_1211)
);

OAI21xp33_ASAP7_75t_L g1212 ( 
.A1(n_1162),
.A2(n_600),
.B(n_598),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1146),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1135),
.B(n_628),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1140),
.B(n_634),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1040),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1125),
.B(n_634),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1199),
.A2(n_823),
.B(n_818),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1161),
.B(n_644),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1058),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1128),
.B(n_644),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1149),
.B(n_878),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_L g1223 ( 
.A(n_1131),
.B(n_878),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1171),
.B(n_678),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1157),
.B(n_832),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1043),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1085),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1044),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1045),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1166),
.A2(n_610),
.B(n_611),
.C(n_603),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1050),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1059),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1179),
.B(n_680),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1171),
.B(n_1153),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1134),
.B(n_682),
.Y(n_1235)
);

NOR3xp33_ASAP7_75t_L g1236 ( 
.A(n_1090),
.B(n_639),
.C(n_627),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1134),
.B(n_690),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1057),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1054),
.B(n_664),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1180),
.B(n_699),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1116),
.B(n_700),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1065),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1074),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1154),
.B(n_704),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1085),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1095),
.B(n_705),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1095),
.B(n_706),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1055),
.B(n_694),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1036),
.B(n_710),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1080),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1082),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1108),
.B(n_1130),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1084),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1089),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1108),
.B(n_711),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1093),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1094),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1136),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1203),
.A2(n_614),
.B1(n_620),
.B2(n_612),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1064),
.B(n_738),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1100),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_SL g1262 ( 
.A(n_1066),
.B(n_894),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_SL g1263 ( 
.A(n_1129),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1060),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1063),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1068),
.B(n_752),
.Y(n_1266)
);

NAND3xp33_ASAP7_75t_L g1267 ( 
.A(n_1173),
.B(n_760),
.C(n_693),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1070),
.B(n_1088),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1071),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1039),
.B(n_754),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1102),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1068),
.B(n_784),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1087),
.B(n_629),
.Y(n_1273)
);

OR2x6_ASAP7_75t_L g1274 ( 
.A(n_1155),
.B(n_1127),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1087),
.B(n_788),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1066),
.A2(n_667),
.B1(n_763),
.B2(n_760),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1124),
.B(n_759),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1101),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1099),
.B(n_800),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1099),
.B(n_1168),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1181),
.B(n_834),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1105),
.B(n_837),
.Y(n_1282)
);

OAI21xp33_ASAP7_75t_L g1283 ( 
.A1(n_1129),
.A2(n_637),
.B(n_630),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1098),
.B(n_846),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1103),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1048),
.B(n_856),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1110),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1049),
.B(n_1203),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1111),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1107),
.B(n_646),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1112),
.B(n_875),
.Y(n_1291)
);

AO221x1_ASAP7_75t_L g1292 ( 
.A1(n_1090),
.A2(n_638),
.B1(n_653),
.B2(n_617),
.C(n_607),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1119),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1151),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1035),
.B(n_862),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1151),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_SL g1297 ( 
.A(n_1204),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1051),
.B(n_922),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1202),
.B(n_763),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1155),
.B(n_879),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1151),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1073),
.B(n_870),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1120),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1193),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1194),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1062),
.B(n_919),
.Y(n_1306)
);

BUFx5_ASAP7_75t_L g1307 ( 
.A(n_1192),
.Y(n_1307)
);

NOR2xp67_ASAP7_75t_L g1308 ( 
.A(n_1141),
.B(n_873),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1062),
.B(n_873),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1113),
.B(n_874),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1138),
.B(n_874),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1079),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1197),
.B(n_887),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1138),
.B(n_876),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1197),
.B(n_877),
.C(n_876),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1077),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1077),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1081),
.B(n_720),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1132),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1109),
.Y(n_1320)
);

AO221x1_ASAP7_75t_L g1321 ( 
.A1(n_1127),
.A2(n_653),
.B1(n_654),
.B2(n_638),
.C(n_607),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1132),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1189),
.B(n_822),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1187),
.B(n_877),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1205),
.B(n_880),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1205),
.B(n_880),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1037),
.B(n_885),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1109),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1150),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1123),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1038),
.B(n_1042),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1042),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1150),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1156),
.B(n_593),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1047),
.Y(n_1335)
);

OR2x6_ASAP7_75t_L g1336 ( 
.A(n_1127),
.B(n_633),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1052),
.B(n_886),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1156),
.B(n_599),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1163),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1053),
.B(n_891),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1200),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1177),
.B(n_601),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1056),
.B(n_1061),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1172),
.B(n_899),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1056),
.B(n_681),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_R g1346 ( 
.A(n_1046),
.B(n_654),
.Y(n_1346)
);

AO221x1_ASAP7_75t_L g1347 ( 
.A1(n_1163),
.A2(n_691),
.B1(n_717),
.B2(n_684),
.C(n_668),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1067),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1075),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1075),
.B(n_715),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1195),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1178),
.A2(n_684),
.B1(n_691),
.B2(n_668),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1196),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1178),
.B(n_602),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1198),
.B(n_718),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1190),
.B(n_605),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1184),
.B(n_718),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1191),
.B(n_745),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1201),
.B(n_857),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1152),
.B(n_745),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1152),
.Y(n_1361)
);

NOR3xp33_ASAP7_75t_L g1362 ( 
.A(n_1079),
.B(n_785),
.C(n_751),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1165),
.B(n_921),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1195),
.B(n_609),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1121),
.B(n_651),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1165),
.B(n_767),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1165),
.Y(n_1367)
);

BUFx8_ASAP7_75t_L g1368 ( 
.A(n_1159),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1122),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1122),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1076),
.B(n_767),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_SL g1372 ( 
.A(n_1159),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1159),
.B(n_658),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1175),
.B(n_660),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1126),
.A2(n_650),
.B1(n_656),
.B2(n_652),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1188),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1133),
.B(n_666),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1175),
.B(n_669),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1137),
.A2(n_742),
.B1(n_756),
.B2(n_717),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1137),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1186),
.B(n_672),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1139),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1139),
.Y(n_1383)
);

NOR2xp67_ASAP7_75t_L g1384 ( 
.A(n_1142),
.B(n_23),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1143),
.Y(n_1385)
);

NAND3xp33_ASAP7_75t_L g1386 ( 
.A(n_1144),
.B(n_676),
.C(n_673),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1144),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1147),
.B(n_721),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1186),
.B(n_679),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1148),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_SL g1391 ( 
.A(n_1188),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1148),
.B(n_712),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1076),
.B(n_791),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1188),
.Y(n_1394)
);

AND2x2_ASAP7_75t_SL g1395 ( 
.A(n_1158),
.B(n_816),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1164),
.B(n_687),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1167),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1169),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1078),
.B(n_871),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1169),
.B(n_698),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1170),
.B(n_702),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1170),
.A2(n_756),
.B1(n_757),
.B2(n_742),
.Y(n_1402)
);

NAND2xp33_ASAP7_75t_SL g1403 ( 
.A(n_1188),
.B(n_757),
.Y(n_1403)
);

NOR3xp33_ASAP7_75t_L g1404 ( 
.A(n_1174),
.B(n_865),
.C(n_825),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1083),
.B(n_897),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1185),
.B(n_24),
.Y(n_1406)
);

BUFx5_ASAP7_75t_L g1407 ( 
.A(n_1086),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1176),
.B(n_707),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1234),
.B(n_780),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1206),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1213),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1206),
.B(n_709),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1216),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1208),
.B(n_1209),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1226),
.Y(n_1415)
);

NOR2xp67_ASAP7_75t_L g1416 ( 
.A(n_1264),
.B(n_21),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1296),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1208),
.B(n_714),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1211),
.B(n_780),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1232),
.B(n_797),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1228),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1209),
.B(n_1210),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1359),
.A2(n_1092),
.B(n_1091),
.Y(n_1423)
);

BUFx4f_ASAP7_75t_L g1424 ( 
.A(n_1339),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1229),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1355),
.A2(n_1096),
.B(n_1092),
.Y(n_1426)
);

BUFx12f_ASAP7_75t_L g1427 ( 
.A(n_1312),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1296),
.B(n_724),
.Y(n_1428)
);

O2A1O1Ixp5_ASAP7_75t_L g1429 ( 
.A1(n_1306),
.A2(n_924),
.B(n_927),
.C(n_910),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1231),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1355),
.A2(n_1104),
.B(n_1097),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1334),
.A2(n_1342),
.B(n_1338),
.C(n_1238),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1210),
.B(n_725),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1288),
.A2(n_1317),
.B(n_1316),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1296),
.B(n_729),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1252),
.B(n_731),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1357),
.A2(n_1106),
.B(n_1104),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1222),
.B(n_735),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1368),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1220),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1258),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1273),
.B(n_737),
.Y(n_1442)
);

OAI21xp33_ASAP7_75t_L g1443 ( 
.A1(n_1258),
.A2(n_925),
.B(n_923),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1368),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1222),
.B(n_1217),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1352),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1358),
.A2(n_1117),
.B(n_1115),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1225),
.A2(n_1183),
.B(n_1182),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1273),
.B(n_739),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1242),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1403),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1243),
.A2(n_671),
.B(n_685),
.C(n_677),
.Y(n_1452)
);

CKINVDCx6p67_ASAP7_75t_R g1453 ( 
.A(n_1265),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1230),
.A2(n_686),
.B(n_695),
.C(n_689),
.Y(n_1454)
);

INVx4_ASAP7_75t_L g1455 ( 
.A(n_1297),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1269),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1280),
.B(n_741),
.Y(n_1457)
);

BUFx4f_ASAP7_75t_L g1458 ( 
.A(n_1274),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1250),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1221),
.B(n_744),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1324),
.B(n_797),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1341),
.B(n_696),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1251),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1219),
.B(n_746),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1354),
.B(n_805),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1225),
.A2(n_1185),
.B(n_1183),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1253),
.B(n_749),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1343),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1254),
.B(n_750),
.Y(n_1469)
);

OAI21xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1257),
.A2(n_701),
.B(n_697),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1331),
.A2(n_708),
.B(n_703),
.Y(n_1471)
);

OAI321xp33_ASAP7_75t_L g1472 ( 
.A1(n_1336),
.A2(n_730),
.A3(n_716),
.B1(n_734),
.B2(n_727),
.C(n_713),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1286),
.A2(n_747),
.B(n_743),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1261),
.B(n_753),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1285),
.B(n_755),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1207),
.B(n_805),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1287),
.B(n_758),
.Y(n_1477)
);

NAND2x1p5_ASAP7_75t_L g1478 ( 
.A(n_1351),
.B(n_927),
.Y(n_1478)
);

INVx11_ASAP7_75t_L g1479 ( 
.A(n_1278),
.Y(n_1479)
);

OAI321xp33_ASAP7_75t_L g1480 ( 
.A1(n_1336),
.A2(n_781),
.A3(n_764),
.B1(n_782),
.B2(n_774),
.C(n_770),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1289),
.B(n_1212),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1256),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1244),
.B(n_762),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1227),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1259),
.B(n_765),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1283),
.A2(n_792),
.B(n_795),
.C(n_789),
.Y(n_1486)
);

AND2x6_ASAP7_75t_L g1487 ( 
.A(n_1351),
.B(n_812),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1356),
.B(n_809),
.Y(n_1488)
);

BUFx4f_ASAP7_75t_L g1489 ( 
.A(n_1274),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1218),
.A2(n_829),
.B(n_828),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1271),
.Y(n_1491)
);

INVxp67_ASAP7_75t_SL g1492 ( 
.A(n_1402),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1218),
.A2(n_835),
.B(n_831),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1233),
.A2(n_839),
.B(n_836),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1305),
.A2(n_849),
.B(n_847),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1377),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1315),
.A2(n_853),
.B(n_852),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1313),
.A2(n_860),
.B(n_855),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1240),
.A2(n_869),
.B(n_866),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1377),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1352),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1236),
.A2(n_882),
.B(n_883),
.C(n_872),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1290),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1346),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1263),
.A2(n_1323),
.B1(n_1344),
.B2(n_1223),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1239),
.B(n_1404),
.C(n_1267),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1263),
.A2(n_768),
.B1(n_771),
.B2(n_766),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1241),
.B(n_772),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1297),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1309),
.A2(n_821),
.B1(n_838),
.B2(n_810),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1408),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1325),
.B(n_776),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1245),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1293),
.B(n_888),
.Y(n_1514)
);

OAI321xp33_ASAP7_75t_L g1515 ( 
.A1(n_1336),
.A2(n_900),
.A3(n_895),
.B1(n_902),
.B2(n_896),
.C(n_890),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1319),
.A2(n_909),
.B(n_904),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1322),
.A2(n_915),
.B(n_912),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1294),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1329),
.A2(n_778),
.B(n_777),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1299),
.B(n_779),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1332),
.A2(n_898),
.B(n_786),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1326),
.B(n_783),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1333),
.A2(n_793),
.B(n_787),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1301),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1376),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1327),
.B(n_794),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1379),
.B(n_798),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1214),
.A2(n_801),
.B(n_799),
.Y(n_1528)
);

INVxp33_ASAP7_75t_SL g1529 ( 
.A(n_1262),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1215),
.A2(n_803),
.B(n_802),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1304),
.A2(n_807),
.B(n_806),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1262),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1345),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1337),
.B(n_811),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1320),
.B(n_814),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1340),
.B(n_815),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1302),
.B(n_817),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1335),
.A2(n_824),
.B(n_820),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1290),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1274),
.B(n_810),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1277),
.B(n_827),
.Y(n_1541)
);

INVx6_ASAP7_75t_L g1542 ( 
.A(n_1392),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1291),
.B(n_833),
.Y(n_1543)
);

BUFx4f_ASAP7_75t_L g1544 ( 
.A(n_1328),
.Y(n_1544)
);

O2A1O1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1310),
.A2(n_838),
.B(n_868),
.C(n_821),
.Y(n_1545)
);

AOI21xp33_ASAP7_75t_L g1546 ( 
.A1(n_1318),
.A2(n_842),
.B(n_840),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1291),
.B(n_843),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1330),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1345),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1303),
.B(n_844),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1376),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1284),
.B(n_848),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1276),
.A2(n_851),
.B1(n_858),
.B2(n_850),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1350),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1395),
.A2(n_1282),
.B1(n_1246),
.B2(n_1255),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1350),
.Y(n_1556)
);

INVx4_ASAP7_75t_L g1557 ( 
.A(n_1391),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1292),
.B(n_868),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1376),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1348),
.A2(n_863),
.B(n_861),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1353),
.A2(n_905),
.B(n_901),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1224),
.B(n_911),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1364),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1247),
.B(n_916),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1321),
.B(n_892),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1349),
.A2(n_920),
.B(n_917),
.Y(n_1566)
);

BUFx4f_ASAP7_75t_L g1567 ( 
.A(n_1392),
.Y(n_1567)
);

O2A1O1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1311),
.A2(n_1314),
.B(n_1281),
.C(n_1270),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1249),
.A2(n_892),
.B(n_926),
.C(n_28),
.Y(n_1569)
);

AOI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1295),
.A2(n_580),
.B(n_578),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1260),
.B(n_25),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1300),
.A2(n_28),
.B(n_25),
.C(n_26),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1266),
.B(n_29),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1272),
.B(n_29),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1391),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1275),
.A2(n_1279),
.B(n_1298),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1347),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1366),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1366),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1360),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1371),
.A2(n_520),
.B(n_519),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1392),
.Y(n_1582)
);

NAND2x1p5_ASAP7_75t_L g1583 ( 
.A(n_1235),
.B(n_30),
.Y(n_1583)
);

CKINVDCx10_ASAP7_75t_R g1584 ( 
.A(n_1362),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1375),
.B(n_32),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1248),
.B(n_33),
.Y(n_1586)
);

NOR2x1_ASAP7_75t_L g1587 ( 
.A(n_1308),
.B(n_34),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1268),
.B(n_34),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1237),
.B(n_35),
.Y(n_1589)
);

BUFx8_ASAP7_75t_SL g1590 ( 
.A(n_1361),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1386),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1367),
.B(n_40),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1365),
.B(n_41),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1373),
.B(n_42),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1394),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1396),
.B(n_43),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1374),
.Y(n_1597)
);

OAI321xp33_ASAP7_75t_L g1598 ( 
.A1(n_1371),
.A2(n_47),
.A3(n_49),
.B1(n_44),
.B2(n_45),
.C(n_48),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1400),
.B(n_44),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1378),
.B(n_45),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1401),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1393),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_SL g1603 ( 
.A(n_1372),
.B(n_531),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1393),
.Y(n_1604)
);

OAI22x1_ASAP7_75t_L g1605 ( 
.A1(n_1363),
.A2(n_53),
.B1(n_50),
.B2(n_51),
.Y(n_1605)
);

BUFx2_ASAP7_75t_SL g1606 ( 
.A(n_1384),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1381),
.B(n_53),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1389),
.B(n_54),
.Y(n_1608)
);

NAND2xp33_ASAP7_75t_L g1609 ( 
.A(n_1307),
.B(n_535),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1399),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1405),
.B(n_55),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1388),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1406),
.Y(n_1613)
);

AOI21xp33_ASAP7_75t_L g1614 ( 
.A1(n_1388),
.A2(n_60),
.B(n_61),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1369),
.A2(n_538),
.B(n_537),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1307),
.B(n_61),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1407),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1307),
.B(n_63),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1407),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1380),
.Y(n_1620)
);

BUFx4f_ASAP7_75t_L g1621 ( 
.A(n_1394),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1383),
.Y(n_1622)
);

NOR2x2_ASAP7_75t_L g1623 ( 
.A(n_1370),
.B(n_65),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1307),
.A2(n_69),
.B1(n_66),
.B2(n_67),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1407),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1407),
.A2(n_71),
.B1(n_67),
.B2(n_70),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1387),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1390),
.A2(n_1398),
.B(n_1397),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1394),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1382),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1385),
.B(n_75),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1206),
.B(n_76),
.Y(n_1632)
);

NOR2xp67_ASAP7_75t_L g1633 ( 
.A(n_1264),
.B(n_77),
.Y(n_1633)
);

A2O1A1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1213),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1206),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1206),
.B(n_81),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1206),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1206),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1206),
.B(n_82),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1206),
.B(n_83),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1234),
.B(n_83),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1206),
.B(n_84),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1206),
.B(n_84),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1206),
.B(n_85),
.Y(n_1644)
);

OR2x2_ASAP7_75t_SL g1645 ( 
.A(n_1278),
.B(n_85),
.Y(n_1645)
);

BUFx10_ASAP7_75t_L g1646 ( 
.A(n_1297),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1206),
.A2(n_91),
.B1(n_86),
.B2(n_90),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1234),
.B(n_90),
.Y(n_1648)
);

BUFx12f_ASAP7_75t_L g1649 ( 
.A(n_1312),
.Y(n_1649)
);

O2A1O1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1232),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1206),
.B(n_92),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1637),
.B(n_93),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1410),
.B(n_95),
.Y(n_1653)
);

AOI221x1_ASAP7_75t_L g1654 ( 
.A1(n_1432),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.C(n_103),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1410),
.B(n_98),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1635),
.B(n_99),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1638),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1441),
.B(n_100),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1446),
.B(n_103),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1411),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1413),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1548),
.Y(n_1662)
);

AOI21xp33_ASAP7_75t_L g1663 ( 
.A1(n_1608),
.A2(n_104),
.B(n_105),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_SL g1664 ( 
.A(n_1529),
.B(n_105),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1501),
.B(n_106),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1468),
.B(n_107),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1414),
.A2(n_1422),
.B(n_1445),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1502),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.C(n_111),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1453),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1503),
.B(n_112),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1533),
.B(n_112),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1549),
.B(n_113),
.Y(n_1672)
);

OAI22x1_ASAP7_75t_L g1673 ( 
.A1(n_1540),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1554),
.B(n_114),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1439),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1557),
.B(n_117),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1415),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1419),
.B(n_117),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1421),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1632),
.A2(n_1636),
.B1(n_1644),
.B2(n_1639),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1557),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1556),
.B(n_118),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1425),
.B(n_1430),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1450),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1461),
.B(n_121),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1490),
.A2(n_122),
.B(n_123),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1439),
.B(n_124),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1459),
.Y(n_1688)
);

BUFx4_ASAP7_75t_SL g1689 ( 
.A(n_1504),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_SL g1690 ( 
.A1(n_1615),
.A2(n_126),
.B(n_127),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1424),
.B(n_130),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1629),
.A2(n_130),
.B(n_132),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1465),
.B(n_133),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1409),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1625),
.A2(n_137),
.B(n_138),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1420),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1476),
.B(n_137),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1625),
.A2(n_138),
.B(n_139),
.Y(n_1698)
);

AO21x2_ASAP7_75t_L g1699 ( 
.A1(n_1490),
.A2(n_139),
.B(n_140),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1463),
.B(n_1492),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1426),
.A2(n_140),
.B(n_141),
.Y(n_1701)
);

AO31x2_ASAP7_75t_L g1702 ( 
.A1(n_1616),
.A2(n_144),
.A3(n_142),
.B(n_143),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1651),
.A2(n_148),
.B1(n_145),
.B2(n_147),
.Y(n_1703)
);

INVx3_ASAP7_75t_SL g1704 ( 
.A(n_1646),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1494),
.A2(n_150),
.B(n_145),
.C(n_149),
.Y(n_1705)
);

OAI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1493),
.A2(n_150),
.B(n_151),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1479),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1434),
.B(n_151),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1434),
.B(n_152),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1482),
.Y(n_1710)
);

AO31x2_ASAP7_75t_L g1711 ( 
.A1(n_1618),
.A2(n_1486),
.A3(n_1555),
.B(n_1605),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1424),
.B(n_154),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1623),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1491),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1431),
.A2(n_154),
.B(n_155),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1444),
.B(n_156),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1578),
.Y(n_1717)
);

OAI22x1_ASAP7_75t_L g1718 ( 
.A1(n_1540),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1602),
.A2(n_1604),
.B(n_1580),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1506),
.B(n_161),
.C(n_162),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1525),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1444),
.B(n_164),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1499),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_1723)
);

BUFx12f_ASAP7_75t_L g1724 ( 
.A(n_1646),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1544),
.B(n_167),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1496),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1437),
.A2(n_168),
.B(n_169),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_L g1728 ( 
.A(n_1525),
.B(n_170),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1454),
.A2(n_174),
.B1(n_171),
.B2(n_173),
.C(n_175),
.Y(n_1729)
);

INVx4_ASAP7_75t_L g1730 ( 
.A(n_1458),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1500),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1601),
.B(n_173),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1458),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1488),
.B(n_179),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1427),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1544),
.B(n_182),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1514),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1576),
.A2(n_183),
.B(n_184),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1510),
.Y(n_1739)
);

INVx4_ASAP7_75t_L g1740 ( 
.A(n_1489),
.Y(n_1740)
);

INVx2_ASAP7_75t_SL g1741 ( 
.A(n_1455),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1579),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1489),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1628),
.A2(n_186),
.B(n_187),
.Y(n_1744)
);

BUFx10_ASAP7_75t_L g1745 ( 
.A(n_1487),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1481),
.A2(n_187),
.B(n_188),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1473),
.B(n_188),
.Y(n_1747)
);

INVx4_ASAP7_75t_SL g1748 ( 
.A(n_1487),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1447),
.A2(n_193),
.B(n_194),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1448),
.A2(n_193),
.B(n_194),
.Y(n_1750)
);

OR2x6_ASAP7_75t_L g1751 ( 
.A(n_1455),
.B(n_1456),
.Y(n_1751)
);

NAND3xp33_ASAP7_75t_SL g1752 ( 
.A(n_1577),
.B(n_195),
.C(n_196),
.Y(n_1752)
);

AO21x1_ASAP7_75t_L g1753 ( 
.A1(n_1581),
.A2(n_196),
.B(n_197),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1641),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_1754)
);

AOI21xp33_ASAP7_75t_L g1755 ( 
.A1(n_1586),
.A2(n_199),
.B(n_200),
.Y(n_1755)
);

NAND2x1_ASAP7_75t_L g1756 ( 
.A(n_1551),
.B(n_200),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1509),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1514),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1649),
.Y(n_1759)
);

NAND2x1_ASAP7_75t_L g1760 ( 
.A(n_1559),
.B(n_202),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1487),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1539),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_SL g1763 ( 
.A1(n_1581),
.A2(n_203),
.B(n_204),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1610),
.Y(n_1764)
);

AOI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1611),
.A2(n_205),
.B(n_206),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1412),
.B(n_205),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_1532),
.B(n_208),
.C(n_209),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1563),
.B(n_208),
.Y(n_1768)
);

NOR2xp67_ASAP7_75t_L g1769 ( 
.A(n_1472),
.B(n_209),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1466),
.A2(n_210),
.B(n_211),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1620),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1596),
.A2(n_210),
.B(n_211),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1511),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1511),
.B(n_212),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1599),
.A2(n_212),
.B(n_213),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1590),
.Y(n_1776)
);

AOI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1470),
.A2(n_216),
.B1(n_213),
.B2(n_215),
.C(n_217),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1624),
.A2(n_218),
.B1(n_215),
.B2(n_216),
.Y(n_1778)
);

INVx3_ASAP7_75t_SL g1779 ( 
.A(n_1645),
.Y(n_1779)
);

AOI22x1_ASAP7_75t_L g1780 ( 
.A1(n_1570),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1460),
.A2(n_223),
.B(n_224),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1418),
.A2(n_225),
.B(n_226),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1622),
.Y(n_1783)
);

BUFx8_ASAP7_75t_SL g1784 ( 
.A(n_1567),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1495),
.B(n_229),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1433),
.A2(n_230),
.B(n_231),
.Y(n_1786)
);

CKINVDCx20_ASAP7_75t_R g1787 ( 
.A(n_1567),
.Y(n_1787)
);

OAI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1516),
.A2(n_232),
.B(n_233),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1527),
.B(n_239),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1438),
.A2(n_240),
.B(n_241),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1442),
.B(n_243),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1521),
.B(n_244),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1495),
.B(n_245),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1462),
.B(n_246),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1462),
.B(n_247),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1558),
.A2(n_1565),
.B1(n_1648),
.B2(n_1607),
.Y(n_1796)
);

NAND2x1p5_ASAP7_75t_L g1797 ( 
.A(n_1575),
.B(n_249),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1627),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1630),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1517),
.A2(n_250),
.B(n_251),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1640),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_SL g1802 ( 
.A1(n_1452),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.C(n_255),
.Y(n_1802)
);

AND3x4_ASAP7_75t_L g1803 ( 
.A(n_1584),
.B(n_252),
.C(n_256),
.Y(n_1803)
);

NAND2x1p5_ASAP7_75t_L g1804 ( 
.A(n_1575),
.B(n_256),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1487),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1423),
.A2(n_257),
.B(n_259),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1497),
.B(n_261),
.Y(n_1807)
);

OA22x2_ASAP7_75t_L g1808 ( 
.A1(n_1505),
.A2(n_265),
.B1(n_262),
.B2(n_264),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1521),
.B(n_262),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1571),
.A2(n_265),
.B(n_267),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1478),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1573),
.A2(n_267),
.B(n_268),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1449),
.B(n_1535),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1478),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1574),
.A2(n_269),
.B(n_270),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1621),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1595),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1609),
.A2(n_269),
.B(n_271),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1543),
.A2(n_271),
.B(n_272),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1642),
.Y(n_1820)
);

AO21x1_ASAP7_75t_L g1821 ( 
.A1(n_1643),
.A2(n_273),
.B(n_274),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1595),
.Y(n_1822)
);

AO21x1_ASAP7_75t_L g1823 ( 
.A1(n_1631),
.A2(n_278),
.B(n_279),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1542),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1592),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1607),
.A2(n_286),
.B1(n_283),
.B2(n_285),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1429),
.A2(n_287),
.B(n_288),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1440),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1498),
.B(n_289),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1585),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1498),
.B(n_292),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1547),
.B(n_293),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1595),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1512),
.A2(n_293),
.B(n_294),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1518),
.B(n_1524),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1436),
.B(n_294),
.Y(n_1836)
);

OAI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1471),
.A2(n_295),
.B(n_296),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1560),
.B(n_296),
.Y(n_1838)
);

NOR2x1_ASAP7_75t_SL g1839 ( 
.A(n_1606),
.B(n_297),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1417),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1417),
.Y(n_1841)
);

INVx1_ASAP7_75t_SL g1842 ( 
.A(n_1542),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1560),
.B(n_300),
.Y(n_1843)
);

AND3x4_ASAP7_75t_L g1844 ( 
.A(n_1587),
.B(n_301),
.C(n_302),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1566),
.B(n_303),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1428),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1568),
.A2(n_303),
.B(n_305),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1518),
.B(n_306),
.Y(n_1848)
);

OAI21x1_ASAP7_75t_L g1849 ( 
.A1(n_1613),
.A2(n_306),
.B(n_307),
.Y(n_1849)
);

OAI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1467),
.A2(n_1474),
.B(n_1469),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1553),
.B(n_307),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1537),
.A2(n_308),
.B(n_309),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1566),
.B(n_1538),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1451),
.A2(n_1612),
.B1(n_1634),
.B2(n_1633),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1483),
.B(n_1562),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1475),
.Y(n_1856)
);

BUFx8_ASAP7_75t_L g1857 ( 
.A(n_1582),
.Y(n_1857)
);

A2O1A1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1572),
.A2(n_311),
.B(n_312),
.C(n_313),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1484),
.A2(n_315),
.B(n_316),
.Y(n_1859)
);

OAI21x1_ASAP7_75t_L g1860 ( 
.A1(n_1513),
.A2(n_315),
.B(n_316),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1477),
.Y(n_1861)
);

OAI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1561),
.A2(n_318),
.B(n_319),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1435),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1522),
.B(n_1526),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1534),
.A2(n_319),
.B(n_320),
.Y(n_1865)
);

BUFx5_ASAP7_75t_L g1866 ( 
.A(n_1621),
.Y(n_1866)
);

OAI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1519),
.A2(n_322),
.B(n_323),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1451),
.Y(n_1868)
);

OAI21x1_ASAP7_75t_L g1869 ( 
.A1(n_1524),
.A2(n_322),
.B(n_324),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1523),
.A2(n_324),
.B(n_325),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1536),
.A2(n_326),
.B(n_327),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1588),
.B(n_326),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1619),
.Y(n_1873)
);

OA21x2_ASAP7_75t_L g1874 ( 
.A1(n_1598),
.A2(n_328),
.B(n_329),
.Y(n_1874)
);

NAND3xp33_ASAP7_75t_SL g1875 ( 
.A(n_1650),
.B(n_1569),
.C(n_1545),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1583),
.Y(n_1876)
);

AOI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1443),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1564),
.B(n_335),
.Y(n_1878)
);

OAI21x1_ASAP7_75t_L g1879 ( 
.A1(n_1583),
.A2(n_336),
.B(n_337),
.Y(n_1879)
);

BUFx4f_ASAP7_75t_L g1880 ( 
.A(n_1594),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1597),
.Y(n_1881)
);

AOI21x1_ASAP7_75t_L g1882 ( 
.A1(n_1600),
.A2(n_336),
.B(n_338),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1541),
.B(n_339),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1589),
.B(n_339),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1507),
.B(n_340),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1593),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1485),
.B(n_341),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1531),
.A2(n_344),
.B(n_345),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1546),
.B(n_344),
.Y(n_1889)
);

AOI221x1_ASAP7_75t_L g1890 ( 
.A1(n_1591),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.C(n_349),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1550),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1617),
.Y(n_1892)
);

INVx3_ASAP7_75t_L g1893 ( 
.A(n_1603),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1520),
.B(n_348),
.Y(n_1894)
);

AND3x4_ASAP7_75t_L g1895 ( 
.A(n_1416),
.B(n_350),
.C(n_352),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1464),
.A2(n_352),
.B(n_353),
.Y(n_1896)
);

OAI21xp33_ASAP7_75t_SL g1897 ( 
.A1(n_1614),
.A2(n_353),
.B(n_354),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1508),
.B(n_355),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1457),
.B(n_355),
.Y(n_1899)
);

A2O1A1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1472),
.A2(n_356),
.B(n_357),
.C(n_358),
.Y(n_1900)
);

OAI21x1_ASAP7_75t_L g1901 ( 
.A1(n_1647),
.A2(n_356),
.B(n_357),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1552),
.B(n_358),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_SL g1903 ( 
.A1(n_1480),
.A2(n_359),
.B(n_360),
.Y(n_1903)
);

OAI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1528),
.A2(n_361),
.B(n_362),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1530),
.A2(n_361),
.B(n_363),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1480),
.A2(n_364),
.B(n_365),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1515),
.B(n_365),
.Y(n_1907)
);

NAND2x1p5_ASAP7_75t_L g1908 ( 
.A(n_1515),
.B(n_366),
.Y(n_1908)
);

OR2x6_ASAP7_75t_L g1909 ( 
.A(n_1626),
.B(n_501),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1410),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1410),
.B(n_367),
.Y(n_1911)
);

AO21x2_ASAP7_75t_L g1912 ( 
.A1(n_1490),
.A2(n_370),
.B(n_371),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1414),
.A2(n_373),
.B(n_375),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1479),
.Y(n_1914)
);

AOI21xp33_ASAP7_75t_L g1915 ( 
.A1(n_1608),
.A2(n_375),
.B(n_376),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1410),
.B(n_377),
.Y(n_1916)
);

NAND2x1p5_ASAP7_75t_L g1917 ( 
.A(n_1410),
.B(n_378),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1410),
.B(n_378),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1432),
.A2(n_379),
.B(n_381),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1637),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1637),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1410),
.B(n_379),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1410),
.B(n_382),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1432),
.A2(n_383),
.B(n_384),
.Y(n_1924)
);

AOI21xp33_ASAP7_75t_L g1925 ( 
.A1(n_1608),
.A2(n_386),
.B(n_387),
.Y(n_1925)
);

AOI221xp5_ASAP7_75t_L g1926 ( 
.A1(n_1446),
.A2(n_386),
.B1(n_388),
.B2(n_389),
.C(n_390),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1432),
.A2(n_388),
.B(n_389),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1410),
.B(n_392),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1410),
.B(n_393),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1432),
.A2(n_393),
.B(n_394),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1446),
.B(n_395),
.Y(n_1931)
);

NOR2x1_ASAP7_75t_L g1932 ( 
.A(n_1455),
.B(n_396),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1432),
.A2(n_397),
.B(n_398),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1410),
.B(n_397),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1432),
.A2(n_399),
.B(n_401),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1637),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1432),
.A2(n_403),
.B(n_404),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1410),
.B(n_403),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1637),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1410),
.A2(n_404),
.B1(n_406),
.B2(n_407),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1637),
.B(n_408),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1637),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1637),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_SL g1944 ( 
.A1(n_1635),
.A2(n_410),
.B(n_411),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1414),
.A2(n_411),
.B(n_412),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1410),
.B(n_413),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1414),
.A2(n_413),
.B(n_414),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1525),
.Y(n_1948)
);

INVx4_ASAP7_75t_L g1949 ( 
.A(n_1439),
.Y(n_1949)
);

AOI21xp33_ASAP7_75t_L g1950 ( 
.A1(n_1608),
.A2(n_416),
.B(n_417),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1635),
.Y(n_1951)
);

OR2x6_ASAP7_75t_L g1952 ( 
.A(n_1637),
.B(n_501),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1646),
.Y(n_1953)
);

A2O1A1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1635),
.A2(n_418),
.B(n_419),
.C(n_420),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1502),
.A2(n_418),
.B1(n_420),
.B2(n_422),
.C(n_424),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1479),
.Y(n_1956)
);

NAND2x1p5_ASAP7_75t_L g1957 ( 
.A(n_1410),
.B(n_425),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1525),
.Y(n_1958)
);

OAI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1432),
.A2(n_427),
.B(n_428),
.Y(n_1959)
);

OAI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1432),
.A2(n_427),
.B(n_431),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1637),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1637),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1410),
.B(n_432),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1637),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1637),
.B(n_433),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1410),
.B(n_433),
.Y(n_1966)
);

O2A1O1Ixp5_ASAP7_75t_L g1967 ( 
.A1(n_1432),
.A2(n_434),
.B(n_435),
.C(n_436),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1432),
.A2(n_434),
.B(n_435),
.Y(n_1968)
);

NAND2x1p5_ASAP7_75t_L g1969 ( 
.A(n_1410),
.B(n_437),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1637),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1410),
.A2(n_439),
.B1(n_441),
.B2(n_442),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1432),
.A2(n_442),
.B(n_443),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1410),
.B(n_445),
.Y(n_1973)
);

AO31x2_ASAP7_75t_L g1974 ( 
.A1(n_1432),
.A2(n_446),
.A3(n_447),
.B(n_448),
.Y(n_1974)
);

AO21x1_ASAP7_75t_L g1975 ( 
.A1(n_1615),
.A2(n_447),
.B(n_448),
.Y(n_1975)
);

AOI21xp33_ASAP7_75t_L g1976 ( 
.A1(n_1608),
.A2(n_449),
.B(n_450),
.Y(n_1976)
);

O2A1O1Ixp5_ASAP7_75t_L g1977 ( 
.A1(n_1432),
.A2(n_449),
.B(n_450),
.C(n_451),
.Y(n_1977)
);

OAI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1432),
.A2(n_451),
.B(n_452),
.Y(n_1978)
);

OAI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1432),
.A2(n_453),
.B(n_454),
.Y(n_1979)
);

INVxp67_ASAP7_75t_L g1980 ( 
.A(n_1637),
.Y(n_1980)
);

BUFx3_ASAP7_75t_L g1981 ( 
.A(n_1439),
.Y(n_1981)
);

AOI21xp33_ASAP7_75t_L g1982 ( 
.A1(n_1608),
.A2(n_456),
.B(n_457),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1432),
.A2(n_458),
.B(n_459),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1410),
.B(n_459),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1432),
.A2(n_461),
.B(n_462),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1410),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1637),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1432),
.A2(n_463),
.B(n_464),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1432),
.A2(n_464),
.B(n_465),
.Y(n_1989)
);

AOI21xp33_ASAP7_75t_L g1990 ( 
.A1(n_1608),
.A2(n_467),
.B(n_468),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1637),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1414),
.A2(n_469),
.B(n_471),
.Y(n_1992)
);

OR2x4_ASAP7_75t_L g1993 ( 
.A(n_1419),
.B(n_469),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1410),
.B(n_471),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1410),
.A2(n_472),
.B1(n_473),
.B2(n_474),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1637),
.Y(n_1996)
);

OAI21x1_ASAP7_75t_SL g1997 ( 
.A1(n_1635),
.A2(n_474),
.B(n_476),
.Y(n_1997)
);

OAI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1432),
.A2(n_476),
.B(n_477),
.Y(n_1998)
);

BUFx2_ASAP7_75t_L g1999 ( 
.A(n_1637),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1432),
.A2(n_477),
.B(n_478),
.Y(n_2000)
);

CKINVDCx6p67_ASAP7_75t_R g2001 ( 
.A(n_1453),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1637),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1635),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1410),
.B(n_479),
.Y(n_2004)
);

OAI21x1_ASAP7_75t_SL g2005 ( 
.A1(n_1635),
.A2(n_480),
.B(n_481),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1986),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1921),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1936),
.Y(n_2008)
);

A2O1A1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1667),
.A2(n_482),
.B(n_483),
.C(n_484),
.Y(n_2009)
);

NAND2x1p5_ASAP7_75t_L g2010 ( 
.A(n_1730),
.B(n_1740),
.Y(n_2010)
);

BUFx2_ASAP7_75t_SL g2011 ( 
.A(n_1669),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1667),
.B(n_485),
.Y(n_2012)
);

AO21x2_ASAP7_75t_L g2013 ( 
.A1(n_1763),
.A2(n_487),
.B(n_489),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1764),
.Y(n_2014)
);

AOI22x1_ASAP7_75t_L g2015 ( 
.A1(n_1847),
.A2(n_490),
.B1(n_491),
.B2(n_492),
.Y(n_2015)
);

INVx4_ASAP7_75t_L g2016 ( 
.A(n_2001),
.Y(n_2016)
);

NAND3xp33_ASAP7_75t_L g2017 ( 
.A(n_1654),
.B(n_491),
.C(n_492),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1745),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1657),
.Y(n_2019)
);

OAI21x1_ASAP7_75t_SL g2020 ( 
.A1(n_1686),
.A2(n_493),
.B(n_494),
.Y(n_2020)
);

BUFx4f_ASAP7_75t_L g2021 ( 
.A(n_1724),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1730),
.B(n_495),
.Y(n_2022)
);

INVx2_ASAP7_75t_SL g2023 ( 
.A(n_1704),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1920),
.B(n_496),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1951),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1784),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1942),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1689),
.Y(n_2028)
);

NOR2xp67_ASAP7_75t_L g2029 ( 
.A(n_1707),
.B(n_497),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1893),
.B(n_497),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_R g2031 ( 
.A(n_1745),
.B(n_498),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_1816),
.Y(n_2032)
);

INVx2_ASAP7_75t_SL g2033 ( 
.A(n_1939),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1943),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1696),
.B(n_498),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1962),
.Y(n_2036)
);

O2A1O1Ixp33_ASAP7_75t_L g2037 ( 
.A1(n_1864),
.A2(n_499),
.B(n_500),
.C(n_1875),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1961),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1964),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1999),
.B(n_1980),
.Y(n_2040)
);

AOI22x1_ASAP7_75t_L g2041 ( 
.A1(n_1919),
.A2(n_1927),
.B1(n_1930),
.B2(n_1924),
.Y(n_2041)
);

NOR2xp67_ASAP7_75t_L g2042 ( 
.A(n_1914),
.B(n_1956),
.Y(n_2042)
);

NAND2x1p5_ASAP7_75t_L g2043 ( 
.A(n_1740),
.B(n_1816),
.Y(n_2043)
);

AO21x2_ASAP7_75t_L g2044 ( 
.A1(n_1959),
.A2(n_1978),
.B(n_1960),
.Y(n_2044)
);

HB1xp67_ASAP7_75t_L g2045 ( 
.A(n_1986),
.Y(n_2045)
);

NAND3xp33_ASAP7_75t_L g2046 ( 
.A(n_1720),
.B(n_1955),
.C(n_1890),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1970),
.Y(n_2047)
);

NAND2x1p5_ASAP7_75t_L g2048 ( 
.A(n_1761),
.B(n_1805),
.Y(n_2048)
);

NOR2x1_ASAP7_75t_R g2049 ( 
.A(n_1735),
.B(n_1759),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_1739),
.B(n_1864),
.Y(n_2050)
);

BUFx4f_ASAP7_75t_L g2051 ( 
.A(n_1952),
.Y(n_2051)
);

INVx4_ASAP7_75t_L g2052 ( 
.A(n_1748),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_SL g2053 ( 
.A1(n_1706),
.A2(n_1998),
.B(n_1979),
.Y(n_2053)
);

OR3x4_ASAP7_75t_SL g2054 ( 
.A(n_1803),
.B(n_1779),
.C(n_1844),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_SL g2055 ( 
.A(n_1713),
.B(n_1776),
.Y(n_2055)
);

INVx2_ASAP7_75t_SL g2056 ( 
.A(n_1675),
.Y(n_2056)
);

AO21x2_ASAP7_75t_L g2057 ( 
.A1(n_1975),
.A2(n_1753),
.B(n_1709),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1773),
.B(n_1987),
.Y(n_2058)
);

BUFx8_ASAP7_75t_L g2059 ( 
.A(n_1811),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_1787),
.Y(n_2060)
);

NOR2x1_ASAP7_75t_R g2061 ( 
.A(n_1687),
.B(n_1716),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1991),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2003),
.Y(n_2063)
);

HB1xp67_ASAP7_75t_L g2064 ( 
.A(n_1952),
.Y(n_2064)
);

AO21x2_ASAP7_75t_L g2065 ( 
.A1(n_1708),
.A2(n_1709),
.B(n_1919),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_1856),
.B(n_1861),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1717),
.Y(n_2067)
);

AO21x2_ASAP7_75t_L g2068 ( 
.A1(n_1708),
.A2(n_1927),
.B(n_1924),
.Y(n_2068)
);

AO21x2_ASAP7_75t_L g2069 ( 
.A1(n_1930),
.A2(n_1935),
.B(n_1933),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1742),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1996),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2002),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1684),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1661),
.Y(n_2074)
);

AO21x2_ASAP7_75t_L g2075 ( 
.A1(n_1933),
.A2(n_1937),
.B(n_1935),
.Y(n_2075)
);

INVx1_ASAP7_75t_SL g2076 ( 
.A(n_1881),
.Y(n_2076)
);

OAI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_1680),
.A2(n_1850),
.B(n_1700),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1677),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1866),
.Y(n_2079)
);

BUFx2_ASAP7_75t_L g2080 ( 
.A(n_1662),
.Y(n_2080)
);

INVx3_ASAP7_75t_L g2081 ( 
.A(n_1866),
.Y(n_2081)
);

AND2x6_ASAP7_75t_L g2082 ( 
.A(n_1973),
.B(n_1748),
.Y(n_2082)
);

OA21x2_ASAP7_75t_L g2083 ( 
.A1(n_1859),
.A2(n_1860),
.B(n_1749),
.Y(n_2083)
);

NAND2x1p5_ASAP7_75t_L g2084 ( 
.A(n_1949),
.B(n_1848),
.Y(n_2084)
);

NAND3xp33_ASAP7_75t_L g2085 ( 
.A(n_1967),
.B(n_1977),
.C(n_1802),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_1789),
.B(n_1952),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1748),
.B(n_1719),
.Y(n_2087)
);

AOI22x1_ASAP7_75t_L g2088 ( 
.A1(n_1937),
.A2(n_1972),
.B1(n_1983),
.B2(n_1968),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1679),
.Y(n_2089)
);

OA21x2_ASAP7_75t_L g2090 ( 
.A1(n_1806),
.A2(n_1972),
.B(n_1968),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1973),
.Y(n_2091)
);

OAI21xp5_ASAP7_75t_SL g2092 ( 
.A1(n_1676),
.A2(n_1743),
.B(n_1733),
.Y(n_2092)
);

BUFx2_ASAP7_75t_R g2093 ( 
.A(n_1824),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1891),
.B(n_1737),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1909),
.A2(n_1931),
.B1(n_1659),
.B2(n_1808),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1758),
.B(n_1825),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1981),
.Y(n_2097)
);

AND2x4_ASAP7_75t_L g2098 ( 
.A(n_1783),
.B(n_1798),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_1866),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1688),
.Y(n_2100)
);

BUFx2_ASAP7_75t_L g2101 ( 
.A(n_1814),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1700),
.B(n_1683),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1660),
.Y(n_2103)
);

AO21x1_ASAP7_75t_L g2104 ( 
.A1(n_1917),
.A2(n_1969),
.B(n_1957),
.Y(n_2104)
);

INVx3_ASAP7_75t_L g2105 ( 
.A(n_1866),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1817),
.Y(n_2106)
);

OA21x2_ASAP7_75t_L g2107 ( 
.A1(n_1983),
.A2(n_1988),
.B(n_1985),
.Y(n_2107)
);

OR2x6_ASAP7_75t_L g2108 ( 
.A(n_1670),
.B(n_1676),
.Y(n_2108)
);

OA21x2_ASAP7_75t_L g2109 ( 
.A1(n_1985),
.A2(n_1989),
.B(n_1988),
.Y(n_2109)
);

AO31x2_ASAP7_75t_L g2110 ( 
.A1(n_1989),
.A2(n_2000),
.A3(n_1854),
.B(n_1821),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1683),
.B(n_1697),
.Y(n_2111)
);

AO21x2_ASAP7_75t_L g2112 ( 
.A1(n_2000),
.A2(n_1827),
.B(n_1818),
.Y(n_2112)
);

INVx2_ASAP7_75t_SL g2113 ( 
.A(n_1953),
.Y(n_2113)
);

INVx3_ASAP7_75t_L g2114 ( 
.A(n_1866),
.Y(n_2114)
);

BUFx3_ASAP7_75t_L g2115 ( 
.A(n_1866),
.Y(n_2115)
);

BUFx3_ASAP7_75t_L g2116 ( 
.A(n_1873),
.Y(n_2116)
);

BUFx10_ASAP7_75t_L g2117 ( 
.A(n_1687),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1710),
.Y(n_2118)
);

CKINVDCx14_ASAP7_75t_R g2119 ( 
.A(n_1733),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1714),
.Y(n_2120)
);

INVx2_ASAP7_75t_SL g2121 ( 
.A(n_1762),
.Y(n_2121)
);

OAI21x1_ASAP7_75t_L g2122 ( 
.A1(n_1869),
.A2(n_1882),
.B(n_1698),
.Y(n_2122)
);

AO22x1_ASAP7_75t_L g2123 ( 
.A1(n_1895),
.A2(n_1743),
.B1(n_1826),
.B2(n_1670),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1652),
.B(n_1941),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_1855),
.B(n_1853),
.Y(n_2125)
);

BUFx4f_ASAP7_75t_L g2126 ( 
.A(n_1716),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1817),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1822),
.Y(n_2128)
);

HB1xp67_ASAP7_75t_L g2129 ( 
.A(n_1848),
.Y(n_2129)
);

BUFx6f_ASAP7_75t_L g2130 ( 
.A(n_1822),
.Y(n_2130)
);

AO21x1_ASAP7_75t_L g2131 ( 
.A1(n_1917),
.A2(n_1969),
.B(n_1957),
.Y(n_2131)
);

OR2x6_ASAP7_75t_L g2132 ( 
.A(n_1751),
.B(n_1797),
.Y(n_2132)
);

INVx4_ASAP7_75t_L g2133 ( 
.A(n_1751),
.Y(n_2133)
);

AO21x1_ASAP7_75t_L g2134 ( 
.A1(n_1908),
.A2(n_1778),
.B(n_1907),
.Y(n_2134)
);

OA21x2_ASAP7_75t_L g2135 ( 
.A1(n_1695),
.A2(n_1692),
.B(n_1849),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_SL g2136 ( 
.A1(n_1785),
.A2(n_1793),
.B(n_1839),
.Y(n_2136)
);

OR2x6_ASAP7_75t_L g2137 ( 
.A(n_1751),
.B(n_1797),
.Y(n_2137)
);

OAI21x1_ASAP7_75t_L g2138 ( 
.A1(n_1756),
.A2(n_1760),
.B(n_1876),
.Y(n_2138)
);

OA21x2_ASAP7_75t_L g2139 ( 
.A1(n_1901),
.A2(n_1780),
.B(n_1715),
.Y(n_2139)
);

AO21x2_ASAP7_75t_L g2140 ( 
.A1(n_1738),
.A2(n_1888),
.B(n_1765),
.Y(n_2140)
);

OAI21x1_ASAP7_75t_L g2141 ( 
.A1(n_1879),
.A2(n_1715),
.B(n_1701),
.Y(n_2141)
);

A2O1A1Ixp33_ASAP7_75t_L g2142 ( 
.A1(n_1769),
.A2(n_1777),
.B(n_1729),
.C(n_1830),
.Y(n_2142)
);

AO21x2_ASAP7_75t_L g2143 ( 
.A1(n_1701),
.A2(n_1727),
.B(n_1750),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1771),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1965),
.B(n_1685),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_1727),
.A2(n_1770),
.B(n_1750),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1656),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1813),
.B(n_1799),
.Y(n_2148)
);

NAND3xp33_ASAP7_75t_L g2149 ( 
.A(n_1767),
.B(n_1897),
.C(n_1796),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1732),
.Y(n_2150)
);

AO21x2_ASAP7_75t_L g2151 ( 
.A1(n_1770),
.A2(n_1912),
.B(n_1699),
.Y(n_2151)
);

BUFx2_ASAP7_75t_R g2152 ( 
.A(n_1691),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1665),
.B(n_1693),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1734),
.B(n_1722),
.Y(n_2154)
);

INVx6_ASAP7_75t_L g2155 ( 
.A(n_1949),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1732),
.Y(n_2156)
);

BUFx3_ASAP7_75t_L g2157 ( 
.A(n_1873),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1774),
.Y(n_2158)
);

AOI22x1_ASAP7_75t_L g2159 ( 
.A1(n_1896),
.A2(n_1834),
.B1(n_1865),
.B2(n_1871),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1774),
.Y(n_2160)
);

OAI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_1832),
.A2(n_1878),
.B(n_1836),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1671),
.Y(n_2162)
);

BUFx10_ASAP7_75t_L g2163 ( 
.A(n_1722),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_1678),
.A2(n_1909),
.B1(n_1768),
.B2(n_1791),
.Y(n_2164)
);

INVxp67_ASAP7_75t_SL g2165 ( 
.A(n_1833),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_1873),
.Y(n_2166)
);

OAI21x1_ASAP7_75t_L g2167 ( 
.A1(n_1810),
.A2(n_1815),
.B(n_1812),
.Y(n_2167)
);

OR2x6_ASAP7_75t_L g2168 ( 
.A(n_1804),
.B(n_1909),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1658),
.B(n_1885),
.Y(n_2169)
);

AOI21x1_ASAP7_75t_L g2170 ( 
.A1(n_1872),
.A2(n_1845),
.B(n_1838),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1792),
.B(n_1809),
.Y(n_2171)
);

OAI21x1_ASAP7_75t_L g2172 ( 
.A1(n_1810),
.A2(n_1815),
.B(n_1812),
.Y(n_2172)
);

AOI221xp5_ASAP7_75t_L g2173 ( 
.A1(n_1826),
.A2(n_1731),
.B1(n_1726),
.B2(n_1778),
.C(n_1889),
.Y(n_2173)
);

BUFx8_ASAP7_75t_L g2174 ( 
.A(n_1741),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1671),
.Y(n_2175)
);

OAI21x1_ASAP7_75t_L g2176 ( 
.A1(n_1772),
.A2(n_1775),
.B(n_1674),
.Y(n_2176)
);

AOI22xp33_ASAP7_75t_L g2177 ( 
.A1(n_1808),
.A2(n_1777),
.B1(n_1668),
.B2(n_1729),
.Y(n_2177)
);

INVxp67_ASAP7_75t_SL g2178 ( 
.A(n_1833),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1791),
.B(n_1851),
.Y(n_2179)
);

AO21x2_ASAP7_75t_L g2180 ( 
.A1(n_1785),
.A2(n_1845),
.B(n_1838),
.Y(n_2180)
);

BUFx3_ASAP7_75t_L g2181 ( 
.A(n_1948),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1766),
.B(n_1843),
.Y(n_2182)
);

BUFx3_ASAP7_75t_L g2183 ( 
.A(n_1948),
.Y(n_2183)
);

BUFx3_ASAP7_75t_L g2184 ( 
.A(n_1948),
.Y(n_2184)
);

OAI21x1_ASAP7_75t_L g2185 ( 
.A1(n_1772),
.A2(n_1775),
.B(n_1674),
.Y(n_2185)
);

AO21x2_ASAP7_75t_L g2186 ( 
.A1(n_1944),
.A2(n_2005),
.B(n_1997),
.Y(n_2186)
);

NAND2x1p5_ASAP7_75t_L g2187 ( 
.A(n_1958),
.B(n_1681),
.Y(n_2187)
);

OA21x2_ASAP7_75t_L g2188 ( 
.A1(n_1858),
.A2(n_1867),
.B(n_1862),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1672),
.Y(n_2189)
);

OAI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_1653),
.A2(n_1655),
.B(n_1984),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_1958),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_1958),
.Y(n_2192)
);

HB1xp67_ASAP7_75t_L g2193 ( 
.A(n_1666),
.Y(n_2193)
);

OAI21x1_ASAP7_75t_L g2194 ( 
.A1(n_1682),
.A2(n_1819),
.B(n_1896),
.Y(n_2194)
);

INVx4_ASAP7_75t_L g2195 ( 
.A(n_1681),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1835),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1813),
.B(n_1794),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_SL g2198 ( 
.A1(n_1906),
.A2(n_1653),
.B(n_1655),
.Y(n_2198)
);

OR2x6_ASAP7_75t_L g2199 ( 
.A(n_1804),
.B(n_1757),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1911),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1911),
.Y(n_2201)
);

OAI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_1916),
.A2(n_2004),
.B(n_1918),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1908),
.B(n_1880),
.Y(n_2203)
);

BUFx2_ASAP7_75t_L g2204 ( 
.A(n_1857),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1835),
.B(n_1828),
.Y(n_2205)
);

OA21x2_ASAP7_75t_L g2206 ( 
.A1(n_1870),
.A2(n_1904),
.B(n_1837),
.Y(n_2206)
);

BUFx2_ASAP7_75t_SL g2207 ( 
.A(n_1842),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1874),
.Y(n_2208)
);

OAI21x1_ASAP7_75t_L g2209 ( 
.A1(n_1819),
.A2(n_1746),
.B(n_1871),
.Y(n_2209)
);

AO21x2_ASAP7_75t_L g2210 ( 
.A1(n_1872),
.A2(n_1752),
.B(n_1807),
.Y(n_2210)
);

OAI21x1_ASAP7_75t_L g2211 ( 
.A1(n_1834),
.A2(n_1865),
.B(n_1666),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_1857),
.Y(n_2212)
);

HB1xp67_ASAP7_75t_L g2213 ( 
.A(n_1916),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_1892),
.B(n_1801),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1918),
.Y(n_2215)
);

BUFx3_ASAP7_75t_L g2216 ( 
.A(n_1841),
.Y(n_2216)
);

OAI21x1_ASAP7_75t_L g2217 ( 
.A1(n_1747),
.A2(n_1744),
.B(n_1820),
.Y(n_2217)
);

INVx4_ASAP7_75t_L g2218 ( 
.A(n_1840),
.Y(n_2218)
);

AND2x4_ASAP7_75t_L g2219 ( 
.A(n_1846),
.B(n_1863),
.Y(n_2219)
);

OAI21x1_ASAP7_75t_L g2220 ( 
.A1(n_1747),
.A2(n_1945),
.B(n_1913),
.Y(n_2220)
);

OAI21x1_ASAP7_75t_L g2221 ( 
.A1(n_1947),
.A2(n_1992),
.B(n_1823),
.Y(n_2221)
);

AO31x2_ASAP7_75t_L g2222 ( 
.A1(n_1900),
.A2(n_1807),
.A3(n_1703),
.B(n_1954),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1922),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1922),
.Y(n_2224)
);

OAI21x1_ASAP7_75t_L g2225 ( 
.A1(n_1887),
.A2(n_1782),
.B(n_1786),
.Y(n_2225)
);

AO21x2_ASAP7_75t_L g2226 ( 
.A1(n_1902),
.A2(n_1788),
.B(n_1800),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1923),
.Y(n_2227)
);

INVx2_ASAP7_75t_SL g2228 ( 
.A(n_1993),
.Y(n_2228)
);

OAI21x1_ASAP7_75t_L g2229 ( 
.A1(n_1887),
.A2(n_1790),
.B(n_1984),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1794),
.B(n_1795),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_1993),
.B(n_1883),
.Y(n_2231)
);

NOR2xp67_ASAP7_75t_L g2232 ( 
.A(n_1673),
.B(n_1718),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_1902),
.A2(n_1880),
.B(n_1884),
.Y(n_2233)
);

BUFx3_ASAP7_75t_L g2234 ( 
.A(n_1840),
.Y(n_2234)
);

NAND2x1p5_ASAP7_75t_L g2235 ( 
.A(n_1712),
.B(n_1868),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1899),
.B(n_1898),
.Y(n_2236)
);

OAI21x1_ASAP7_75t_SL g2237 ( 
.A1(n_1928),
.A2(n_1946),
.B(n_1934),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_1795),
.B(n_1938),
.Y(n_2238)
);

BUFx4f_ASAP7_75t_L g2239 ( 
.A(n_1664),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_1963),
.Y(n_2240)
);

INVx3_ASAP7_75t_SL g2241 ( 
.A(n_1725),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_1898),
.B(n_1899),
.Y(n_2242)
);

HB1xp67_ASAP7_75t_L g2243 ( 
.A(n_1963),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1966),
.B(n_1894),
.Y(n_2244)
);

AO21x2_ASAP7_75t_L g2245 ( 
.A1(n_1829),
.A2(n_1831),
.B(n_1884),
.Y(n_2245)
);

OAI21x1_ASAP7_75t_L g2246 ( 
.A1(n_1966),
.A2(n_1852),
.B(n_1905),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_1711),
.B(n_1736),
.Y(n_2247)
);

OAI21x1_ASAP7_75t_L g2248 ( 
.A1(n_1929),
.A2(n_1994),
.B(n_1781),
.Y(n_2248)
);

INVx3_ASAP7_75t_L g2249 ( 
.A(n_1711),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1668),
.B(n_1711),
.Y(n_2250)
);

OAI21x1_ASAP7_75t_L g2251 ( 
.A1(n_1703),
.A2(n_1995),
.B(n_1971),
.Y(n_2251)
);

AO21x2_ASAP7_75t_L g2252 ( 
.A1(n_1663),
.A2(n_1990),
.B(n_1982),
.Y(n_2252)
);

INVx1_ASAP7_75t_SL g2253 ( 
.A(n_1932),
.Y(n_2253)
);

OA21x2_ASAP7_75t_L g2254 ( 
.A1(n_1663),
.A2(n_1915),
.B(n_1990),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_1926),
.B(n_1694),
.Y(n_2255)
);

OAI21x1_ASAP7_75t_L g2256 ( 
.A1(n_1910),
.A2(n_1995),
.B(n_1971),
.Y(n_2256)
);

CKINVDCx20_ASAP7_75t_R g2257 ( 
.A(n_1910),
.Y(n_2257)
);

OAI21x1_ASAP7_75t_L g2258 ( 
.A1(n_1940),
.A2(n_1903),
.B(n_1877),
.Y(n_2258)
);

AO31x2_ASAP7_75t_L g2259 ( 
.A1(n_1940),
.A2(n_1705),
.A3(n_1723),
.B(n_1974),
.Y(n_2259)
);

OA21x2_ASAP7_75t_L g2260 ( 
.A1(n_1915),
.A2(n_1982),
.B(n_1976),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1702),
.Y(n_2261)
);

NAND3xp33_ASAP7_75t_L g2262 ( 
.A(n_1925),
.B(n_1950),
.C(n_1976),
.Y(n_2262)
);

OAI21x1_ASAP7_75t_L g2263 ( 
.A1(n_1886),
.A2(n_1754),
.B(n_1926),
.Y(n_2263)
);

BUFx4_ASAP7_75t_SL g2264 ( 
.A(n_1728),
.Y(n_2264)
);

CKINVDCx20_ASAP7_75t_R g2265 ( 
.A(n_1755),
.Y(n_2265)
);

BUFx2_ASAP7_75t_L g2266 ( 
.A(n_1702),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_1702),
.Y(n_2267)
);

OAI21x1_ASAP7_75t_SL g2268 ( 
.A1(n_1690),
.A2(n_1763),
.B(n_1706),
.Y(n_2268)
);

BUFx3_ASAP7_75t_L g2269 ( 
.A(n_1724),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1921),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1921),
.Y(n_2271)
);

INVx4_ASAP7_75t_L g2272 ( 
.A(n_2001),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1721),
.Y(n_2273)
);

BUFx4_ASAP7_75t_SL g2274 ( 
.A(n_1669),
.Y(n_2274)
);

OAI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_1667),
.A2(n_1422),
.B(n_1414),
.Y(n_2275)
);

AOI22x1_ASAP7_75t_L g2276 ( 
.A1(n_1847),
.A2(n_1410),
.B1(n_1924),
.B2(n_1919),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1764),
.Y(n_2277)
);

INVx8_ASAP7_75t_L g2278 ( 
.A(n_1724),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1921),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_1730),
.B(n_1635),
.Y(n_2280)
);

OAI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_1667),
.A2(n_1422),
.B(n_1414),
.Y(n_2281)
);

INVx4_ASAP7_75t_L g2282 ( 
.A(n_2001),
.Y(n_2282)
);

INVx5_ASAP7_75t_L g2283 ( 
.A(n_1745),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_1680),
.A2(n_1667),
.B(n_1432),
.Y(n_2284)
);

OAI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_1880),
.A2(n_1410),
.B1(n_1637),
.B2(n_1635),
.Y(n_2285)
);

OR2x2_ASAP7_75t_L g2286 ( 
.A(n_1920),
.B(n_1637),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_1745),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1764),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_1920),
.B(n_1637),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1921),
.Y(n_2290)
);

AOI22x1_ASAP7_75t_L g2291 ( 
.A1(n_1847),
.A2(n_1410),
.B1(n_1924),
.B2(n_1919),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_1986),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1667),
.B(n_1637),
.Y(n_2293)
);

OR2x6_ASAP7_75t_L g2294 ( 
.A(n_1952),
.B(n_1730),
.Y(n_2294)
);

BUFx8_ASAP7_75t_L g2295 ( 
.A(n_1724),
.Y(n_2295)
);

NAND2x1p5_ASAP7_75t_L g2296 ( 
.A(n_1730),
.B(n_1410),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1921),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1921),
.Y(n_2298)
);

OAI21x1_ASAP7_75t_SL g2299 ( 
.A1(n_1690),
.A2(n_1763),
.B(n_1706),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2019),
.Y(n_2300)
);

OR2x6_ASAP7_75t_L g2301 ( 
.A(n_2168),
.B(n_2294),
.Y(n_2301)
);

BUFx2_ASAP7_75t_L g2302 ( 
.A(n_2059),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2019),
.Y(n_2303)
);

OAI22xp5_ASAP7_75t_L g2304 ( 
.A1(n_2119),
.A2(n_2092),
.B1(n_2257),
.B2(n_2051),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2007),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_2295),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2208),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2008),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2027),
.Y(n_2309)
);

CKINVDCx6p67_ASAP7_75t_R g2310 ( 
.A(n_2278),
.Y(n_2310)
);

BUFx12f_ASAP7_75t_L g2311 ( 
.A(n_2295),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2034),
.Y(n_2312)
);

OAI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_2119),
.A2(n_2257),
.B1(n_2051),
.B2(n_2168),
.Y(n_2313)
);

HB1xp67_ASAP7_75t_L g2314 ( 
.A(n_2006),
.Y(n_2314)
);

INVx4_ASAP7_75t_L g2315 ( 
.A(n_2278),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2025),
.Y(n_2316)
);

OAI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2168),
.A2(n_2102),
.B1(n_2293),
.B2(n_2177),
.Y(n_2317)
);

AOI221xp5_ASAP7_75t_L g2318 ( 
.A1(n_2050),
.A2(n_2123),
.B1(n_2177),
.B2(n_2066),
.C(n_2077),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_2232),
.A2(n_2255),
.B1(n_2050),
.B2(n_2125),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2038),
.Y(n_2320)
);

BUFx12f_ASAP7_75t_L g2321 ( 
.A(n_2295),
.Y(n_2321)
);

CKINVDCx10_ASAP7_75t_R g2322 ( 
.A(n_2274),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2289),
.B(n_2066),
.Y(n_2323)
);

AO21x1_ASAP7_75t_SL g2324 ( 
.A1(n_2129),
.A2(n_2064),
.B(n_2091),
.Y(n_2324)
);

BUFx2_ASAP7_75t_L g2325 ( 
.A(n_2059),
.Y(n_2325)
);

AOI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2125),
.A2(n_2265),
.B1(n_2095),
.B2(n_2179),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_2006),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2208),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2039),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_2052),
.Y(n_2330)
);

OAI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2142),
.A2(n_2284),
.B(n_2262),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2047),
.Y(n_2332)
);

HB1xp67_ASAP7_75t_L g2333 ( 
.A(n_2045),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2062),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_2174),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2169),
.B(n_2286),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2071),
.Y(n_2337)
);

INVx6_ASAP7_75t_L g2338 ( 
.A(n_2174),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2072),
.Y(n_2339)
);

INVx2_ASAP7_75t_SL g2340 ( 
.A(n_2278),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2270),
.Y(n_2341)
);

INVx4_ASAP7_75t_L g2342 ( 
.A(n_2021),
.Y(n_2342)
);

INVxp67_ASAP7_75t_L g2343 ( 
.A(n_2061),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2271),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2098),
.B(n_2154),
.Y(n_2345)
);

BUFx3_ASAP7_75t_L g2346 ( 
.A(n_2174),
.Y(n_2346)
);

INVx4_ASAP7_75t_L g2347 ( 
.A(n_2021),
.Y(n_2347)
);

HB1xp67_ASAP7_75t_L g2348 ( 
.A(n_2045),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2279),
.Y(n_2349)
);

CKINVDCx11_ASAP7_75t_R g2350 ( 
.A(n_2016),
.Y(n_2350)
);

INVx6_ASAP7_75t_L g2351 ( 
.A(n_2059),
.Y(n_2351)
);

AO21x1_ASAP7_75t_L g2352 ( 
.A1(n_2203),
.A2(n_2030),
.B(n_2037),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2290),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2297),
.Y(n_2354)
);

HB1xp67_ASAP7_75t_L g2355 ( 
.A(n_2292),
.Y(n_2355)
);

INVx3_ASAP7_75t_L g2356 ( 
.A(n_2052),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2298),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_2280),
.Y(n_2358)
);

BUFx10_ASAP7_75t_L g2359 ( 
.A(n_2028),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2074),
.Y(n_2360)
);

INVx3_ASAP7_75t_L g2361 ( 
.A(n_2280),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2171),
.B(n_2147),
.Y(n_2362)
);

INVx2_ASAP7_75t_SL g2363 ( 
.A(n_2274),
.Y(n_2363)
);

AO21x1_ASAP7_75t_SL g2364 ( 
.A1(n_2129),
.A2(n_2064),
.B(n_2091),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2078),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_2280),
.Y(n_2366)
);

AO21x2_ASAP7_75t_L g2367 ( 
.A1(n_2237),
.A2(n_2198),
.B(n_2053),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2089),
.Y(n_2368)
);

INVx2_ASAP7_75t_SL g2369 ( 
.A(n_2269),
.Y(n_2369)
);

INVx4_ASAP7_75t_L g2370 ( 
.A(n_2016),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2098),
.B(n_2058),
.Y(n_2371)
);

AO21x1_ASAP7_75t_SL g2372 ( 
.A1(n_2095),
.A2(n_2082),
.B(n_2086),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2098),
.B(n_2040),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2100),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2126),
.B(n_2024),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_2028),
.Y(n_2376)
);

AOI22xp33_ASAP7_75t_L g2377 ( 
.A1(n_2265),
.A2(n_2239),
.B1(n_2149),
.B2(n_2173),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2126),
.B(n_2145),
.Y(n_2378)
);

OR2x2_ASAP7_75t_L g2379 ( 
.A(n_2080),
.B(n_2111),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2144),
.Y(n_2380)
);

INVx3_ASAP7_75t_L g2381 ( 
.A(n_2283),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2118),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_2026),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2120),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2073),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2103),
.Y(n_2386)
);

AOI22xp33_ASAP7_75t_L g2387 ( 
.A1(n_2239),
.A2(n_2231),
.B1(n_2236),
.B2(n_2294),
.Y(n_2387)
);

HB1xp67_ASAP7_75t_L g2388 ( 
.A(n_2292),
.Y(n_2388)
);

INVx1_ASAP7_75t_SL g2389 ( 
.A(n_2076),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2063),
.Y(n_2390)
);

BUFx4f_ASAP7_75t_SL g2391 ( 
.A(n_2272),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_2231),
.A2(n_2236),
.B1(n_2294),
.B2(n_2242),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2101),
.B(n_2182),
.Y(n_2393)
);

INVx3_ASAP7_75t_L g2394 ( 
.A(n_2283),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_2155),
.Y(n_2395)
);

INVxp67_ASAP7_75t_L g2396 ( 
.A(n_2108),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2014),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2067),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2033),
.B(n_2036),
.Y(n_2399)
);

AOI22xp33_ASAP7_75t_L g2400 ( 
.A1(n_2236),
.A2(n_2242),
.B1(n_2108),
.B2(n_2175),
.Y(n_2400)
);

BUFx12f_ASAP7_75t_L g2401 ( 
.A(n_2272),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2067),
.Y(n_2402)
);

INVx6_ASAP7_75t_SL g2403 ( 
.A(n_2132),
.Y(n_2403)
);

AOI21x1_ASAP7_75t_L g2404 ( 
.A1(n_2104),
.A2(n_2131),
.B(n_2170),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2070),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2070),
.Y(n_2406)
);

INVxp67_ASAP7_75t_L g2407 ( 
.A(n_2108),
.Y(n_2407)
);

AOI22xp33_ASAP7_75t_L g2408 ( 
.A1(n_2162),
.A2(n_2189),
.B1(n_2156),
.B2(n_2150),
.Y(n_2408)
);

AO21x2_ASAP7_75t_L g2409 ( 
.A1(n_2268),
.A2(n_2299),
.B(n_2261),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2094),
.B(n_2035),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2094),
.B(n_2035),
.Y(n_2411)
);

INVx3_ASAP7_75t_L g2412 ( 
.A(n_2283),
.Y(n_2412)
);

NAND3xp33_ASAP7_75t_L g2413 ( 
.A(n_2159),
.B(n_2009),
.C(n_2267),
.Y(n_2413)
);

AOI22xp33_ASAP7_75t_SL g2414 ( 
.A1(n_2082),
.A2(n_2031),
.B1(n_2133),
.B2(n_2251),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2277),
.Y(n_2415)
);

BUFx3_ASAP7_75t_L g2416 ( 
.A(n_2155),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2275),
.B(n_2281),
.Y(n_2417)
);

AOI22xp33_ASAP7_75t_L g2418 ( 
.A1(n_2263),
.A2(n_2244),
.B1(n_2134),
.B2(n_2161),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2132),
.B(n_2137),
.Y(n_2419)
);

INVx5_ASAP7_75t_L g2420 ( 
.A(n_2132),
.Y(n_2420)
);

BUFx3_ASAP7_75t_L g2421 ( 
.A(n_2155),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2148),
.B(n_2117),
.Y(n_2422)
);

OR2x2_ASAP7_75t_L g2423 ( 
.A(n_2121),
.B(n_2285),
.Y(n_2423)
);

NAND2x1p5_ASAP7_75t_L g2424 ( 
.A(n_2283),
.B(n_2282),
.Y(n_2424)
);

INVx3_ASAP7_75t_L g2425 ( 
.A(n_2099),
.Y(n_2425)
);

INVx2_ASAP7_75t_SL g2426 ( 
.A(n_2269),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2288),
.Y(n_2427)
);

HB1xp67_ASAP7_75t_L g2428 ( 
.A(n_2165),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2012),
.Y(n_2429)
);

INVx3_ASAP7_75t_L g2430 ( 
.A(n_2099),
.Y(n_2430)
);

AOI22xp33_ASAP7_75t_L g2431 ( 
.A1(n_2238),
.A2(n_2252),
.B1(n_2164),
.B2(n_2228),
.Y(n_2431)
);

BUFx2_ASAP7_75t_L g2432 ( 
.A(n_2137),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2096),
.Y(n_2433)
);

INVx1_ASAP7_75t_SL g2434 ( 
.A(n_2093),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2148),
.B(n_2117),
.Y(n_2435)
);

BUFx2_ASAP7_75t_SL g2436 ( 
.A(n_2282),
.Y(n_2436)
);

BUFx4f_ASAP7_75t_SL g2437 ( 
.A(n_2204),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2096),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2022),
.Y(n_2439)
);

CKINVDCx6p67_ASAP7_75t_R g2440 ( 
.A(n_2011),
.Y(n_2440)
);

BUFx2_ASAP7_75t_L g2441 ( 
.A(n_2137),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2254),
.A2(n_2260),
.B1(n_2210),
.B2(n_2088),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2142),
.A2(n_2046),
.B(n_2085),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2148),
.B(n_2117),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2022),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_2026),
.Y(n_2446)
);

BUFx2_ASAP7_75t_L g2447 ( 
.A(n_2199),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2022),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2199),
.Y(n_2449)
);

INVx4_ASAP7_75t_L g2450 ( 
.A(n_2212),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2199),
.Y(n_2451)
);

BUFx3_ASAP7_75t_L g2452 ( 
.A(n_2296),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2296),
.Y(n_2453)
);

OAI21xp33_ASAP7_75t_SL g2454 ( 
.A1(n_2203),
.A2(n_2030),
.B(n_2256),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2200),
.B(n_2201),
.Y(n_2455)
);

OR2x6_ASAP7_75t_L g2456 ( 
.A(n_2084),
.B(n_2087),
.Y(n_2456)
);

HB1xp67_ASAP7_75t_L g2457 ( 
.A(n_2165),
.Y(n_2457)
);

INVxp67_ASAP7_75t_L g2458 ( 
.A(n_2082),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2214),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2214),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2193),
.Y(n_2461)
);

INVx4_ASAP7_75t_SL g2462 ( 
.A(n_2082),
.Y(n_2462)
);

INVxp67_ASAP7_75t_SL g2463 ( 
.A(n_2084),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2193),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2083),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2163),
.B(n_2216),
.Y(n_2466)
);

OR2x6_ASAP7_75t_L g2467 ( 
.A(n_2087),
.B(n_2133),
.Y(n_2467)
);

AOI22xp33_ASAP7_75t_SL g2468 ( 
.A1(n_2082),
.A2(n_2031),
.B1(n_2020),
.B2(n_2256),
.Y(n_2468)
);

OR2x2_ASAP7_75t_L g2469 ( 
.A(n_2153),
.B(n_2124),
.Y(n_2469)
);

INVx11_ASAP7_75t_L g2470 ( 
.A(n_2049),
.Y(n_2470)
);

AOI22xp33_ASAP7_75t_L g2471 ( 
.A1(n_2254),
.A2(n_2260),
.B1(n_2210),
.B2(n_2041),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_L g2472 ( 
.A(n_2197),
.B(n_2230),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2213),
.Y(n_2473)
);

INVx2_ASAP7_75t_SL g2474 ( 
.A(n_2023),
.Y(n_2474)
);

BUFx2_ASAP7_75t_L g2475 ( 
.A(n_2010),
.Y(n_2475)
);

AOI21xp33_ASAP7_75t_SL g2476 ( 
.A1(n_2212),
.A2(n_2010),
.B(n_2241),
.Y(n_2476)
);

BUFx2_ASAP7_75t_L g2477 ( 
.A(n_2043),
.Y(n_2477)
);

HB1xp67_ASAP7_75t_L g2478 ( 
.A(n_2178),
.Y(n_2478)
);

BUFx2_ASAP7_75t_L g2479 ( 
.A(n_2043),
.Y(n_2479)
);

NOR2xp67_ASAP7_75t_L g2480 ( 
.A(n_2113),
.B(n_2056),
.Y(n_2480)
);

INVx1_ASAP7_75t_SL g2481 ( 
.A(n_2207),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2213),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2243),
.Y(n_2483)
);

INVx2_ASAP7_75t_SL g2484 ( 
.A(n_2163),
.Y(n_2484)
);

BUFx10_ASAP7_75t_L g2485 ( 
.A(n_2060),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2243),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2219),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2163),
.B(n_2216),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2219),
.Y(n_2489)
);

INVx2_ASAP7_75t_SL g2490 ( 
.A(n_2097),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2158),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2219),
.Y(n_2492)
);

AOI22xp33_ASAP7_75t_L g2493 ( 
.A1(n_2260),
.A2(n_2044),
.B1(n_2250),
.B2(n_2223),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2160),
.Y(n_2494)
);

BUFx2_ASAP7_75t_L g2495 ( 
.A(n_2116),
.Y(n_2495)
);

BUFx3_ASAP7_75t_L g2496 ( 
.A(n_2116),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2205),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2267),
.Y(n_2498)
);

AOI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_2055),
.A2(n_2241),
.B1(n_2224),
.B2(n_2215),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2227),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2266),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2205),
.B(n_2157),
.Y(n_2502)
);

INVx3_ASAP7_75t_SL g2503 ( 
.A(n_2060),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2235),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_2205),
.B(n_2157),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_2178),
.Y(n_2506)
);

AO22x1_ASAP7_75t_L g2507 ( 
.A1(n_2087),
.A2(n_2253),
.B1(n_2054),
.B2(n_2287),
.Y(n_2507)
);

BUFx3_ASAP7_75t_L g2508 ( 
.A(n_2166),
.Y(n_2508)
);

HB1xp67_ASAP7_75t_L g2509 ( 
.A(n_2240),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2235),
.Y(n_2510)
);

NAND2x1p5_ASAP7_75t_L g2511 ( 
.A(n_2115),
.B(n_2195),
.Y(n_2511)
);

HB1xp67_ASAP7_75t_L g2512 ( 
.A(n_2240),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2032),
.Y(n_2513)
);

AOI22xp33_ASAP7_75t_SL g2514 ( 
.A1(n_2136),
.A2(n_2044),
.B1(n_2206),
.B2(n_2291),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2032),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2029),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2013),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2013),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2233),
.A2(n_2017),
.B1(n_2206),
.B2(n_2048),
.Y(n_2519)
);

OAI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2206),
.A2(n_2048),
.B1(n_2190),
.B2(n_2202),
.Y(n_2520)
);

OAI22xp33_ASAP7_75t_L g2521 ( 
.A1(n_2195),
.A2(n_2188),
.B1(n_2054),
.B2(n_2115),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2166),
.Y(n_2522)
);

AOI222xp33_ASAP7_75t_L g2523 ( 
.A1(n_2247),
.A2(n_2042),
.B1(n_2167),
.B2(n_2172),
.C1(n_2258),
.C2(n_2185),
.Y(n_2523)
);

AND2x4_ASAP7_75t_L g2524 ( 
.A(n_2462),
.B(n_2247),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2305),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2323),
.B(n_2196),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2336),
.B(n_2196),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2371),
.B(n_2393),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2373),
.B(n_2196),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2417),
.B(n_2247),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2345),
.B(n_2378),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2469),
.B(n_2196),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2379),
.B(n_2234),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2410),
.B(n_2234),
.Y(n_2534)
);

INVx3_ASAP7_75t_L g2535 ( 
.A(n_2511),
.Y(n_2535)
);

INVx3_ASAP7_75t_L g2536 ( 
.A(n_2511),
.Y(n_2536)
);

INVxp67_ASAP7_75t_L g2537 ( 
.A(n_2428),
.Y(n_2537)
);

AND2x4_ASAP7_75t_SL g2538 ( 
.A(n_2315),
.B(n_2018),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2411),
.B(n_2375),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2362),
.B(n_2187),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2308),
.Y(n_2541)
);

INVx1_ASAP7_75t_SL g2542 ( 
.A(n_2437),
.Y(n_2542)
);

OR2x2_ASAP7_75t_L g2543 ( 
.A(n_2304),
.B(n_2245),
.Y(n_2543)
);

AOI22xp33_ASAP7_75t_L g2544 ( 
.A1(n_2318),
.A2(n_2276),
.B1(n_2015),
.B2(n_2226),
.Y(n_2544)
);

OR2x2_ASAP7_75t_L g2545 ( 
.A(n_2304),
.B(n_2259),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2362),
.B(n_2187),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2433),
.B(n_2438),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2307),
.Y(n_2548)
);

OAI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2313),
.A2(n_2188),
.B1(n_2152),
.B2(n_2109),
.Y(n_2549)
);

OAI21xp5_ASAP7_75t_SL g2550 ( 
.A1(n_2313),
.A2(n_2018),
.B(n_2287),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2309),
.Y(n_2551)
);

HB1xp67_ASAP7_75t_L g2552 ( 
.A(n_2428),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2312),
.Y(n_2553)
);

INVx4_ASAP7_75t_L g2554 ( 
.A(n_2338),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2335),
.B(n_2218),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2320),
.Y(n_2556)
);

INVx3_ASAP7_75t_L g2557 ( 
.A(n_2452),
.Y(n_2557)
);

NOR2xp33_ASAP7_75t_L g2558 ( 
.A(n_2472),
.B(n_2423),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_2311),
.Y(n_2559)
);

AOI22xp33_ASAP7_75t_SL g2560 ( 
.A1(n_2317),
.A2(n_2188),
.B1(n_2258),
.B2(n_2226),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2329),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2335),
.B(n_2218),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2332),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2346),
.B(n_2167),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2346),
.B(n_2172),
.Y(n_2565)
);

BUFx2_ASAP7_75t_L g2566 ( 
.A(n_2403),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2475),
.B(n_2186),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2334),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2389),
.B(n_2259),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2477),
.B(n_2186),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2337),
.Y(n_2571)
);

AOI22xp33_ASAP7_75t_L g2572 ( 
.A1(n_2318),
.A2(n_2069),
.B1(n_2075),
.B2(n_2068),
.Y(n_2572)
);

INVx3_ASAP7_75t_L g2573 ( 
.A(n_2452),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2479),
.B(n_2249),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2319),
.B(n_2249),
.Y(n_2575)
);

OR2x2_ASAP7_75t_L g2576 ( 
.A(n_2461),
.B(n_2259),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2339),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2319),
.B(n_2259),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2328),
.Y(n_2579)
);

HB1xp67_ASAP7_75t_L g2580 ( 
.A(n_2457),
.Y(n_2580)
);

BUFx3_ASAP7_75t_L g2581 ( 
.A(n_2338),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2341),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2472),
.B(n_2110),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2344),
.B(n_2110),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2349),
.B(n_2110),
.Y(n_2585)
);

INVx3_ASAP7_75t_L g2586 ( 
.A(n_2381),
.Y(n_2586)
);

INVx1_ASAP7_75t_SL g2587 ( 
.A(n_2437),
.Y(n_2587)
);

NAND3xp33_ASAP7_75t_L g2588 ( 
.A(n_2377),
.B(n_2109),
.C(n_2107),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2353),
.B(n_2110),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2354),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2357),
.B(n_2176),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2360),
.Y(n_2592)
);

OR2x2_ASAP7_75t_L g2593 ( 
.A(n_2464),
.B(n_2180),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_2310),
.Y(n_2594)
);

OAI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2317),
.A2(n_2107),
.B1(n_2109),
.B2(n_2105),
.Y(n_2595)
);

INVxp67_ASAP7_75t_SL g2596 ( 
.A(n_2457),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2478),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2365),
.Y(n_2598)
);

AND2x4_ASAP7_75t_L g2599 ( 
.A(n_2462),
.B(n_2181),
.Y(n_2599)
);

AOI22xp33_ASAP7_75t_L g2600 ( 
.A1(n_2326),
.A2(n_2075),
.B1(n_2069),
.B2(n_2068),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2368),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2331),
.B(n_2180),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2374),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2380),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2382),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2473),
.B(n_2065),
.Y(n_2606)
);

OR2x2_ASAP7_75t_L g2607 ( 
.A(n_2482),
.B(n_2483),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2384),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2326),
.B(n_2176),
.Y(n_2609)
);

NAND2x1_ASAP7_75t_L g2610 ( 
.A(n_2301),
.B(n_2079),
.Y(n_2610)
);

BUFx3_ASAP7_75t_L g2611 ( 
.A(n_2338),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2386),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2385),
.Y(n_2613)
);

HB1xp67_ASAP7_75t_L g2614 ( 
.A(n_2478),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2465),
.Y(n_2615)
);

INVx1_ASAP7_75t_SL g2616 ( 
.A(n_2436),
.Y(n_2616)
);

AOI22xp33_ASAP7_75t_SL g2617 ( 
.A1(n_2419),
.A2(n_2107),
.B1(n_2139),
.B2(n_2112),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2502),
.B(n_2185),
.Y(n_2618)
);

BUFx2_ASAP7_75t_L g2619 ( 
.A(n_2403),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2408),
.B(n_2065),
.Y(n_2620)
);

INVx2_ASAP7_75t_SL g2621 ( 
.A(n_2315),
.Y(n_2621)
);

HB1xp67_ASAP7_75t_L g2622 ( 
.A(n_2506),
.Y(n_2622)
);

INVx2_ASAP7_75t_SL g2623 ( 
.A(n_2351),
.Y(n_2623)
);

BUFx2_ASAP7_75t_L g2624 ( 
.A(n_2302),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2500),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2491),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2494),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2505),
.B(n_2194),
.Y(n_2628)
);

AOI22xp33_ASAP7_75t_L g2629 ( 
.A1(n_2377),
.A2(n_2112),
.B1(n_2143),
.B2(n_2057),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2486),
.Y(n_2630)
);

OR2x2_ASAP7_75t_L g2631 ( 
.A(n_2399),
.B(n_2390),
.Y(n_2631)
);

AND2x4_ASAP7_75t_SL g2632 ( 
.A(n_2370),
.B(n_2079),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2455),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2325),
.B(n_2194),
.Y(n_2634)
);

AND2x2_ASAP7_75t_L g2635 ( 
.A(n_2466),
.B(n_2488),
.Y(n_2635)
);

BUFx3_ASAP7_75t_L g2636 ( 
.A(n_2424),
.Y(n_2636)
);

BUFx3_ASAP7_75t_L g2637 ( 
.A(n_2424),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2455),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2358),
.B(n_2211),
.Y(n_2639)
);

NOR2x1_ASAP7_75t_L g2640 ( 
.A(n_2370),
.B(n_2081),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2358),
.B(n_2211),
.Y(n_2641)
);

INVx5_ASAP7_75t_L g2642 ( 
.A(n_2351),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2361),
.B(n_2209),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2408),
.B(n_2057),
.Y(n_2644)
);

BUFx2_ASAP7_75t_L g2645 ( 
.A(n_2301),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2397),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2429),
.B(n_2222),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2398),
.Y(n_2648)
);

INVxp67_ASAP7_75t_SL g2649 ( 
.A(n_2506),
.Y(n_2649)
);

HB1xp67_ASAP7_75t_L g2650 ( 
.A(n_2314),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2361),
.B(n_2209),
.Y(n_2651)
);

BUFx2_ASAP7_75t_L g2652 ( 
.A(n_2301),
.Y(n_2652)
);

BUFx3_ASAP7_75t_L g2653 ( 
.A(n_2351),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2402),
.Y(n_2654)
);

AOI22xp5_ASAP7_75t_SL g2655 ( 
.A1(n_2434),
.A2(n_2105),
.B1(n_2114),
.B2(n_2081),
.Y(n_2655)
);

AND2x2_ASAP7_75t_L g2656 ( 
.A(n_2366),
.B(n_2143),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2366),
.B(n_2217),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_2391),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2405),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2490),
.B(n_2481),
.Y(n_2660)
);

AND2x4_ASAP7_75t_L g2661 ( 
.A(n_2462),
.B(n_2183),
.Y(n_2661)
);

AND2x4_ASAP7_75t_L g2662 ( 
.A(n_2420),
.B(n_2183),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2418),
.B(n_2222),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2406),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2392),
.B(n_2217),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2415),
.Y(n_2666)
);

INVx3_ASAP7_75t_L g2667 ( 
.A(n_2381),
.Y(n_2667)
);

HB1xp67_ASAP7_75t_L g2668 ( 
.A(n_2314),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2427),
.Y(n_2669)
);

BUFx3_ASAP7_75t_L g2670 ( 
.A(n_2395),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2300),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2303),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_2327),
.Y(n_2673)
);

INVx3_ASAP7_75t_L g2674 ( 
.A(n_2394),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2392),
.B(n_2181),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2316),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2418),
.B(n_2222),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2419),
.B(n_2184),
.Y(n_2678)
);

INVx4_ASAP7_75t_L g2679 ( 
.A(n_2391),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2493),
.B(n_2222),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2495),
.B(n_2191),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2480),
.B(n_2191),
.Y(n_2682)
);

HB1xp67_ASAP7_75t_L g2683 ( 
.A(n_2333),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_SL g2684 ( 
.A1(n_2432),
.A2(n_2139),
.B1(n_2151),
.B2(n_2135),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2447),
.B(n_2184),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2463),
.B(n_2225),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2420),
.B(n_2114),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2463),
.B(n_2225),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2321),
.Y(n_2689)
);

AOI21xp5_ASAP7_75t_SL g2690 ( 
.A1(n_2458),
.A2(n_2135),
.B(n_2264),
.Y(n_2690)
);

OAI22xp5_ASAP7_75t_L g2691 ( 
.A1(n_2414),
.A2(n_2135),
.B1(n_2139),
.B2(n_2090),
.Y(n_2691)
);

OAI21xp33_ASAP7_75t_L g2692 ( 
.A1(n_2431),
.A2(n_2221),
.B(n_2146),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2348),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2395),
.B(n_2229),
.Y(n_2694)
);

INVx3_ASAP7_75t_L g2695 ( 
.A(n_2394),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2306),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2416),
.B(n_2229),
.Y(n_2697)
);

AND2x4_ASAP7_75t_L g2698 ( 
.A(n_2420),
.B(n_2273),
.Y(n_2698)
);

HB1xp67_ASAP7_75t_L g2699 ( 
.A(n_2348),
.Y(n_2699)
);

OAI21xp33_ASAP7_75t_L g2700 ( 
.A1(n_2431),
.A2(n_2221),
.B(n_2220),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2416),
.B(n_2128),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2421),
.B(n_2127),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2355),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2421),
.B(n_2127),
.Y(n_2704)
);

AO21x1_ASAP7_75t_L g2705 ( 
.A1(n_2521),
.A2(n_2122),
.B(n_2141),
.Y(n_2705)
);

BUFx2_ASAP7_75t_L g2706 ( 
.A(n_2496),
.Y(n_2706)
);

AND2x4_ASAP7_75t_L g2707 ( 
.A(n_2420),
.B(n_2192),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2548),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2528),
.B(n_2509),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2539),
.B(n_2509),
.Y(n_2710)
);

AND2x4_ASAP7_75t_SL g2711 ( 
.A(n_2679),
.B(n_2456),
.Y(n_2711)
);

AOI22xp33_ASAP7_75t_L g2712 ( 
.A1(n_2558),
.A2(n_2372),
.B1(n_2400),
.B2(n_2414),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2525),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2541),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2583),
.B(n_2498),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2551),
.Y(n_2716)
);

OR2x2_ASAP7_75t_L g2717 ( 
.A(n_2631),
.B(n_2388),
.Y(n_2717)
);

OR2x2_ASAP7_75t_L g2718 ( 
.A(n_2607),
.B(n_2388),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2553),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2556),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2526),
.B(n_2512),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2584),
.B(n_2501),
.Y(n_2722)
);

AOI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2549),
.A2(n_2400),
.B1(n_2387),
.B2(n_2499),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2579),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2527),
.B(n_2512),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2635),
.B(n_2324),
.Y(n_2726)
);

INVx4_ASAP7_75t_L g2727 ( 
.A(n_2642),
.Y(n_2727)
);

INVx2_ASAP7_75t_SL g2728 ( 
.A(n_2594),
.Y(n_2728)
);

INVxp67_ASAP7_75t_SL g2729 ( 
.A(n_2596),
.Y(n_2729)
);

AOI22xp33_ASAP7_75t_L g2730 ( 
.A1(n_2558),
.A2(n_2387),
.B1(n_2343),
.B2(n_2468),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2585),
.B(n_2520),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2589),
.B(n_2520),
.Y(n_2732)
);

NOR2xp33_ASAP7_75t_L g2733 ( 
.A(n_2633),
.B(n_2343),
.Y(n_2733)
);

BUFx6f_ASAP7_75t_SL g2734 ( 
.A(n_2679),
.Y(n_2734)
);

OR2x2_ASAP7_75t_L g2735 ( 
.A(n_2552),
.B(n_2459),
.Y(n_2735)
);

HB1xp67_ASAP7_75t_L g2736 ( 
.A(n_2552),
.Y(n_2736)
);

BUFx3_ASAP7_75t_L g2737 ( 
.A(n_2636),
.Y(n_2737)
);

AOI22xp33_ASAP7_75t_SL g2738 ( 
.A1(n_2549),
.A2(n_2441),
.B1(n_2407),
.B2(n_2396),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2561),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2563),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2568),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2531),
.B(n_2364),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2571),
.Y(n_2743)
);

NOR2x1_ASAP7_75t_L g2744 ( 
.A(n_2554),
.B(n_2342),
.Y(n_2744)
);

AND2x2_ASAP7_75t_L g2745 ( 
.A(n_2532),
.B(n_2487),
.Y(n_2745)
);

AND2x4_ASAP7_75t_SL g2746 ( 
.A(n_2554),
.B(n_2456),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_2634),
.B(n_2467),
.Y(n_2747)
);

INVx1_ASAP7_75t_SL g2748 ( 
.A(n_2706),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2529),
.B(n_2489),
.Y(n_2749)
);

AND2x4_ASAP7_75t_L g2750 ( 
.A(n_2564),
.B(n_2467),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2577),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2638),
.B(n_2517),
.Y(n_2752)
);

OR2x2_ASAP7_75t_L g2753 ( 
.A(n_2580),
.B(n_2460),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2547),
.B(n_2492),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2582),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2591),
.B(n_2518),
.Y(n_2756)
);

AOI22xp33_ASAP7_75t_L g2757 ( 
.A1(n_2534),
.A2(n_2468),
.B1(n_2352),
.B2(n_2521),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2533),
.B(n_2497),
.Y(n_2758)
);

BUFx3_ASAP7_75t_L g2759 ( 
.A(n_2636),
.Y(n_2759)
);

OR2x6_ASAP7_75t_SL g2760 ( 
.A(n_2594),
.B(n_2376),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2540),
.B(n_2522),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2590),
.Y(n_2762)
);

HB1xp67_ASAP7_75t_L g2763 ( 
.A(n_2597),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2546),
.B(n_2449),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2592),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2598),
.Y(n_2766)
);

OAI222xp33_ASAP7_75t_L g2767 ( 
.A1(n_2545),
.A2(n_2543),
.B1(n_2467),
.B2(n_2456),
.C1(n_2560),
.C2(n_2655),
.Y(n_2767)
);

OR2x2_ASAP7_75t_L g2768 ( 
.A(n_2597),
.B(n_2614),
.Y(n_2768)
);

NOR2xp33_ASAP7_75t_L g2769 ( 
.A(n_2645),
.B(n_2507),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2601),
.B(n_2603),
.Y(n_2770)
);

BUFx12f_ASAP7_75t_L g2771 ( 
.A(n_2559),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2604),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2605),
.Y(n_2773)
);

BUFx2_ASAP7_75t_L g2774 ( 
.A(n_2637),
.Y(n_2774)
);

INVx1_ASAP7_75t_SL g2775 ( 
.A(n_2614),
.Y(n_2775)
);

NOR2x1p5_ASAP7_75t_L g2776 ( 
.A(n_2581),
.B(n_2342),
.Y(n_2776)
);

INVx3_ASAP7_75t_SL g2777 ( 
.A(n_2696),
.Y(n_2777)
);

OR2x2_ASAP7_75t_L g2778 ( 
.A(n_2622),
.B(n_2596),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2608),
.B(n_2451),
.Y(n_2779)
);

INVx1_ASAP7_75t_SL g2780 ( 
.A(n_2622),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2612),
.B(n_2439),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2613),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2678),
.B(n_2445),
.Y(n_2783)
);

OR2x2_ASAP7_75t_L g2784 ( 
.A(n_2649),
.B(n_2363),
.Y(n_2784)
);

AND2x4_ASAP7_75t_SL g2785 ( 
.A(n_2535),
.B(n_2536),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2593),
.B(n_2443),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2660),
.B(n_2448),
.Y(n_2787)
);

AND2x2_ASAP7_75t_L g2788 ( 
.A(n_2626),
.B(n_2496),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2625),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2630),
.Y(n_2790)
);

INVx4_ASAP7_75t_L g2791 ( 
.A(n_2642),
.Y(n_2791)
);

OAI221xp5_ASAP7_75t_SL g2792 ( 
.A1(n_2550),
.A2(n_2407),
.B1(n_2396),
.B2(n_2458),
.C(n_2440),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2627),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_2637),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2681),
.B(n_2508),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2650),
.B(n_2443),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2701),
.B(n_2508),
.Y(n_2797)
);

AND2x2_ASAP7_75t_SL g2798 ( 
.A(n_2524),
.B(n_2347),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2693),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2702),
.B(n_2453),
.Y(n_2800)
);

BUFx2_ASAP7_75t_L g2801 ( 
.A(n_2624),
.Y(n_2801)
);

OR2x2_ASAP7_75t_L g2802 ( 
.A(n_2649),
.B(n_2537),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2650),
.B(n_2442),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2668),
.B(n_2673),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2703),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2646),
.Y(n_2806)
);

BUFx2_ASAP7_75t_L g2807 ( 
.A(n_2581),
.Y(n_2807)
);

BUFx2_ASAP7_75t_L g2808 ( 
.A(n_2611),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2611),
.Y(n_2809)
);

AND2x2_ASAP7_75t_SL g2810 ( 
.A(n_2524),
.B(n_2632),
.Y(n_2810)
);

HB1xp67_ASAP7_75t_L g2811 ( 
.A(n_2537),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2668),
.B(n_2471),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2648),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2654),
.Y(n_2814)
);

BUFx2_ASAP7_75t_L g2815 ( 
.A(n_2653),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2615),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2659),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2683),
.B(n_2471),
.Y(n_2818)
);

AND2x4_ASAP7_75t_L g2819 ( 
.A(n_2565),
.B(n_2409),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2704),
.B(n_2504),
.Y(n_2820)
);

INVx2_ASAP7_75t_SL g2821 ( 
.A(n_2616),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2683),
.B(n_2523),
.Y(n_2822)
);

AOI222xp33_ASAP7_75t_L g2823 ( 
.A1(n_2542),
.A2(n_2350),
.B1(n_2503),
.B2(n_2347),
.C1(n_2401),
.C2(n_2516),
.Y(n_2823)
);

NOR2x1_ASAP7_75t_L g2824 ( 
.A(n_2653),
.B(n_2450),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2664),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2699),
.B(n_2367),
.Y(n_2826)
);

INVx4_ASAP7_75t_R g2827 ( 
.A(n_2658),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2666),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2669),
.Y(n_2829)
);

AOI22xp33_ASAP7_75t_L g2830 ( 
.A1(n_2575),
.A2(n_2413),
.B1(n_2510),
.B2(n_2435),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2675),
.B(n_2685),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2699),
.Y(n_2832)
);

AOI22xp5_ASAP7_75t_L g2833 ( 
.A1(n_2652),
.A2(n_2422),
.B1(n_2444),
.B2(n_2350),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2770),
.B(n_2578),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2713),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2831),
.B(n_2656),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2731),
.B(n_2732),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2731),
.B(n_2609),
.Y(n_2838)
);

HB1xp67_ASAP7_75t_L g2839 ( 
.A(n_2736),
.Y(n_2839)
);

OR2x2_ASAP7_75t_L g2840 ( 
.A(n_2796),
.B(n_2569),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2714),
.Y(n_2841)
);

INVx3_ASAP7_75t_L g2842 ( 
.A(n_2810),
.Y(n_2842)
);

OR2x2_ASAP7_75t_L g2843 ( 
.A(n_2717),
.B(n_2530),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2715),
.B(n_2530),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2716),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2816),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2732),
.B(n_2628),
.Y(n_2847)
);

INVxp67_ASAP7_75t_SL g2848 ( 
.A(n_2729),
.Y(n_2848)
);

NAND2x1p5_ASAP7_75t_L g2849 ( 
.A(n_2810),
.B(n_2642),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2719),
.Y(n_2850)
);

INVxp67_ASAP7_75t_L g2851 ( 
.A(n_2801),
.Y(n_2851)
);

INVx2_ASAP7_75t_SL g2852 ( 
.A(n_2737),
.Y(n_2852)
);

HB1xp67_ASAP7_75t_L g2853 ( 
.A(n_2736),
.Y(n_2853)
);

NAND4xp25_ASAP7_75t_L g2854 ( 
.A(n_2730),
.B(n_2560),
.C(n_2572),
.D(n_2600),
.Y(n_2854)
);

INVx4_ASAP7_75t_L g2855 ( 
.A(n_2727),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2720),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2708),
.Y(n_2857)
);

OR2x2_ASAP7_75t_L g2858 ( 
.A(n_2796),
.B(n_2576),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2715),
.B(n_2572),
.Y(n_2859)
);

AND2x2_ASAP7_75t_L g2860 ( 
.A(n_2819),
.B(n_2618),
.Y(n_2860)
);

BUFx2_ASAP7_75t_L g2861 ( 
.A(n_2726),
.Y(n_2861)
);

INVxp67_ASAP7_75t_L g2862 ( 
.A(n_2748),
.Y(n_2862)
);

OR2x2_ASAP7_75t_L g2863 ( 
.A(n_2804),
.B(n_2647),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2710),
.B(n_2567),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2709),
.B(n_2570),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2819),
.B(n_2665),
.Y(n_2866)
);

AND2x4_ASAP7_75t_L g2867 ( 
.A(n_2750),
.B(n_2643),
.Y(n_2867)
);

NOR2x1p5_ASAP7_75t_L g2868 ( 
.A(n_2727),
.B(n_2610),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2754),
.B(n_2799),
.Y(n_2869)
);

AND2x4_ASAP7_75t_L g2870 ( 
.A(n_2750),
.B(n_2651),
.Y(n_2870)
);

HB1xp67_ASAP7_75t_L g2871 ( 
.A(n_2763),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2805),
.B(n_2647),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2822),
.B(n_2639),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2748),
.B(n_2606),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2739),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2718),
.B(n_2671),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2822),
.B(n_2641),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2756),
.B(n_2686),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2756),
.B(n_2688),
.Y(n_2879)
);

HB1xp67_ASAP7_75t_L g2880 ( 
.A(n_2763),
.Y(n_2880)
);

AND2x4_ASAP7_75t_SL g2881 ( 
.A(n_2791),
.B(n_2557),
.Y(n_2881)
);

BUFx3_ASAP7_75t_L g2882 ( 
.A(n_2774),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2722),
.B(n_2657),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2740),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2779),
.B(n_2672),
.Y(n_2885)
);

AND2x2_ASAP7_75t_L g2886 ( 
.A(n_2722),
.B(n_2694),
.Y(n_2886)
);

OR2x2_ASAP7_75t_L g2887 ( 
.A(n_2804),
.B(n_2602),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2741),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2786),
.B(n_2697),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2793),
.B(n_2676),
.Y(n_2890)
);

NOR2xp33_ASAP7_75t_L g2891 ( 
.A(n_2733),
.B(n_2623),
.Y(n_2891)
);

AND2x4_ASAP7_75t_SL g2892 ( 
.A(n_2791),
.B(n_2557),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2743),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2751),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2786),
.B(n_2680),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2724),
.Y(n_2896)
);

AND2x4_ASAP7_75t_L g2897 ( 
.A(n_2747),
.B(n_2409),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2832),
.B(n_2790),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2755),
.Y(n_2899)
);

NAND2x1_ASAP7_75t_L g2900 ( 
.A(n_2827),
.B(n_2690),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2762),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2835),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2895),
.B(n_2765),
.Y(n_2903)
);

NAND3x1_ASAP7_75t_L g2904 ( 
.A(n_2842),
.B(n_2742),
.C(n_2824),
.Y(n_2904)
);

AND2x2_ASAP7_75t_L g2905 ( 
.A(n_2861),
.B(n_2721),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2841),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2836),
.B(n_2725),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2836),
.B(n_2747),
.Y(n_2908)
);

NOR2xp67_ASAP7_75t_R g2909 ( 
.A(n_2842),
.B(n_2642),
.Y(n_2909)
);

OR2x2_ASAP7_75t_L g2910 ( 
.A(n_2843),
.B(n_2768),
.Y(n_2910)
);

AND2x4_ASAP7_75t_L g2911 ( 
.A(n_2897),
.B(n_2729),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2895),
.B(n_2837),
.Y(n_2912)
);

OR2x2_ASAP7_75t_L g2913 ( 
.A(n_2887),
.B(n_2775),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2837),
.B(n_2766),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2873),
.B(n_2877),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2873),
.B(n_2772),
.Y(n_2916)
);

HB1xp67_ASAP7_75t_L g2917 ( 
.A(n_2839),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2877),
.B(n_2773),
.Y(n_2918)
);

OR2x2_ASAP7_75t_L g2919 ( 
.A(n_2887),
.B(n_2863),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2860),
.B(n_2795),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2882),
.Y(n_2921)
);

BUFx2_ASAP7_75t_L g2922 ( 
.A(n_2855),
.Y(n_2922)
);

OR2x2_ASAP7_75t_L g2923 ( 
.A(n_2863),
.B(n_2889),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2845),
.Y(n_2924)
);

NAND2x1_ASAP7_75t_L g2925 ( 
.A(n_2855),
.B(n_2821),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2850),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2860),
.B(n_2764),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2856),
.Y(n_2928)
);

NAND2x1p5_ASAP7_75t_L g2929 ( 
.A(n_2855),
.B(n_2798),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2875),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2882),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2846),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2884),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2838),
.B(n_2782),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2847),
.B(n_2761),
.Y(n_2935)
);

HB1xp67_ASAP7_75t_L g2936 ( 
.A(n_2853),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2847),
.B(n_2787),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2888),
.Y(n_2938)
);

HB1xp67_ASAP7_75t_L g2939 ( 
.A(n_2871),
.Y(n_2939)
);

OR2x2_ASAP7_75t_L g2940 ( 
.A(n_2889),
.B(n_2775),
.Y(n_2940)
);

A2O1A1Ixp33_ASAP7_75t_L g2941 ( 
.A1(n_2842),
.A2(n_2711),
.B(n_2621),
.C(n_2792),
.Y(n_2941)
);

OR2x2_ASAP7_75t_L g2942 ( 
.A(n_2840),
.B(n_2858),
.Y(n_2942)
);

AND2x2_ASAP7_75t_SL g2943 ( 
.A(n_2881),
.B(n_2798),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2893),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2894),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2886),
.B(n_2883),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2899),
.Y(n_2947)
);

OR2x6_ASAP7_75t_L g2948 ( 
.A(n_2900),
.B(n_2737),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2838),
.B(n_2858),
.Y(n_2949)
);

INVxp67_ASAP7_75t_L g2950 ( 
.A(n_2880),
.Y(n_2950)
);

NAND2x1_ASAP7_75t_L g2951 ( 
.A(n_2852),
.B(n_2897),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2901),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2898),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2885),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2846),
.Y(n_2955)
);

AND2x4_ASAP7_75t_L g2956 ( 
.A(n_2897),
.B(n_2811),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2890),
.Y(n_2957)
);

INVx3_ASAP7_75t_R g2958 ( 
.A(n_2849),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2942),
.Y(n_2959)
);

INVx1_ASAP7_75t_SL g2960 ( 
.A(n_2943),
.Y(n_2960)
);

OR2x2_ASAP7_75t_L g2961 ( 
.A(n_2919),
.B(n_2840),
.Y(n_2961)
);

AND2x2_ASAP7_75t_L g2962 ( 
.A(n_2908),
.B(n_2866),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2917),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2922),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2946),
.B(n_2866),
.Y(n_2965)
);

NAND4xp75_ASAP7_75t_L g2966 ( 
.A(n_2958),
.B(n_2744),
.C(n_2769),
.D(n_2852),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2912),
.B(n_2878),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2920),
.B(n_2862),
.Y(n_2968)
);

OR2x2_ASAP7_75t_L g2969 ( 
.A(n_2923),
.B(n_2869),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2912),
.B(n_2878),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2936),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2905),
.B(n_2851),
.Y(n_2972)
);

AOI21xp5_ASAP7_75t_L g2973 ( 
.A1(n_2909),
.A2(n_2767),
.B(n_2792),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2939),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2939),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2953),
.B(n_2879),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2907),
.B(n_2927),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2932),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2913),
.Y(n_2979)
);

O2A1O1Ixp33_ASAP7_75t_L g2980 ( 
.A1(n_2925),
.A2(n_2823),
.B(n_2777),
.C(n_2587),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2955),
.Y(n_2981)
);

OR2x2_ASAP7_75t_L g2982 ( 
.A(n_2949),
.B(n_2874),
.Y(n_2982)
);

AOI22xp33_ASAP7_75t_L g2983 ( 
.A1(n_2911),
.A2(n_2854),
.B1(n_2730),
.B2(n_2712),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2949),
.Y(n_2984)
);

AND2x2_ASAP7_75t_L g2985 ( 
.A(n_2937),
.B(n_2935),
.Y(n_2985)
);

AND2x4_ASAP7_75t_L g2986 ( 
.A(n_2948),
.B(n_2867),
.Y(n_2986)
);

OAI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2904),
.A2(n_2738),
.B(n_2767),
.Y(n_2987)
);

AOI22xp5_ASAP7_75t_L g2988 ( 
.A1(n_2903),
.A2(n_2738),
.B1(n_2712),
.B2(n_2733),
.Y(n_2988)
);

NOR2xp33_ASAP7_75t_L g2989 ( 
.A(n_2957),
.B(n_2777),
.Y(n_2989)
);

AOI32xp33_ASAP7_75t_L g2990 ( 
.A1(n_2911),
.A2(n_2892),
.A3(n_2881),
.B1(n_2769),
.B2(n_2711),
.Y(n_2990)
);

O2A1O1Ixp33_ASAP7_75t_L g2991 ( 
.A1(n_2941),
.A2(n_2823),
.B(n_2689),
.C(n_2474),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2915),
.B(n_2879),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_SL g2993 ( 
.A1(n_2929),
.A2(n_2734),
.B1(n_2794),
.B2(n_2759),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2902),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2915),
.B(n_2883),
.Y(n_2995)
);

AOI31xp33_ASAP7_75t_L g2996 ( 
.A1(n_2929),
.A2(n_2849),
.A3(n_2728),
.B(n_2891),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2906),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2903),
.B(n_2859),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_L g2999 ( 
.A1(n_2956),
.A2(n_2757),
.B1(n_2723),
.B2(n_2830),
.Y(n_2999)
);

NAND2x1p5_ASAP7_75t_L g3000 ( 
.A(n_2909),
.B(n_2759),
.Y(n_3000)
);

AOI21xp5_ASAP7_75t_L g3001 ( 
.A1(n_2948),
.A2(n_2757),
.B(n_2848),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2924),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_2921),
.B(n_2867),
.Y(n_3003)
);

AND2x2_ASAP7_75t_L g3004 ( 
.A(n_2931),
.B(n_2867),
.Y(n_3004)
);

OR2x2_ASAP7_75t_L g3005 ( 
.A(n_2916),
.B(n_2834),
.Y(n_3005)
);

AOI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2916),
.A2(n_2734),
.B1(n_2891),
.B2(n_2830),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_SL g3007 ( 
.A(n_2956),
.B(n_2892),
.Y(n_3007)
);

NAND3xp33_ASAP7_75t_L g3008 ( 
.A(n_2950),
.B(n_2811),
.C(n_2784),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2961),
.Y(n_3009)
);

INVxp67_ASAP7_75t_SL g3010 ( 
.A(n_2980),
.Y(n_3010)
);

OAI222xp33_ASAP7_75t_L g3011 ( 
.A1(n_2960),
.A2(n_2951),
.B1(n_2948),
.B2(n_2918),
.C1(n_2934),
.C2(n_2940),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2978),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2975),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2983),
.B(n_2950),
.Y(n_3014)
);

OAI221xp5_ASAP7_75t_L g3015 ( 
.A1(n_2987),
.A2(n_2918),
.B1(n_2914),
.B2(n_2934),
.C(n_2954),
.Y(n_3015)
);

AOI22xp5_ASAP7_75t_L g3016 ( 
.A1(n_2988),
.A2(n_2914),
.B1(n_2844),
.B2(n_2886),
.Y(n_3016)
);

NAND4xp25_ASAP7_75t_L g3017 ( 
.A(n_2987),
.B(n_2450),
.C(n_2619),
.D(n_2566),
.Y(n_3017)
);

INVx1_ASAP7_75t_SL g3018 ( 
.A(n_2964),
.Y(n_3018)
);

OR2x2_ASAP7_75t_L g3019 ( 
.A(n_2982),
.B(n_2910),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2994),
.Y(n_3020)
);

OA21x2_ASAP7_75t_L g3021 ( 
.A1(n_2973),
.A2(n_3001),
.B(n_2966),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2981),
.Y(n_3022)
);

OAI21xp5_ASAP7_75t_L g3023 ( 
.A1(n_2980),
.A2(n_2640),
.B(n_2794),
.Y(n_3023)
);

OAI21xp33_ASAP7_75t_SL g3024 ( 
.A1(n_2996),
.A2(n_2868),
.B(n_2776),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2998),
.B(n_2926),
.Y(n_3025)
);

NAND3xp33_ASAP7_75t_L g3026 ( 
.A(n_3001),
.B(n_2952),
.C(n_2930),
.Y(n_3026)
);

AOI32xp33_ASAP7_75t_L g3027 ( 
.A1(n_2993),
.A2(n_2746),
.A3(n_2809),
.B1(n_2815),
.B2(n_2807),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2986),
.B(n_2870),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2974),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2973),
.A2(n_2632),
.B(n_2746),
.Y(n_3030)
);

AOI22xp5_ASAP7_75t_L g3031 ( 
.A1(n_2999),
.A2(n_2870),
.B1(n_2933),
.B2(n_2928),
.Y(n_3031)
);

OAI321xp33_ASAP7_75t_L g3032 ( 
.A1(n_2991),
.A2(n_2990),
.A3(n_3006),
.B1(n_3000),
.B2(n_2989),
.C(n_3008),
.Y(n_3032)
);

AOI32xp33_ASAP7_75t_L g3033 ( 
.A1(n_2986),
.A2(n_2972),
.A3(n_2968),
.B1(n_2985),
.B2(n_2977),
.Y(n_3033)
);

AOI21xp33_ASAP7_75t_L g3034 ( 
.A1(n_2963),
.A2(n_2426),
.B(n_2369),
.Y(n_3034)
);

AOI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_2998),
.A2(n_2870),
.B1(n_2944),
.B2(n_2938),
.Y(n_3035)
);

BUFx2_ASAP7_75t_L g3036 ( 
.A(n_3000),
.Y(n_3036)
);

AOI21xp33_ASAP7_75t_L g3037 ( 
.A1(n_2971),
.A2(n_2808),
.B(n_2682),
.Y(n_3037)
);

OAI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_3007),
.A2(n_2588),
.B(n_2945),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_3003),
.B(n_2947),
.Y(n_3039)
);

AOI322xp5_ASAP7_75t_L g3040 ( 
.A1(n_2992),
.A2(n_2864),
.A3(n_2865),
.B1(n_2789),
.B2(n_2600),
.C1(n_2876),
.C2(n_2780),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_3016),
.B(n_2984),
.Y(n_3041)
);

AOI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_3017),
.A2(n_2979),
.B1(n_2959),
.B2(n_2976),
.Y(n_3042)
);

NAND3xp33_ASAP7_75t_L g3043 ( 
.A(n_3010),
.B(n_3002),
.C(n_2997),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_3009),
.Y(n_3044)
);

OAI31xp33_ASAP7_75t_L g3045 ( 
.A1(n_3017),
.A2(n_3004),
.A3(n_2976),
.B(n_2992),
.Y(n_3045)
);

NAND2xp33_ASAP7_75t_SL g3046 ( 
.A(n_3036),
.B(n_2503),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_3028),
.B(n_2965),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_3014),
.B(n_2995),
.Y(n_3048)
);

NOR2xp67_ASAP7_75t_L g3049 ( 
.A(n_3024),
.B(n_2771),
.Y(n_3049)
);

OAI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_3033),
.A2(n_2995),
.B1(n_2970),
.B2(n_2967),
.Y(n_3050)
);

AOI21xp33_ASAP7_75t_L g3051 ( 
.A1(n_3021),
.A2(n_2562),
.B(n_2555),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_3020),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_3032),
.B(n_2696),
.Y(n_3053)
);

NAND2xp33_ASAP7_75t_SL g3054 ( 
.A(n_3023),
.B(n_2967),
.Y(n_3054)
);

NAND3xp33_ASAP7_75t_L g3055 ( 
.A(n_3021),
.B(n_2544),
.C(n_2629),
.Y(n_3055)
);

AOI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_3032),
.A2(n_2970),
.B(n_2340),
.Y(n_3056)
);

OA22x2_ASAP7_75t_L g3057 ( 
.A1(n_3031),
.A2(n_2833),
.B1(n_2785),
.B2(n_2538),
.Y(n_3057)
);

INVxp67_ASAP7_75t_L g3058 ( 
.A(n_3018),
.Y(n_3058)
);

AOI211xp5_ASAP7_75t_L g3059 ( 
.A1(n_3011),
.A2(n_2476),
.B(n_2595),
.C(n_2322),
.Y(n_3059)
);

AOI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_3030),
.A2(n_2538),
.B(n_2785),
.Y(n_3060)
);

OAI21xp33_ASAP7_75t_SL g3061 ( 
.A1(n_3027),
.A2(n_2962),
.B(n_2969),
.Y(n_3061)
);

AOI21xp33_ASAP7_75t_L g3062 ( 
.A1(n_3023),
.A2(n_2670),
.B(n_2826),
.Y(n_3062)
);

AOI21xp5_ASAP7_75t_SL g3063 ( 
.A1(n_3026),
.A2(n_2470),
.B(n_2446),
.Y(n_3063)
);

NAND3xp33_ASAP7_75t_SL g3064 ( 
.A(n_3015),
.B(n_2383),
.C(n_2760),
.Y(n_3064)
);

AOI311xp33_ASAP7_75t_L g3065 ( 
.A1(n_3037),
.A2(n_3034),
.A3(n_3038),
.B(n_3013),
.C(n_3025),
.Y(n_3065)
);

AOI31xp33_ASAP7_75t_L g3066 ( 
.A1(n_3018),
.A2(n_3005),
.A3(n_2661),
.B(n_2599),
.Y(n_3066)
);

AOI221xp5_ASAP7_75t_L g3067 ( 
.A1(n_3035),
.A2(n_2814),
.B1(n_2806),
.B2(n_2813),
.C(n_2829),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_3040),
.B(n_2872),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_3012),
.A2(n_2826),
.B(n_2780),
.Y(n_3069)
);

OAI211xp5_ASAP7_75t_L g3070 ( 
.A1(n_3019),
.A2(n_2629),
.B(n_2544),
.C(n_2692),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_SL g3071 ( 
.A(n_3022),
.B(n_2359),
.Y(n_3071)
);

OAI21xp33_ASAP7_75t_L g3072 ( 
.A1(n_3039),
.A2(n_3029),
.B(n_2812),
.Y(n_3072)
);

NAND4xp25_ASAP7_75t_L g3073 ( 
.A(n_3017),
.B(n_2595),
.C(n_2670),
.D(n_2617),
.Y(n_3073)
);

OAI311xp33_ASAP7_75t_L g3074 ( 
.A1(n_3017),
.A2(n_2700),
.A3(n_2812),
.B1(n_2818),
.C1(n_2803),
.Y(n_3074)
);

NOR2xp33_ASAP7_75t_L g3075 ( 
.A(n_3053),
.B(n_2359),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_L g3076 ( 
.A(n_3049),
.B(n_2485),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_L g3077 ( 
.A(n_3064),
.B(n_2485),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_3058),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_3048),
.B(n_2817),
.Y(n_3079)
);

AOI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_3046),
.A2(n_3063),
.B(n_3064),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_3044),
.B(n_2825),
.Y(n_3081)
);

AOI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_3061),
.A2(n_2783),
.B1(n_2788),
.B2(n_2797),
.Y(n_3082)
);

XNOR2xp5_ASAP7_75t_L g3083 ( 
.A(n_3059),
.B(n_2820),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_3052),
.Y(n_3084)
);

OAI211xp5_ASAP7_75t_L g3085 ( 
.A1(n_3065),
.A2(n_2617),
.B(n_2454),
.C(n_2573),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_3041),
.B(n_2828),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_3067),
.B(n_2781),
.Y(n_3087)
);

O2A1O1Ixp33_ASAP7_75t_L g3088 ( 
.A1(n_3056),
.A2(n_2484),
.B(n_2513),
.C(n_2515),
.Y(n_3088)
);

AOI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_3066),
.A2(n_2818),
.B(n_2803),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_3068),
.B(n_3050),
.Y(n_3090)
);

INVxp67_ASAP7_75t_L g3091 ( 
.A(n_3071),
.Y(n_3091)
);

AOI21xp33_ASAP7_75t_L g3092 ( 
.A1(n_3043),
.A2(n_2667),
.B(n_2586),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_3042),
.Y(n_3093)
);

AO21x1_ASAP7_75t_L g3094 ( 
.A1(n_3054),
.A2(n_2519),
.B(n_2687),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_3047),
.B(n_2758),
.Y(n_3095)
);

OAI21xp33_ASAP7_75t_SL g3096 ( 
.A1(n_3045),
.A2(n_2778),
.B(n_2802),
.Y(n_3096)
);

AOI21xp33_ASAP7_75t_SL g3097 ( 
.A1(n_3057),
.A2(n_2412),
.B(n_2599),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_3051),
.B(n_2573),
.Y(n_3098)
);

NAND3xp33_ASAP7_75t_L g3099 ( 
.A(n_3055),
.B(n_2514),
.C(n_2684),
.Y(n_3099)
);

NOR2xp33_ASAP7_75t_L g3100 ( 
.A(n_3057),
.B(n_2586),
.Y(n_3100)
);

AND5x1_ASAP7_75t_L g3101 ( 
.A(n_3080),
.B(n_3074),
.C(n_3060),
.D(n_3069),
.E(n_3073),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_3093),
.B(n_3072),
.Y(n_3102)
);

OA22x2_ASAP7_75t_L g3103 ( 
.A1(n_3090),
.A2(n_3070),
.B1(n_3062),
.B2(n_2661),
.Y(n_3103)
);

NOR2x1_ASAP7_75t_L g3104 ( 
.A(n_3077),
.B(n_2412),
.Y(n_3104)
);

NOR3xp33_ASAP7_75t_L g3105 ( 
.A(n_3078),
.B(n_2674),
.C(n_2667),
.Y(n_3105)
);

AOI22x1_ASAP7_75t_L g3106 ( 
.A1(n_3083),
.A2(n_3091),
.B1(n_3084),
.B2(n_3089),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_3075),
.B(n_2800),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_3094),
.B(n_3096),
.Y(n_3108)
);

NAND3xp33_ASAP7_75t_SL g3109 ( 
.A(n_3088),
.B(n_2264),
.C(n_2705),
.Y(n_3109)
);

OA22x2_ASAP7_75t_L g3110 ( 
.A1(n_3082),
.A2(n_2536),
.B1(n_2535),
.B2(n_2695),
.Y(n_3110)
);

AND4x1_ASAP7_75t_L g3111 ( 
.A(n_3076),
.B(n_2663),
.C(n_2677),
.D(n_2574),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_3081),
.Y(n_3112)
);

AND2x4_ASAP7_75t_L g3113 ( 
.A(n_3098),
.B(n_2749),
.Y(n_3113)
);

AOI22xp5_ASAP7_75t_L g3114 ( 
.A1(n_3100),
.A2(n_2745),
.B1(n_2677),
.B2(n_2663),
.Y(n_3114)
);

INVx1_ASAP7_75t_SL g3115 ( 
.A(n_3079),
.Y(n_3115)
);

NOR3xp33_ASAP7_75t_SL g3116 ( 
.A(n_3085),
.B(n_2519),
.C(n_2691),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_3086),
.Y(n_3117)
);

OAI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_3099),
.A2(n_2514),
.B(n_2644),
.Y(n_3118)
);

HB1xp67_ASAP7_75t_L g3119 ( 
.A(n_3087),
.Y(n_3119)
);

AOI21xp5_ASAP7_75t_L g3120 ( 
.A1(n_3097),
.A2(n_2602),
.B(n_2752),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3095),
.Y(n_3121)
);

NOR3xp33_ASAP7_75t_L g3122 ( 
.A(n_3109),
.B(n_3102),
.C(n_3108),
.Y(n_3122)
);

AND2x2_ASAP7_75t_SL g3123 ( 
.A(n_3119),
.B(n_2330),
.Y(n_3123)
);

NAND3xp33_ASAP7_75t_SL g3124 ( 
.A(n_3116),
.B(n_3092),
.C(n_2644),
.Y(n_3124)
);

NOR2x1_ASAP7_75t_L g3125 ( 
.A(n_3104),
.B(n_2330),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_3115),
.B(n_3092),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_3113),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_3112),
.Y(n_3128)
);

NOR3xp33_ASAP7_75t_L g3129 ( 
.A(n_3104),
.B(n_2356),
.C(n_2674),
.Y(n_3129)
);

NOR2x1_ASAP7_75t_L g3130 ( 
.A(n_3117),
.B(n_2356),
.Y(n_3130)
);

OA21x2_ASAP7_75t_L g3131 ( 
.A1(n_3106),
.A2(n_3121),
.B(n_3114),
.Y(n_3131)
);

INVxp67_ASAP7_75t_SL g3132 ( 
.A(n_3101),
.Y(n_3132)
);

NAND3xp33_ASAP7_75t_L g3133 ( 
.A(n_3105),
.B(n_2695),
.C(n_2684),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_3113),
.B(n_2857),
.Y(n_3134)
);

NAND3xp33_ASAP7_75t_SL g3135 ( 
.A(n_3111),
.B(n_3118),
.C(n_3103),
.Y(n_3135)
);

NOR3xp33_ASAP7_75t_L g3136 ( 
.A(n_3120),
.B(n_2248),
.C(n_2404),
.Y(n_3136)
);

NAND3xp33_ASAP7_75t_L g3137 ( 
.A(n_3107),
.B(n_2130),
.C(n_2106),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_3110),
.B(n_2752),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_3115),
.B(n_2896),
.Y(n_3139)
);

XOR2xp5_ASAP7_75t_L g3140 ( 
.A(n_3132),
.B(n_2662),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3128),
.Y(n_3141)
);

NOR2x1_ASAP7_75t_L g3142 ( 
.A(n_3135),
.B(n_2367),
.Y(n_3142)
);

NOR2x1p5_ASAP7_75t_L g3143 ( 
.A(n_3127),
.B(n_2662),
.Y(n_3143)
);

NOR2x1_ASAP7_75t_L g3144 ( 
.A(n_3131),
.B(n_2140),
.Y(n_3144)
);

BUFx2_ASAP7_75t_L g3145 ( 
.A(n_3130),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_3139),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_3134),
.Y(n_3147)
);

XNOR2xp5_ASAP7_75t_L g3148 ( 
.A(n_3122),
.B(n_2687),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_3123),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_3138),
.Y(n_3150)
);

NOR2x1_ASAP7_75t_L g3151 ( 
.A(n_3131),
.B(n_3124),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_3151),
.B(n_3126),
.Y(n_3152)
);

NOR3xp33_ASAP7_75t_L g3153 ( 
.A(n_3141),
.B(n_3133),
.C(n_3137),
.Y(n_3153)
);

AND2x4_ASAP7_75t_L g3154 ( 
.A(n_3143),
.B(n_3125),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3146),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3141),
.Y(n_3156)
);

XNOR2xp5_ASAP7_75t_L g3157 ( 
.A(n_3140),
.B(n_3129),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_3147),
.Y(n_3158)
);

XOR2xp5_ASAP7_75t_L g3159 ( 
.A(n_3148),
.B(n_2735),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3150),
.Y(n_3160)
);

OAI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_3152),
.A2(n_3142),
.B(n_3149),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_3158),
.B(n_3145),
.Y(n_3162)
);

BUFx2_ASAP7_75t_L g3163 ( 
.A(n_3155),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3156),
.Y(n_3164)
);

OAI22x1_ASAP7_75t_L g3165 ( 
.A1(n_3157),
.A2(n_3144),
.B1(n_3136),
.B2(n_2707),
.Y(n_3165)
);

OAI21x1_ASAP7_75t_L g3166 ( 
.A1(n_3162),
.A2(n_3160),
.B(n_3159),
.Y(n_3166)
);

AOI211xp5_ASAP7_75t_L g3167 ( 
.A1(n_3161),
.A2(n_3153),
.B(n_3154),
.C(n_2691),
.Y(n_3167)
);

XNOR2x2_ASAP7_75t_L g3168 ( 
.A(n_3164),
.B(n_3154),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3163),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_3161),
.Y(n_3170)
);

OAI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_3169),
.A2(n_3165),
.B1(n_2620),
.B2(n_2753),
.Y(n_3171)
);

OA21x2_ASAP7_75t_L g3172 ( 
.A1(n_3170),
.A2(n_2248),
.B(n_2138),
.Y(n_3172)
);

AOI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_3167),
.A2(n_2140),
.B1(n_2707),
.B2(n_2698),
.Y(n_3173)
);

INVx5_ASAP7_75t_L g3174 ( 
.A(n_3168),
.Y(n_3174)
);

INVx3_ASAP7_75t_L g3175 ( 
.A(n_3174),
.Y(n_3175)
);

OAI21x1_ASAP7_75t_L g3176 ( 
.A1(n_3173),
.A2(n_3166),
.B(n_2246),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_3175),
.B(n_3171),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_3177),
.A2(n_3175),
.B(n_3176),
.Y(n_3178)
);

OR2x2_ASAP7_75t_L g3179 ( 
.A(n_3178),
.B(n_3172),
.Y(n_3179)
);

AOI22xp33_ASAP7_75t_L g3180 ( 
.A1(n_3179),
.A2(n_2698),
.B1(n_2425),
.B2(n_2430),
.Y(n_3180)
);


endmodule