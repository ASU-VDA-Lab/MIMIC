module fake_jpeg_16863_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_11),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_45),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_34),
.B1(n_20),
.B2(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_48),
.B1(n_59),
.B2(n_63),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_18),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_52),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_28),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_53),
.B(n_28),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_18),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_28),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_44),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_20),
.B1(n_26),
.B2(n_35),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_22),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_26),
.B1(n_25),
.B2(n_30),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_65),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_86),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_69),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_68),
.B(n_77),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_81),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_20),
.B1(n_35),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_74),
.A2(n_93),
.B1(n_97),
.B2(n_105),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_19),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_80),
.B(n_90),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_83),
.A2(n_102),
.B(n_61),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_19),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

NAND2x1_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_16),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_87),
.B(n_100),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_94),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_44),
.B(n_42),
.C(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_31),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_98),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_31),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_16),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_61),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_16),
.B(n_27),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_42),
.B1(n_17),
.B2(n_21),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_19),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_108),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_19),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_21),
.B1(n_17),
.B2(n_32),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_74),
.B1(n_73),
.B2(n_105),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_86),
.C(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_119),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_61),
.C(n_16),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_82),
.A2(n_17),
.B1(n_24),
.B2(n_27),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_98),
.B1(n_27),
.B2(n_24),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_133),
.B(n_101),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_79),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g187 ( 
.A(n_136),
.B(n_144),
.C(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_138),
.B1(n_149),
.B2(n_151),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_90),
.B1(n_82),
.B2(n_71),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_96),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_80),
.B(n_78),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_150),
.B(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_69),
.Y(n_148)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_90),
.B(n_87),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_72),
.B1(n_95),
.B2(n_94),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_89),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_153),
.B(n_155),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_24),
.B1(n_104),
.B2(n_81),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_157),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_129),
.B(n_33),
.Y(n_195)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_164),
.Y(n_198)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_92),
.B1(n_91),
.B2(n_85),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_163),
.A2(n_119),
.B1(n_110),
.B2(n_111),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_126),
.B(n_10),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_33),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_114),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_16),
.B(n_33),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_143),
.B1(n_142),
.B2(n_144),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_123),
.B1(n_113),
.B2(n_124),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_168),
.A2(n_200),
.B1(n_166),
.B2(n_146),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_135),
.B1(n_113),
.B2(n_126),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_140),
.B1(n_16),
.B2(n_33),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_184),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_108),
.C(n_124),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_179),
.C(n_163),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_135),
.B(n_131),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_192),
.B(n_194),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_126),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_147),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_162),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_123),
.B(n_121),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_186),
.A2(n_195),
.B(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_134),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_115),
.B(n_134),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_159),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_29),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_160),
.B1(n_139),
.B2(n_141),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_150),
.A2(n_129),
.B1(n_85),
.B2(n_114),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_204),
.C(n_210),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_143),
.C(n_136),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_218),
.B1(n_170),
.B2(n_171),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_219),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_143),
.C(n_149),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_164),
.C(n_140),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_214),
.C(n_220),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_140),
.C(n_60),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_221),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_60),
.C(n_29),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_223),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_224),
.A2(n_176),
.B1(n_183),
.B2(n_180),
.Y(n_243)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_225),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_181),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_171),
.A2(n_85),
.B1(n_29),
.B2(n_22),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_227),
.A2(n_185),
.B1(n_176),
.B2(n_182),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_183),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_29),
.C(n_22),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_200),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_230),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_184),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_177),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_233),
.C(n_246),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_202),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_234),
.B(n_235),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_202),
.A2(n_169),
.B(n_192),
.C(n_178),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_212),
.B1(n_215),
.B2(n_229),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_250),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_212),
.A2(n_195),
.B1(n_169),
.B2(n_168),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_222),
.Y(n_263)
);

INVxp33_ASAP7_75t_SL g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NOR4xp25_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_194),
.C(n_187),
.D(n_198),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_169),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_252),
.B(n_3),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_253),
.A2(n_257),
.B1(n_258),
.B2(n_243),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_210),
.C(n_207),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_259),
.C(n_269),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_208),
.B1(n_214),
.B2(n_223),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_213),
.B1(n_215),
.B2(n_217),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_220),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_218),
.B1(n_215),
.B2(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_240),
.B(n_247),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_264),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_271),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_29),
.C(n_22),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_240),
.A2(n_9),
.B1(n_14),
.B2(n_12),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_3),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_240),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_11),
.B1(n_9),
.B2(n_8),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_256),
.B(n_244),
.Y(n_274)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_276),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_251),
.C(n_233),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_279),
.C(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_251),
.C(n_246),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_245),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_286),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_242),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_22),
.C(n_29),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_3),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_253),
.B1(n_267),
.B2(n_266),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_287),
.A2(n_288),
.B1(n_266),
.B2(n_258),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_260),
.A2(n_237),
.B1(n_248),
.B2(n_5),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_261),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_282),
.A2(n_263),
.B1(n_269),
.B2(n_259),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_293),
.B(n_301),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_7),
.B(n_9),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_298),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_300),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_22),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_275),
.B(n_8),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_302),
.B(n_284),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_276),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_311),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_307),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_295),
.A2(n_281),
.B1(n_277),
.B2(n_279),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_290),
.B(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_273),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_296),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_296),
.C(n_298),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_313),
.B(n_314),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_316),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_302),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_295),
.Y(n_318)
);

AOI31xp67_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_319),
.A3(n_4),
.B(n_5),
.Y(n_323)
);

A2O1A1O1Ixp25_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_293),
.B(n_5),
.C(n_6),
.D(n_4),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_320),
.A2(n_308),
.B(n_307),
.Y(n_322)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_326),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_324),
.A3(n_321),
.B1(n_317),
.B2(n_315),
.C1(n_325),
.C2(n_318),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_4),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_6),
.Y(n_330)
);


endmodule