module fake_jpeg_266_n_214 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_214);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_28),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_1),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_20),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx5_ASAP7_75t_SL g89 ( 
.A(n_78),
.Y(n_89)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_70),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_84),
.B1(n_82),
.B2(n_79),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_90),
.B1(n_95),
.B2(n_83),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_58),
.B1(n_54),
.B2(n_67),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_54),
.B1(n_58),
.B2(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_97),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_67),
.B1(n_65),
.B2(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_63),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_114),
.B1(n_59),
.B2(n_53),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_55),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_106),
.C(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_76),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_76),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_82),
.B1(n_84),
.B2(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_64),
.B1(n_71),
.B2(n_73),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_69),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_74),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_64),
.B1(n_75),
.B2(n_62),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_78),
.B1(n_65),
.B2(n_62),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_125),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_95),
.B1(n_96),
.B2(n_57),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_136),
.B1(n_11),
.B2(n_12),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_89),
.B(n_78),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_26),
.B(n_50),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_96),
.B1(n_88),
.B2(n_89),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_135),
.B1(n_137),
.B2(n_13),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_130),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_57),
.B1(n_65),
.B2(n_75),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_73),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_69),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_134),
.B(n_4),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_99),
.A2(n_59),
.B1(n_53),
.B2(n_3),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

AO22x1_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_111),
.B1(n_110),
.B2(n_100),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_143),
.B(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_145),
.B(n_159),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_135),
.A2(n_116),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_148),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_129),
.B1(n_138),
.B2(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_129),
.B1(n_138),
.B2(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_152),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_153),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_136),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_157),
.B1(n_160),
.B2(n_16),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_161),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_125),
.B(n_12),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_31),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_174),
.B1(n_177),
.B2(n_19),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_15),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_170),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_16),
.B(n_17),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_179),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_152),
.C(n_142),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_36),
.C(n_49),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_150),
.B1(n_146),
.B2(n_155),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_185),
.B1(n_188),
.B2(n_190),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_177),
.Y(n_198)
);

XOR2x2_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_35),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_179),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_37),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_175),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_188)
);

OAI321xp33_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_51),
.A3(n_24),
.B1(n_27),
.B2(n_30),
.C(n_32),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_162),
.B1(n_166),
.B2(n_164),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_194),
.C(n_196),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_195),
.Y(n_201)
);

OA21x2_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_165),
.B(n_162),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_198),
.C(n_189),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_203),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_189),
.C(n_186),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_195),
.C(n_192),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_204),
.A2(n_195),
.B(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_182),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_171),
.B(n_163),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_208),
.B(n_204),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_206),
.B(n_193),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_173),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_169),
.B(n_40),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_41),
.B1(n_45),
.B2(n_47),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_48),
.Y(n_214)
);


endmodule