module fake_jpeg_16620_n_269 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_269);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_154;
wire n_76;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_28),
.A2(n_21),
.B1(n_24),
.B2(n_15),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_26),
.Y(n_57)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_21),
.B1(n_24),
.B2(n_15),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_16),
.C(n_14),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_61),
.Y(n_80)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_21),
.B1(n_26),
.B2(n_22),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_22),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_36),
.B1(n_34),
.B2(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_42),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_28),
.B1(n_21),
.B2(n_49),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_28),
.B1(n_39),
.B2(n_36),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_81),
.CI(n_85),
.CON(n_98),
.SN(n_98)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_42),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_57),
.B(n_15),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_88),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_62),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_52),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_74),
.C(n_16),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_94),
.B1(n_72),
.B2(n_85),
.Y(n_106)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_28),
.B1(n_53),
.B2(n_46),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_104),
.B1(n_89),
.B2(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_77),
.B(n_26),
.Y(n_111)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_13),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_13),
.B(n_17),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_53),
.B1(n_60),
.B2(n_58),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_106),
.B(n_120),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_80),
.B1(n_63),
.B2(n_50),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_117),
.B1(n_118),
.B2(n_84),
.Y(n_137)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_94),
.B1(n_98),
.B2(n_97),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_123),
.C(n_101),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_55),
.B1(n_83),
.B2(n_82),
.Y(n_117)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_45),
.B1(n_84),
.B2(n_40),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_122),
.A2(n_98),
.B1(n_93),
.B2(n_104),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_29),
.C(n_48),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_87),
.B(n_88),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_132),
.C(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_95),
.Y(n_131)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_29),
.C(n_66),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_103),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_13),
.B1(n_34),
.B2(n_32),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_140),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_40),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_14),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_145),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_102),
.B1(n_34),
.B2(n_32),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_112),
.B1(n_34),
.B2(n_33),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_8),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

CKINVDCx12_ASAP7_75t_R g147 ( 
.A(n_108),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_122),
.C(n_125),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_151),
.C(n_152),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_114),
.C(n_110),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_110),
.C(n_107),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_170),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_127),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_156),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_120),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_111),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_107),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_169),
.B1(n_144),
.B2(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_76),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_126),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

BUFx4f_ASAP7_75t_SL g173 ( 
.A(n_160),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_129),
.B(n_137),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_185),
.B1(n_169),
.B2(n_161),
.Y(n_195)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_143),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_179),
.A2(n_164),
.B(n_12),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_150),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_148),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_146),
.B1(n_76),
.B2(n_2),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_168),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_23),
.B1(n_20),
.B2(n_17),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_59),
.B1(n_32),
.B2(n_17),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_23),
.B1(n_20),
.B2(n_32),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_23),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_20),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_156),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_8),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_195),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_193),
.C(n_205),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_151),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_152),
.B1(n_154),
.B2(n_163),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_201),
.B1(n_172),
.B2(n_173),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_189),
.B(n_184),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_203),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_206),
.B(n_10),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_181),
.A2(n_59),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_44),
.C(n_31),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_11),
.B(n_10),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_213),
.B1(n_216),
.B2(n_220),
.Y(n_223)
);

NOR2x1_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_198),
.B1(n_174),
.B2(n_190),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_215),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_180),
.B1(n_185),
.B2(n_33),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_195),
.A2(n_33),
.B1(n_30),
.B2(n_18),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_33),
.B1(n_30),
.B2(n_19),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_9),
.B1(n_11),
.B2(n_8),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_44),
.B(n_27),
.C(n_31),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_218),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_5),
.B1(n_7),
.B2(n_6),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_222),
.B(n_224),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_193),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_202),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_44),
.C(n_27),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_232),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_7),
.B(n_6),
.Y(n_227)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_230),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_19),
.Y(n_230)
);

OAI31xp67_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_19),
.A3(n_27),
.B(n_3),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_5),
.B1(n_1),
.B2(n_4),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_16),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_240),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_16),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_243),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_19),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_228),
.C(n_226),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_250),
.C(n_236),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_232),
.B(n_230),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_253),
.B(n_252),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_29),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_25),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_244),
.Y(n_255)
);

NOR2x1_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_0),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_241),
.A3(n_4),
.B1(n_0),
.B2(n_30),
.C1(n_16),
.C2(n_27),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_256),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_257),
.A2(n_258),
.B(n_259),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_16),
.B(n_4),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_246),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g263 ( 
.A1(n_262),
.A2(n_246),
.B(n_4),
.Y(n_263)
);

OAI21x1_ASAP7_75t_SL g265 ( 
.A1(n_263),
.A2(n_264),
.B(n_31),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_261),
.B(n_31),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_SL g267 ( 
.A(n_266),
.B(n_260),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_31),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_31),
.Y(n_269)
);


endmodule