module fake_aes_8537_n_1264 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1264);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1264;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_822;
wire n_706;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_315;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_659;
wire n_432;
wire n_386;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_274;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g274 ( .A(n_273), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_189), .Y(n_275) );
INVxp33_ASAP7_75t_SL g276 ( .A(n_148), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_18), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_117), .Y(n_278) );
CKINVDCx16_ASAP7_75t_R g279 ( .A(n_207), .Y(n_279) );
CKINVDCx16_ASAP7_75t_R g280 ( .A(n_151), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_61), .Y(n_281) );
INVxp67_ASAP7_75t_SL g282 ( .A(n_67), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_39), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_200), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_194), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_149), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_222), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_113), .Y(n_288) );
CKINVDCx16_ASAP7_75t_R g289 ( .A(n_178), .Y(n_289) );
CKINVDCx16_ASAP7_75t_R g290 ( .A(n_225), .Y(n_290) );
CKINVDCx14_ASAP7_75t_R g291 ( .A(n_213), .Y(n_291) );
INVxp33_ASAP7_75t_SL g292 ( .A(n_155), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_263), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_215), .Y(n_294) );
CKINVDCx14_ASAP7_75t_R g295 ( .A(n_210), .Y(n_295) );
INVxp33_ASAP7_75t_SL g296 ( .A(n_159), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_180), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_117), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_137), .Y(n_299) );
INVxp33_ASAP7_75t_SL g300 ( .A(n_59), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_260), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_179), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_26), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_165), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_216), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_230), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_234), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_5), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_171), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_251), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_211), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_186), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_105), .Y(n_314) );
INVxp33_ASAP7_75t_SL g315 ( .A(n_239), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_190), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_198), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_93), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_75), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_59), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g321 ( .A(n_204), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_209), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_250), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_3), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_122), .B(n_205), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_45), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_72), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_99), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_112), .Y(n_329) );
CKINVDCx16_ASAP7_75t_R g330 ( .A(n_65), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_71), .Y(n_331) );
INVxp33_ASAP7_75t_L g332 ( .A(n_152), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_163), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_265), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_68), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_110), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_118), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_157), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_132), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_97), .Y(n_340) );
INVxp33_ASAP7_75t_L g341 ( .A(n_106), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_147), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_129), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_114), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_154), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_1), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_99), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_272), .Y(n_348) );
CKINVDCx16_ASAP7_75t_R g349 ( .A(n_253), .Y(n_349) );
CKINVDCx16_ASAP7_75t_R g350 ( .A(n_17), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_269), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_270), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_96), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_57), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_2), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_71), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_83), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_264), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_110), .Y(n_359) );
INVxp33_ASAP7_75t_L g360 ( .A(n_121), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_241), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_63), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_82), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_182), .Y(n_364) );
XNOR2x1_ASAP7_75t_L g365 ( .A(n_139), .B(n_160), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_156), .Y(n_366) );
INVxp33_ASAP7_75t_SL g367 ( .A(n_123), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_58), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_93), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g370 ( .A(n_252), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_49), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_177), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_62), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_52), .Y(n_374) );
INVxp33_ASAP7_75t_SL g375 ( .A(n_109), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_74), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_249), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_237), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_150), .Y(n_379) );
CKINVDCx16_ASAP7_75t_R g380 ( .A(n_2), .Y(n_380) );
INVxp33_ASAP7_75t_SL g381 ( .A(n_1), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_32), .Y(n_382) );
INVxp33_ASAP7_75t_L g383 ( .A(n_20), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_58), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_124), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_5), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_172), .Y(n_387) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_85), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_28), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_38), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_235), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_248), .Y(n_392) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_158), .B(n_169), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_28), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_41), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_85), .Y(n_396) );
CKINVDCx14_ASAP7_75t_R g397 ( .A(n_267), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_4), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_100), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_50), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_10), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_262), .Y(n_402) );
INVxp33_ASAP7_75t_SL g403 ( .A(n_214), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_300), .A2(n_6), .B1(n_0), .B2(n_3), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_327), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_327), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_311), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_378), .B(n_0), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_368), .B(n_6), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_327), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_378), .B(n_7), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_372), .B(n_7), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_274), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_274), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_372), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_284), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_311), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_368), .B(n_8), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_385), .B(n_8), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_311), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_372), .B(n_9), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_385), .B(n_9), .Y(n_422) );
OAI22xp5_ASAP7_75t_SL g423 ( .A1(n_362), .A2(n_12), .B1(n_10), .B2(n_11), .Y(n_423) );
INVx6_ASAP7_75t_L g424 ( .A(n_379), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_334), .B(n_11), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_358), .B(n_12), .Y(n_426) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_298), .B(n_13), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_311), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_341), .B(n_360), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_311), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_284), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_285), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_285), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_379), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_286), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_332), .B(n_13), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_286), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_283), .B(n_14), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_313), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_383), .B(n_14), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_313), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_429), .B(n_279), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_420), .Y(n_443) );
OR2x6_ASAP7_75t_L g444 ( .A(n_419), .B(n_365), .Y(n_444) );
AND2x2_ASAP7_75t_SL g445 ( .A(n_419), .B(n_280), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_420), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_419), .B(n_415), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_415), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_415), .Y(n_449) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_412), .A2(n_421), .B(n_438), .Y(n_450) );
BUFx10_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_419), .B(n_298), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_415), .B(n_343), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_420), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_439), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_413), .B(n_414), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_405), .B(n_343), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_419), .B(n_319), .Y(n_460) );
BUFx3_ASAP7_75t_L g461 ( .A(n_424), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_424), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_410), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_410), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_429), .B(n_289), .Y(n_465) );
INVx4_ASAP7_75t_L g466 ( .A(n_424), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_429), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_422), .Y(n_468) );
NAND2xp33_ASAP7_75t_L g469 ( .A(n_413), .B(n_325), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_420), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_410), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_439), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_422), .B(n_290), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_439), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_413), .A2(n_288), .B1(n_304), .B2(n_283), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_422), .B(n_321), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_414), .B(n_416), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_409), .B(n_349), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_439), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_441), .Y(n_480) );
AND2x6_ASAP7_75t_L g481 ( .A(n_427), .B(n_287), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_409), .B(n_370), .Y(n_482) );
AND2x6_ASAP7_75t_L g483 ( .A(n_427), .B(n_293), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_441), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_406), .B(n_352), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_409), .A2(n_375), .B1(n_381), .B2(n_300), .Y(n_486) );
AND2x6_ASAP7_75t_L g487 ( .A(n_418), .B(n_293), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_414), .B(n_352), .Y(n_488) );
NOR2x1p5_ASAP7_75t_L g489 ( .A(n_478), .B(n_408), .Y(n_489) );
BUFx4f_ASAP7_75t_SL g490 ( .A(n_467), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_457), .Y(n_491) );
INVx4_ASAP7_75t_L g492 ( .A(n_451), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_447), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_448), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_447), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_451), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_468), .B(n_418), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_451), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_447), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_468), .B(n_418), .Y(n_500) );
BUFx6f_ASAP7_75t_SL g501 ( .A(n_445), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_447), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_448), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_487), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_448), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_444), .A2(n_404), .B1(n_330), .B2(n_350), .Y(n_506) );
AND3x1_ASAP7_75t_SL g507 ( .A(n_486), .B(n_423), .C(n_278), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_447), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_447), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_451), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_460), .B(n_440), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_445), .B(n_408), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_445), .A2(n_411), .B1(n_436), .B2(n_426), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_445), .B(n_411), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_467), .B(n_442), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_487), .B(n_432), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_451), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_477), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_460), .B(n_425), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_444), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_456), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_487), .B(n_432), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_477), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_452), .B(n_426), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_460), .B(n_436), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_456), .Y(n_527) );
INVx4_ASAP7_75t_L g528 ( .A(n_487), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_487), .B(n_433), .Y(n_529) );
OR2x6_ASAP7_75t_L g530 ( .A(n_444), .B(n_423), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_463), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_456), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_444), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_464), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_456), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_456), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_487), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_464), .Y(n_538) );
BUFx3_ASAP7_75t_L g539 ( .A(n_487), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_473), .A2(n_365), .B1(n_375), .B2(n_412), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_471), .Y(n_541) );
INVx5_ASAP7_75t_L g542 ( .A(n_487), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_471), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_449), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_449), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_487), .B(n_433), .Y(n_546) );
AND3x2_ASAP7_75t_SL g547 ( .A(n_444), .B(n_331), .C(n_319), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_487), .B(n_435), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_453), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_453), .Y(n_550) );
AO22x1_ASAP7_75t_L g551 ( .A1(n_487), .A2(n_292), .B1(n_296), .B2(n_276), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_478), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_444), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_472), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_452), .B(n_275), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_452), .A2(n_437), .B1(n_416), .B2(n_431), .Y(n_556) );
INVxp33_ASAP7_75t_SL g557 ( .A(n_473), .Y(n_557) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_472), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_474), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_476), .B(n_416), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_474), .Y(n_561) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_479), .Y(n_562) );
BUFx2_ASAP7_75t_L g563 ( .A(n_476), .Y(n_563) );
BUFx4f_ASAP7_75t_SL g564 ( .A(n_481), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_460), .Y(n_565) );
INVx4_ASAP7_75t_L g566 ( .A(n_452), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_479), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_460), .Y(n_568) );
INVx4_ASAP7_75t_L g569 ( .A(n_452), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_482), .B(n_437), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_482), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_480), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_452), .Y(n_573) );
BUFx2_ASAP7_75t_L g574 ( .A(n_444), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_491), .A2(n_486), .B1(n_460), .B2(n_465), .Y(n_575) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_498), .Y(n_576) );
OR2x6_ASAP7_75t_L g577 ( .A(n_528), .B(n_442), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_490), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_557), .A2(n_465), .B1(n_469), .B2(n_450), .Y(n_579) );
INVx3_ASAP7_75t_L g580 ( .A(n_492), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_493), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_497), .Y(n_582) );
BUFx12f_ASAP7_75t_L g583 ( .A(n_530), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_493), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_573), .Y(n_585) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_498), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_497), .B(n_465), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_493), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_563), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_542), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_498), .B(n_466), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_566), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_573), .Y(n_593) );
BUFx4f_ASAP7_75t_SL g594 ( .A(n_566), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_501), .A2(n_483), .B1(n_481), .B2(n_380), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_501), .A2(n_481), .B1(n_483), .B2(n_450), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_560), .B(n_469), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_489), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_519), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_507), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_569), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_520), .B(n_450), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_524), .A2(n_475), .B1(n_404), .B2(n_454), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_501), .A2(n_481), .B1(n_483), .B2(n_450), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_570), .B(n_450), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_570), .B(n_282), .Y(n_606) );
BUFx2_ASAP7_75t_L g607 ( .A(n_563), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_492), .Y(n_608) );
INVx3_ASAP7_75t_L g609 ( .A(n_492), .Y(n_609) );
BUFx2_ASAP7_75t_L g610 ( .A(n_537), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_557), .A2(n_454), .B1(n_292), .B2(n_296), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_495), .Y(n_612) );
CKINVDCx11_ASAP7_75t_R g613 ( .A(n_530), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_569), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_518), .Y(n_615) );
INVx8_ASAP7_75t_L g616 ( .A(n_542), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_552), .B(n_324), .Y(n_617) );
AO22x1_ASAP7_75t_L g618 ( .A1(n_521), .A2(n_483), .B1(n_481), .B2(n_315), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_504), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_571), .A2(n_483), .B1(n_481), .B2(n_337), .Y(n_620) );
AND2x4_ASAP7_75t_L g621 ( .A(n_511), .B(n_353), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_520), .A2(n_483), .B1(n_481), .B2(n_431), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_498), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_498), .B(n_466), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_SL g625 ( .A1(n_516), .A2(n_488), .B(n_484), .C(n_480), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_530), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_511), .B(n_388), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_518), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_495), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_499), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_520), .B(n_481), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_514), .A2(n_483), .B1(n_481), .B2(n_431), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_518), .B(n_400), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_558), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_540), .B(n_337), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_515), .A2(n_485), .B1(n_459), .B2(n_329), .C(n_335), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_530), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_528), .Y(n_638) );
BUFx12f_ASAP7_75t_L g639 ( .A(n_526), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_537), .A2(n_367), .B1(n_403), .B2(n_276), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_542), .B(n_459), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_542), .B(n_485), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_512), .B(n_367), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_500), .B(n_483), .Y(n_644) );
INVxp33_ASAP7_75t_SL g645 ( .A(n_521), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_499), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_502), .Y(n_647) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_558), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_539), .A2(n_403), .B1(n_295), .B2(n_397), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_502), .Y(n_650) );
BUFx12f_ASAP7_75t_L g651 ( .A(n_526), .Y(n_651) );
OAI21x1_ASAP7_75t_SL g652 ( .A1(n_528), .A2(n_466), .B(n_297), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_514), .A2(n_483), .B1(n_431), .B2(n_406), .Y(n_653) );
AND2x4_ASAP7_75t_L g654 ( .A(n_542), .B(n_277), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_513), .B(n_466), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_539), .B(n_281), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_504), .A2(n_291), .B1(n_431), .B2(n_382), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_558), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_508), .B(n_336), .Y(n_659) );
NAND2x1p5_ASAP7_75t_L g660 ( .A(n_508), .B(n_466), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_496), .B(n_461), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_574), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_509), .Y(n_663) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_554), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_509), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_510), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_558), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_565), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_533), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_568), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_551), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_559), .Y(n_672) );
AOI21x1_ASAP7_75t_L g673 ( .A1(n_551), .A2(n_441), .B(n_443), .Y(n_673) );
OR2x6_ASAP7_75t_L g674 ( .A(n_517), .B(n_288), .Y(n_674) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_558), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_533), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_559), .Y(n_677) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_562), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_554), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_562), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_525), .B(n_340), .Y(n_681) );
INVx4_ASAP7_75t_L g682 ( .A(n_562), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_561), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_506), .A2(n_384), .B1(n_328), .B2(n_371), .Y(n_684) );
INVx6_ASAP7_75t_L g685 ( .A(n_522), .Y(n_685) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_562), .Y(n_686) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_562), .Y(n_687) );
INVx5_ASAP7_75t_SL g688 ( .A(n_522), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_553), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_538), .A2(n_462), .B(n_461), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_564), .A2(n_441), .B1(n_314), .B2(n_318), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_547), .A2(n_314), .B1(n_318), .B2(n_309), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_556), .B(n_376), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_567), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_496), .B(n_461), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_523), .B(n_275), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_572), .B(n_320), .Y(n_697) );
O2A1O1Ixp5_ASAP7_75t_L g698 ( .A1(n_555), .A2(n_377), .B(n_297), .C(n_299), .Y(n_698) );
NOR2xp33_ASAP7_75t_SL g699 ( .A(n_645), .B(n_510), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_575), .A2(n_534), .B1(n_531), .B2(n_541), .C(n_538), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_684), .A2(n_548), .B1(n_546), .B2(n_529), .C(n_541), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_628), .Y(n_702) );
AND2x4_ASAP7_75t_L g703 ( .A(n_599), .B(n_510), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g704 ( .A(n_578), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_634), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_605), .A2(n_527), .B1(n_545), .B2(n_544), .Y(n_706) );
BUFx3_ASAP7_75t_L g707 ( .A(n_628), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_582), .B(n_543), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_697), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_587), .B(n_543), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_634), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_579), .A2(n_550), .B1(n_549), .B2(n_547), .C(n_344), .Y(n_712) );
INVx3_ASAP7_75t_L g713 ( .A(n_628), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_605), .A2(n_532), .B1(n_536), .B2(n_547), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_634), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_589), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_607), .B(n_532), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_594), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_634), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_659), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_648), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_664), .B(n_536), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_692), .A2(n_535), .B1(n_522), .B2(n_494), .Y(n_723) );
OAI21x1_ASAP7_75t_L g724 ( .A1(n_673), .A2(n_503), .B(n_494), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_577), .A2(n_617), .B1(n_676), .B2(n_669), .Y(n_725) );
AOI21xp33_ASAP7_75t_L g726 ( .A1(n_643), .A2(n_505), .B(n_522), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_672), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_644), .A2(n_505), .B(n_535), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_603), .B(n_535), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_577), .A2(n_535), .B1(n_424), .B2(n_347), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_577), .B(n_346), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_648), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_635), .A2(n_424), .B1(n_354), .B2(n_355), .Y(n_733) );
BUFx2_ASAP7_75t_L g734 ( .A(n_639), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_651), .A2(n_424), .B1(n_356), .B2(n_357), .Y(n_735) );
OR2x6_ASAP7_75t_L g736 ( .A(n_616), .B(n_331), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_648), .Y(n_737) );
INVx2_ASAP7_75t_SL g738 ( .A(n_594), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_648), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_662), .A2(n_424), .B1(n_359), .B2(n_369), .Y(n_740) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_583), .A2(n_689), .B1(n_626), .B2(n_637), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_677), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_675), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_580), .B(n_461), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_621), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_613), .A2(n_374), .B1(n_373), .B2(n_326), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_621), .A2(n_326), .B1(n_386), .B2(n_320), .Y(n_747) );
OAI21xp33_ASAP7_75t_SL g748 ( .A1(n_679), .A2(n_299), .B(n_294), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_598), .B(n_386), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_627), .A2(n_390), .B1(n_394), .B2(n_389), .Y(n_750) );
AND2x4_ASAP7_75t_L g751 ( .A(n_580), .B(n_462), .Y(n_751) );
INVx4_ASAP7_75t_L g752 ( .A(n_616), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_675), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_627), .A2(n_390), .B1(n_394), .B2(n_389), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_675), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_681), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_681), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_675), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_606), .A2(n_396), .B1(n_399), .B2(n_398), .C(n_395), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_664), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_683), .B(n_395), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_612), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_600), .A2(n_398), .B1(n_399), .B2(n_396), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_595), .A2(n_401), .B1(n_301), .B2(n_302), .Y(n_764) );
INVx4_ASAP7_75t_L g765 ( .A(n_616), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_629), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_630), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_671), .A2(n_401), .B1(n_351), .B2(n_364), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_646), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_633), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_595), .A2(n_301), .B1(n_302), .B2(n_294), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_694), .B(n_363), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_597), .A2(n_366), .B1(n_317), .B2(n_305), .Y(n_773) );
BUFx2_ASAP7_75t_L g774 ( .A(n_674), .Y(n_774) );
NAND2x1p5_ASAP7_75t_L g775 ( .A(n_608), .B(n_462), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_611), .B(n_462), .Y(n_776) );
BUFx3_ASAP7_75t_L g777 ( .A(n_576), .Y(n_777) );
BUFx2_ASAP7_75t_L g778 ( .A(n_674), .Y(n_778) );
INVx1_ASAP7_75t_SL g779 ( .A(n_656), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_602), .A2(n_455), .B(n_443), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_674), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_678), .Y(n_782) );
NAND2x1p5_ASAP7_75t_L g783 ( .A(n_608), .B(n_303), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_631), .A2(n_305), .B1(n_306), .B2(n_303), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_597), .A2(n_307), .B1(n_308), .B2(n_306), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_647), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_650), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_653), .B(n_307), .Y(n_788) );
OR2x6_ASAP7_75t_L g789 ( .A(n_610), .B(n_308), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_643), .A2(n_312), .B1(n_316), .B2(n_310), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_653), .B(n_663), .Y(n_791) );
AO31x2_ASAP7_75t_L g792 ( .A1(n_655), .A2(n_417), .A3(n_407), .B(n_312), .Y(n_792) );
AOI222xp33_ASAP7_75t_L g793 ( .A1(n_636), .A2(n_310), .B1(n_316), .B2(n_322), .C1(n_323), .C2(n_402), .Y(n_793) );
AND2x6_ASAP7_75t_L g794 ( .A(n_688), .B(n_322), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_665), .Y(n_795) );
OAI222xp33_ASAP7_75t_L g796 ( .A1(n_640), .A2(n_323), .B1(n_392), .B2(n_387), .C1(n_402), .C2(n_348), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_678), .Y(n_797) );
BUFx3_ASAP7_75t_L g798 ( .A(n_576), .Y(n_798) );
OAI21x1_ASAP7_75t_L g799 ( .A1(n_690), .A2(n_698), .B(n_667), .Y(n_799) );
AND2x4_ASAP7_75t_L g800 ( .A(n_609), .B(n_348), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_668), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_670), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_691), .A2(n_392), .B1(n_387), .B2(n_342), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_609), .B(n_393), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_656), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_585), .Y(n_806) );
INVxp67_ASAP7_75t_L g807 ( .A(n_654), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_632), .B(n_338), .Y(n_808) );
OAI22xp5_ASAP7_75t_SL g809 ( .A1(n_596), .A2(n_391), .B1(n_333), .B2(n_345), .Y(n_809) );
NAND2x1p5_ASAP7_75t_L g810 ( .A(n_615), .B(n_339), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_593), .Y(n_811) );
BUFx3_ASAP7_75t_L g812 ( .A(n_586), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_632), .B(n_361), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_586), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_688), .Y(n_815) );
CKINVDCx11_ASAP7_75t_R g816 ( .A(n_586), .Y(n_816) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_623), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_655), .A2(n_434), .B1(n_417), .B2(n_407), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_686), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_686), .Y(n_820) );
BUFx3_ASAP7_75t_L g821 ( .A(n_623), .Y(n_821) );
AOI21x1_ASAP7_75t_L g822 ( .A1(n_690), .A2(n_417), .B(n_407), .Y(n_822) );
AND2x4_ASAP7_75t_L g823 ( .A(n_615), .B(n_15), .Y(n_823) );
AO31x2_ASAP7_75t_L g824 ( .A1(n_658), .A2(n_417), .A3(n_407), .B(n_443), .Y(n_824) );
OR2x2_ASAP7_75t_L g825 ( .A(n_693), .B(n_15), .Y(n_825) );
INVx3_ASAP7_75t_L g826 ( .A(n_623), .Y(n_826) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_620), .A2(n_434), .B1(n_17), .B2(n_16), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_691), .A2(n_434), .B1(n_428), .B2(n_430), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_581), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_618), .Y(n_830) );
AOI22xp33_ASAP7_75t_SL g831 ( .A1(n_657), .A2(n_434), .B1(n_18), .B2(n_16), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_592), .A2(n_434), .B1(n_428), .B2(n_430), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_619), .A2(n_434), .B1(n_428), .B2(n_430), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_686), .Y(n_834) );
BUFx4f_ASAP7_75t_SL g835 ( .A(n_815), .Y(n_835) );
AO31x2_ASAP7_75t_L g836 ( .A1(n_729), .A2(n_785), .A3(n_828), .B(n_728), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_712), .A2(n_604), .B1(n_596), .B2(n_652), .Y(n_837) );
AND2x4_ASAP7_75t_L g838 ( .A(n_752), .B(n_619), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_781), .B(n_622), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g840 ( .A1(n_781), .A2(n_649), .B1(n_623), .B2(n_688), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_809), .A2(n_642), .B1(n_641), .B2(n_666), .Y(n_841) );
OR2x2_ASAP7_75t_L g842 ( .A(n_716), .B(n_601), .Y(n_842) );
BUFx10_ASAP7_75t_L g843 ( .A(n_794), .Y(n_843) );
INVxp67_ASAP7_75t_L g844 ( .A(n_708), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_708), .B(n_614), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_791), .A2(n_604), .B1(n_588), .B2(n_584), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_727), .Y(n_847) );
NOR2x1_ASAP7_75t_SL g848 ( .A(n_736), .B(n_686), .Y(n_848) );
OA21x2_ASAP7_75t_L g849 ( .A1(n_724), .A2(n_680), .B(n_455), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_742), .Y(n_850) );
INVx3_ASAP7_75t_L g851 ( .A(n_752), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_774), .B(n_660), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_791), .A2(n_682), .B1(n_696), .B2(n_666), .Y(n_853) );
AOI22xp33_ASAP7_75t_SL g854 ( .A1(n_778), .A2(n_794), .B1(n_823), .B2(n_830), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_699), .A2(n_638), .B1(n_590), .B2(n_660), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_808), .A2(n_638), .B1(n_695), .B2(n_661), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_736), .A2(n_687), .B1(n_685), .B2(n_695), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g858 ( .A1(n_736), .A2(n_687), .B1(n_685), .B2(n_661), .Y(n_858) );
AND2x4_ASAP7_75t_L g859 ( .A(n_752), .B(n_687), .Y(n_859) );
AO31x2_ASAP7_75t_L g860 ( .A1(n_780), .A2(n_625), .A3(n_455), .B(n_458), .Y(n_860) );
AOI21xp33_ASAP7_75t_L g861 ( .A1(n_725), .A2(n_624), .B(n_591), .Y(n_861) );
AOI222xp33_ASAP7_75t_L g862 ( .A1(n_759), .A2(n_624), .B1(n_591), .B2(n_685), .C1(n_430), .C2(n_428), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_710), .B(n_731), .Y(n_863) );
OA21x2_ASAP7_75t_L g864 ( .A1(n_799), .A2(n_458), .B(n_470), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_808), .A2(n_428), .B1(n_430), .B2(n_420), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g866 ( .A1(n_789), .A2(n_428), .B1(n_430), .B2(n_420), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g867 ( .A(n_831), .B(n_428), .C(n_420), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_762), .Y(n_868) );
AND2x4_ASAP7_75t_L g869 ( .A(n_765), .B(n_19), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g870 ( .A1(n_700), .A2(n_470), .B(n_458), .Y(n_870) );
BUFx6f_ASAP7_75t_L g871 ( .A(n_816), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_761), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_731), .B(n_756), .Y(n_873) );
NAND2xp5_ASAP7_75t_SL g874 ( .A(n_741), .B(n_446), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_757), .B(n_19), .Y(n_875) );
OAI21x1_ASAP7_75t_L g876 ( .A1(n_822), .A2(n_470), .B(n_446), .Y(n_876) );
OAI22xp33_ASAP7_75t_SL g877 ( .A1(n_789), .A2(n_22), .B1(n_20), .B2(n_21), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_813), .A2(n_446), .B1(n_23), .B2(n_21), .Y(n_878) );
OAI211xp5_ASAP7_75t_L g879 ( .A1(n_793), .A2(n_446), .B(n_24), .C(n_22), .Y(n_879) );
AOI221x1_ASAP7_75t_SL g880 ( .A1(n_749), .A2(n_23), .B1(n_24), .B2(n_25), .C(n_26), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_766), .Y(n_881) );
AOI221xp5_ASAP7_75t_L g882 ( .A1(n_749), .A2(n_446), .B1(n_27), .B2(n_29), .C(n_30), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_761), .Y(n_883) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_825), .A2(n_30), .B1(n_25), .B2(n_27), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_745), .Y(n_885) );
AOI21xp33_ASAP7_75t_SL g886 ( .A1(n_704), .A2(n_31), .B(n_32), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_767), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_801), .Y(n_888) );
OAI221xp5_ASAP7_75t_L g889 ( .A1(n_746), .A2(n_446), .B1(n_33), .B2(n_34), .C(n_35), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_813), .A2(n_446), .B1(n_35), .B2(n_31), .Y(n_890) );
OAI221xp5_ASAP7_75t_L g891 ( .A1(n_763), .A2(n_34), .B1(n_36), .B2(n_37), .C(n_38), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_802), .Y(n_892) );
AOI21x1_ASAP7_75t_L g893 ( .A1(n_804), .A2(n_799), .B(n_711), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_723), .A2(n_36), .B1(n_37), .B2(n_40), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_709), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_779), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_788), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_788), .A2(n_46), .B1(n_48), .B2(n_49), .Y(n_898) );
NOR2xp67_ASAP7_75t_L g899 ( .A(n_704), .B(n_50), .Y(n_899) );
AOI21xp33_ASAP7_75t_L g900 ( .A1(n_776), .A2(n_51), .B(n_52), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_764), .A2(n_51), .B1(n_53), .B2(n_54), .Y(n_901) );
BUFx2_ASAP7_75t_L g902 ( .A(n_794), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_714), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_771), .A2(n_56), .B1(n_60), .B2(n_62), .Y(n_904) );
OAI211xp5_ASAP7_75t_L g905 ( .A1(n_768), .A2(n_60), .B(n_63), .C(n_64), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_770), .A2(n_66), .B1(n_69), .B2(n_70), .Y(n_906) );
OAI22xp33_ASAP7_75t_L g907 ( .A1(n_825), .A2(n_69), .B1(n_70), .B2(n_73), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_769), .B(n_73), .Y(n_908) );
OR2x2_ASAP7_75t_L g909 ( .A(n_717), .B(n_74), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_786), .Y(n_910) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_794), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_772), .Y(n_912) );
OAI211xp5_ASAP7_75t_SL g913 ( .A1(n_747), .A2(n_76), .B(n_77), .C(n_78), .Y(n_913) );
AND2x4_ASAP7_75t_L g914 ( .A(n_765), .B(n_79), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_823), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_915) );
AOI222xp33_ASAP7_75t_L g916 ( .A1(n_750), .A2(n_80), .B1(n_81), .B2(n_82), .C1(n_83), .C2(n_84), .Y(n_916) );
AOI22xp5_ASAP7_75t_L g917 ( .A1(n_703), .A2(n_84), .B1(n_86), .B2(n_87), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_787), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_706), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_919) );
OAI221xp5_ASAP7_75t_L g920 ( .A1(n_754), .A2(n_89), .B1(n_90), .B2(n_91), .C(n_92), .Y(n_920) );
OAI22xp5_ASAP7_75t_SL g921 ( .A1(n_734), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_795), .B(n_94), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_772), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_760), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_703), .A2(n_95), .B1(n_97), .B2(n_98), .Y(n_925) );
CKINVDCx11_ASAP7_75t_R g926 ( .A(n_765), .Y(n_926) );
INVx3_ASAP7_75t_L g927 ( .A(n_707), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_823), .A2(n_95), .B1(n_98), .B2(n_100), .Y(n_928) );
AOI22xp33_ASAP7_75t_SL g929 ( .A1(n_794), .A2(n_101), .B1(n_102), .B2(n_103), .Y(n_929) );
AO31x2_ASAP7_75t_L g930 ( .A1(n_705), .A2(n_101), .A3(n_102), .B(n_104), .Y(n_930) );
AOI22xp33_ASAP7_75t_SL g931 ( .A1(n_794), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_720), .B(n_107), .Y(n_932) );
AOI22xp33_ASAP7_75t_SL g933 ( .A1(n_748), .A2(n_107), .B1(n_108), .B2(n_109), .Y(n_933) );
AOI21xp33_ASAP7_75t_L g934 ( .A1(n_776), .A2(n_108), .B(n_111), .Y(n_934) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_726), .A2(n_185), .B(n_268), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_733), .B(n_111), .Y(n_936) );
INVxp67_ASAP7_75t_L g937 ( .A(n_722), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_722), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_718), .B(n_113), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_790), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_940) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_707), .Y(n_941) );
AND2x6_ASAP7_75t_L g942 ( .A(n_817), .B(n_125), .Y(n_942) );
AOI21xp33_ASAP7_75t_L g943 ( .A1(n_773), .A2(n_116), .B(n_118), .Y(n_943) );
OAI221xp5_ASAP7_75t_L g944 ( .A1(n_735), .A2(n_119), .B1(n_120), .B2(n_121), .C(n_126), .Y(n_944) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_810), .A2(n_119), .B1(n_120), .B2(n_127), .Y(n_945) );
INVx2_ASAP7_75t_L g946 ( .A(n_806), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_800), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_805), .A2(n_128), .B1(n_130), .B2(n_131), .Y(n_948) );
AOI222xp33_ASAP7_75t_L g949 ( .A1(n_796), .A2(n_133), .B1(n_134), .B2(n_135), .C1(n_136), .C2(n_138), .Y(n_949) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_702), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_738), .B(n_140), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g952 ( .A1(n_880), .A2(n_827), .B1(n_803), .B2(n_701), .C(n_784), .Y(n_952) );
OAI21xp33_ASAP7_75t_L g953 ( .A1(n_911), .A2(n_931), .B(n_929), .Y(n_953) );
OAI221xp5_ASAP7_75t_L g954 ( .A1(n_841), .A2(n_740), .B1(n_783), .B2(n_807), .C(n_730), .Y(n_954) );
OA21x2_ASAP7_75t_L g955 ( .A1(n_893), .A2(n_818), .B(n_832), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_888), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_892), .Y(n_957) );
BUFx6f_ASAP7_75t_L g958 ( .A(n_926), .Y(n_958) );
AND2x4_ASAP7_75t_L g959 ( .A(n_851), .B(n_702), .Y(n_959) );
AO21x1_ASAP7_75t_SL g960 ( .A1(n_843), .A2(n_811), .B(n_829), .Y(n_960) );
BUFx2_ASAP7_75t_L g961 ( .A(n_835), .Y(n_961) );
OR2x2_ASAP7_75t_L g962 ( .A(n_863), .B(n_800), .Y(n_962) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_869), .Y(n_963) );
AOI211xp5_ASAP7_75t_L g964 ( .A1(n_921), .A2(n_833), .B(n_713), .C(n_751), .Y(n_964) );
NAND2x1_ASAP7_75t_L g965 ( .A(n_942), .B(n_817), .Y(n_965) );
OR2x2_ASAP7_75t_L g966 ( .A(n_909), .B(n_844), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_847), .Y(n_967) );
INVx3_ASAP7_75t_L g968 ( .A(n_851), .Y(n_968) );
INVx3_ASAP7_75t_L g969 ( .A(n_843), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_850), .Y(n_970) );
NAND3xp33_ASAP7_75t_SL g971 ( .A(n_911), .B(n_775), .C(n_820), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_868), .Y(n_972) );
INVxp67_ASAP7_75t_SL g973 ( .A(n_937), .Y(n_973) );
OR2x2_ASAP7_75t_L g974 ( .A(n_844), .B(n_792), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g975 ( .A1(n_884), .A2(n_744), .B1(n_751), .B2(n_826), .C(n_814), .Y(n_975) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_914), .Y(n_976) );
OAI221xp5_ASAP7_75t_L g977 ( .A1(n_841), .A2(n_775), .B1(n_812), .B2(n_777), .C(n_821), .Y(n_977) );
AOI31xp33_ASAP7_75t_L g978 ( .A1(n_854), .A2(n_834), .A3(n_820), .B(n_819), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_881), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g980 ( .A1(n_902), .A2(n_777), .B1(n_812), .B2(n_798), .Y(n_980) );
OR2x2_ASAP7_75t_L g981 ( .A(n_887), .B(n_910), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_872), .B(n_792), .Y(n_982) );
NAND4xp25_ASAP7_75t_L g983 ( .A(n_916), .B(n_899), .C(n_897), .D(n_898), .Y(n_983) );
INVxp67_ASAP7_75t_R g984 ( .A(n_852), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_918), .Y(n_985) );
AOI211xp5_ASAP7_75t_SL g986 ( .A1(n_884), .A2(n_814), .B(n_826), .C(n_758), .Y(n_986) );
AO21x1_ASAP7_75t_SL g987 ( .A1(n_855), .A2(n_814), .B(n_826), .Y(n_987) );
OAI31xp33_ASAP7_75t_L g988 ( .A1(n_879), .A2(n_834), .A3(n_711), .B(n_715), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_873), .B(n_792), .Y(n_989) );
OAI31xp33_ASAP7_75t_L g990 ( .A1(n_907), .A2(n_753), .A3(n_719), .B(n_797), .Y(n_990) );
INVx2_ASAP7_75t_SL g991 ( .A(n_871), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_839), .B(n_824), .Y(n_992) );
OAI31xp33_ASAP7_75t_L g993 ( .A1(n_907), .A2(n_743), .A3(n_721), .B(n_782), .Y(n_993) );
OR2x2_ASAP7_75t_L g994 ( .A(n_924), .B(n_715), .Y(n_994) );
OAI211xp5_ASAP7_75t_L g995 ( .A1(n_929), .A2(n_755), .B(n_732), .C(n_782), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_883), .B(n_721), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_946), .Y(n_997) );
OAI211xp5_ASAP7_75t_L g998 ( .A1(n_931), .A2(n_758), .B(n_755), .C(n_739), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_885), .Y(n_999) );
NAND3xp33_ASAP7_75t_L g1000 ( .A(n_886), .B(n_737), .C(n_817), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_937), .A2(n_824), .B1(n_142), .B2(n_143), .Y(n_1001) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_859), .B(n_824), .Y(n_1002) );
OA21x2_ASAP7_75t_L g1003 ( .A1(n_876), .A2(n_824), .B(n_144), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_842), .Y(n_1004) );
OAI211xp5_ASAP7_75t_L g1005 ( .A1(n_933), .A2(n_141), .B(n_145), .C(n_146), .Y(n_1005) );
OR2x2_ASAP7_75t_L g1006 ( .A(n_938), .B(n_153), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_908), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_912), .B(n_271), .Y(n_1008) );
OAI221xp5_ASAP7_75t_L g1009 ( .A1(n_837), .A2(n_161), .B1(n_162), .B2(n_164), .C(n_166), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_845), .B(n_167), .Y(n_1010) );
OAI211xp5_ASAP7_75t_SL g1011 ( .A1(n_898), .A2(n_168), .B(n_170), .C(n_173), .Y(n_1011) );
OAI21xp33_ASAP7_75t_L g1012 ( .A1(n_895), .A2(n_174), .B(n_175), .Y(n_1012) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_859), .B(n_176), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_923), .B(n_266), .Y(n_1014) );
OAI31xp33_ASAP7_75t_L g1015 ( .A1(n_877), .A2(n_181), .A3(n_183), .B(n_184), .Y(n_1015) );
NAND3xp33_ASAP7_75t_L g1016 ( .A(n_895), .B(n_187), .C(n_188), .Y(n_1016) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_837), .A2(n_191), .B1(n_192), .B2(n_193), .C(n_195), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_947), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_890), .A2(n_196), .B1(n_197), .B2(n_199), .Y(n_1019) );
OAI31xp33_ASAP7_75t_L g1020 ( .A1(n_913), .A2(n_905), .A3(n_891), .B(n_889), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_890), .A2(n_201), .B1(n_202), .B2(n_203), .Y(n_1021) );
OAI211xp5_ASAP7_75t_L g1022 ( .A1(n_945), .A2(n_206), .B(n_208), .C(n_212), .Y(n_1022) );
NOR3xp33_ASAP7_75t_SL g1023 ( .A(n_920), .B(n_217), .C(n_218), .Y(n_1023) );
AOI221xp5_ASAP7_75t_L g1024 ( .A1(n_943), .A2(n_219), .B1(n_220), .B2(n_221), .C(n_223), .Y(n_1024) );
OAI21x1_ASAP7_75t_SL g1025 ( .A1(n_848), .A2(n_224), .B(n_226), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_915), .A2(n_227), .B1(n_228), .B2(n_229), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_936), .A2(n_231), .B1(n_232), .B2(n_233), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_922), .Y(n_1028) );
OAI221xp5_ASAP7_75t_L g1029 ( .A1(n_940), .A2(n_236), .B1(n_238), .B2(n_240), .C(n_242), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g1030 ( .A1(n_940), .A2(n_243), .B1(n_244), .B2(n_245), .C(n_246), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_939), .Y(n_1031) );
INVx2_ASAP7_75t_L g1032 ( .A(n_860), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_950), .Y(n_1033) );
AOI221xp5_ASAP7_75t_L g1034 ( .A1(n_900), .A2(n_247), .B1(n_254), .B2(n_255), .C(n_257), .Y(n_1034) );
OA211x2_ASAP7_75t_L g1035 ( .A1(n_874), .A2(n_258), .B(n_259), .C(n_261), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_871), .B(n_875), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_838), .B(n_932), .Y(n_1037) );
OAI21xp33_ASAP7_75t_L g1038 ( .A1(n_928), .A2(n_917), .B(n_925), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_982), .Y(n_1039) );
INVx3_ASAP7_75t_L g1040 ( .A(n_965), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_974), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_992), .B(n_930), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1032), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_956), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_989), .B(n_930), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_957), .Y(n_1046) );
OAI211xp5_ASAP7_75t_SL g1047 ( .A1(n_1004), .A2(n_882), .B(n_906), .C(n_896), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_999), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_1033), .B(n_941), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1018), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_996), .Y(n_1051) );
OAI31xp33_ASAP7_75t_L g1052 ( .A1(n_953), .A2(n_944), .A3(n_904), .B(n_919), .Y(n_1052) );
OAI221xp5_ASAP7_75t_L g1053 ( .A1(n_983), .A2(n_903), .B1(n_901), .B2(n_861), .C(n_934), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_967), .Y(n_1054) );
OAI31xp33_ASAP7_75t_L g1055 ( .A1(n_954), .A2(n_858), .A3(n_894), .B(n_866), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_970), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_1002), .Y(n_1057) );
INVx2_ASAP7_75t_SL g1058 ( .A(n_1002), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_972), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_979), .Y(n_1060) );
OAI31xp33_ASAP7_75t_L g1061 ( .A1(n_954), .A2(n_858), .A3(n_866), .B(n_867), .Y(n_1061) );
AOI33xp33_ASAP7_75t_L g1062 ( .A1(n_1031), .A2(n_878), .A3(n_846), .B1(n_840), .B2(n_853), .B3(n_856), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_985), .Y(n_1063) );
INVx1_ASAP7_75t_SL g1064 ( .A(n_961), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_997), .B(n_930), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_981), .B(n_846), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_1003), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_973), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_994), .B(n_950), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1007), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_984), .B(n_941), .Y(n_1071) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_969), .B(n_860), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_1003), .Y(n_1073) );
INVx3_ASAP7_75t_L g1074 ( .A(n_969), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1028), .Y(n_1075) );
AOI31xp33_ASAP7_75t_L g1076 ( .A1(n_964), .A2(n_949), .A3(n_951), .B(n_857), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_952), .A2(n_862), .B1(n_942), .B2(n_927), .Y(n_1077) );
INVx3_ASAP7_75t_L g1078 ( .A(n_968), .Y(n_1078) );
BUFx3_ASAP7_75t_L g1079 ( .A(n_958), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_966), .B(n_836), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_968), .Y(n_1081) );
AOI221xp5_ASAP7_75t_L g1082 ( .A1(n_1038), .A2(n_865), .B1(n_870), .B2(n_948), .C(n_935), .Y(n_1082) );
INVx3_ASAP7_75t_L g1083 ( .A(n_1013), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_962), .B(n_860), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1085 ( .A(n_963), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_976), .B(n_836), .Y(n_1086) );
INVx2_ASAP7_75t_L g1087 ( .A(n_955), .Y(n_1087) );
INVx2_ASAP7_75t_L g1088 ( .A(n_955), .Y(n_1088) );
AND2x4_ASAP7_75t_L g1089 ( .A(n_1013), .B(n_860), .Y(n_1089) );
BUFx3_ASAP7_75t_L g1090 ( .A(n_958), .Y(n_1090) );
BUFx3_ASAP7_75t_L g1091 ( .A(n_958), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1025), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1010), .B(n_864), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_1036), .B(n_836), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_977), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_991), .B(n_942), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_959), .B(n_849), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1006), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_977), .Y(n_1099) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_1037), .B(n_849), .Y(n_1100) );
OAI221xp5_ASAP7_75t_SL g1101 ( .A1(n_1020), .A2(n_975), .B1(n_993), .B2(n_990), .C(n_1015), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_971), .B(n_978), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_995), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1008), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_995), .Y(n_1105) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1014), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_998), .Y(n_1107) );
INVxp67_ASAP7_75t_L g1108 ( .A(n_960), .Y(n_1108) );
AND2x2_ASAP7_75t_SL g1109 ( .A(n_986), .B(n_1034), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1044), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1044), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_1109), .A2(n_1017), .B1(n_1009), .B2(n_1029), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1045), .B(n_987), .Y(n_1113) );
OAI31xp33_ASAP7_75t_L g1114 ( .A1(n_1108), .A2(n_1022), .A3(n_1005), .B(n_998), .Y(n_1114) );
AND2x4_ASAP7_75t_L g1115 ( .A(n_1057), .B(n_1000), .Y(n_1115) );
NOR2xp33_ASAP7_75t_L g1116 ( .A(n_1085), .B(n_1005), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1070), .B(n_988), .Y(n_1117) );
AND2x4_ASAP7_75t_L g1118 ( .A(n_1057), .B(n_1023), .Y(n_1118) );
NOR2xp67_ASAP7_75t_L g1119 ( .A(n_1102), .B(n_1022), .Y(n_1119) );
AND2x4_ASAP7_75t_L g1120 ( .A(n_1072), .B(n_1016), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1070), .B(n_980), .Y(n_1121) );
NAND2xp5_ASAP7_75t_SL g1122 ( .A(n_1109), .B(n_1034), .Y(n_1122) );
INVx2_ASAP7_75t_L g1123 ( .A(n_1043), .Y(n_1123) );
INVx2_ASAP7_75t_SL g1124 ( .A(n_1058), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_1109), .A2(n_1030), .B1(n_1012), .B2(n_1011), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1046), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1046), .Y(n_1127) );
AND3x2_ASAP7_75t_L g1128 ( .A(n_1061), .B(n_1024), .C(n_1035), .Y(n_1128) );
INVx2_ASAP7_75t_L g1129 ( .A(n_1043), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1049), .B(n_1001), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1075), .B(n_1019), .Y(n_1131) );
INVx1_ASAP7_75t_SL g1132 ( .A(n_1064), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1049), .B(n_1021), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1075), .B(n_1026), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1045), .B(n_1027), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1048), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1054), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1054), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1042), .B(n_1084), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1056), .Y(n_1140) );
NAND4xp25_ASAP7_75t_L g1141 ( .A(n_1101), .B(n_1052), .C(n_1080), .D(n_1077), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1056), .Y(n_1142) );
AND4x1_ASAP7_75t_L g1143 ( .A(n_1061), .B(n_1052), .C(n_1055), .D(n_1062), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1042), .B(n_1084), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1069), .B(n_1058), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1069), .B(n_1071), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1059), .B(n_1063), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_1053), .A2(n_1095), .B1(n_1099), .B2(n_1047), .Y(n_1148) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_1068), .B(n_1041), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1039), .B(n_1065), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1060), .B(n_1039), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1065), .B(n_1097), .Y(n_1152) );
NAND2xp5_ASAP7_75t_SL g1153 ( .A(n_1083), .B(n_1096), .Y(n_1153) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1050), .Y(n_1154) );
XNOR2x1_ASAP7_75t_L g1155 ( .A(n_1079), .B(n_1091), .Y(n_1155) );
NAND2xp5_ASAP7_75t_SL g1156 ( .A(n_1096), .B(n_1089), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1051), .B(n_1066), .Y(n_1157) );
NAND3xp33_ASAP7_75t_L g1158 ( .A(n_1092), .B(n_1103), .C(n_1107), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1094), .B(n_1100), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1110), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_1159), .B(n_1094), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1111), .Y(n_1162) );
XNOR2xp5_ASAP7_75t_L g1163 ( .A(n_1155), .B(n_1079), .Y(n_1163) );
INVx1_ASAP7_75t_SL g1164 ( .A(n_1155), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1152), .B(n_1072), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1126), .Y(n_1166) );
INVx2_ASAP7_75t_SL g1167 ( .A(n_1124), .Y(n_1167) );
INVx2_ASAP7_75t_SL g1168 ( .A(n_1124), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_1139), .B(n_1086), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1127), .Y(n_1170) );
AND3x2_ASAP7_75t_L g1171 ( .A(n_1114), .B(n_1096), .C(n_1095), .Y(n_1171) );
NAND3xp33_ASAP7_75t_SL g1172 ( .A(n_1143), .B(n_1099), .C(n_1103), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1139), .B(n_1072), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1144), .B(n_1072), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1157), .B(n_1098), .Y(n_1175) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1150), .B(n_1107), .Y(n_1176) );
AOI221xp5_ASAP7_75t_L g1177 ( .A1(n_1141), .A2(n_1076), .B1(n_1105), .B2(n_1091), .C(n_1090), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1136), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1137), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1149), .B(n_1087), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1150), .B(n_1105), .Y(n_1181) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1154), .Y(n_1182) );
NAND3xp33_ASAP7_75t_L g1183 ( .A(n_1122), .B(n_1106), .C(n_1104), .Y(n_1183) );
NOR4xp25_ASAP7_75t_L g1184 ( .A(n_1148), .B(n_1074), .C(n_1104), .D(n_1106), .Y(n_1184) );
AND2x4_ASAP7_75t_L g1185 ( .A(n_1156), .B(n_1040), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1146), .B(n_1088), .Y(n_1186) );
INVx3_ASAP7_75t_L g1187 ( .A(n_1123), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1151), .B(n_1088), .Y(n_1188) );
AND2x4_ASAP7_75t_L g1189 ( .A(n_1156), .B(n_1040), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1113), .B(n_1087), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1138), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1113), .B(n_1093), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1145), .B(n_1093), .Y(n_1193) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1123), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_1112), .A2(n_1096), .B1(n_1081), .B2(n_1078), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1160), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1160), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1162), .Y(n_1198) );
AND2x4_ASAP7_75t_L g1199 ( .A(n_1185), .B(n_1153), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1162), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1165), .B(n_1120), .Y(n_1201) );
NOR2xp33_ASAP7_75t_L g1202 ( .A(n_1164), .B(n_1132), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1176), .B(n_1142), .Y(n_1203) );
INVxp67_ASAP7_75t_L g1204 ( .A(n_1167), .Y(n_1204) );
AOI22xp5_ASAP7_75t_L g1205 ( .A1(n_1172), .A2(n_1177), .B1(n_1119), .B2(n_1171), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1181), .B(n_1140), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1175), .B(n_1147), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1165), .B(n_1120), .Y(n_1208) );
AOI21xp5_ASAP7_75t_L g1209 ( .A1(n_1184), .A2(n_1153), .B(n_1125), .Y(n_1209) );
O2A1O1Ixp5_ASAP7_75t_L g1210 ( .A1(n_1185), .A2(n_1116), .B(n_1117), .C(n_1158), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1169), .B(n_1135), .Y(n_1211) );
INVxp67_ASAP7_75t_L g1212 ( .A(n_1167), .Y(n_1212) );
XNOR2x1_ASAP7_75t_L g1213 ( .A(n_1163), .B(n_1128), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1166), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1161), .B(n_1135), .Y(n_1215) );
XOR2xp5_ASAP7_75t_L g1216 ( .A(n_1163), .B(n_1133), .Y(n_1216) );
XOR2x2_ASAP7_75t_L g1217 ( .A(n_1192), .B(n_1116), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1170), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1170), .Y(n_1219) );
OAI31xp33_ASAP7_75t_L g1220 ( .A1(n_1183), .A2(n_1118), .A3(n_1121), .B(n_1130), .Y(n_1220) );
NAND4xp25_ASAP7_75t_L g1221 ( .A(n_1195), .B(n_1118), .C(n_1131), .D(n_1134), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1178), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1161), .B(n_1129), .Y(n_1223) );
O2A1O1Ixp33_ASAP7_75t_L g1224 ( .A1(n_1168), .A2(n_1115), .B(n_1082), .C(n_1073), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1179), .Y(n_1225) );
XNOR2xp5_ASAP7_75t_L g1226 ( .A(n_1192), .B(n_1067), .Y(n_1226) );
INVx2_ASAP7_75t_SL g1227 ( .A(n_1187), .Y(n_1227) );
AOI221xp5_ASAP7_75t_L g1228 ( .A1(n_1179), .A2(n_1073), .B1(n_1191), .B2(n_1193), .C(n_1173), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1173), .B(n_1174), .Y(n_1229) );
INVxp67_ASAP7_75t_L g1230 ( .A(n_1188), .Y(n_1230) );
INVxp33_ASAP7_75t_SL g1231 ( .A(n_1202), .Y(n_1231) );
OAI22xp33_ASAP7_75t_L g1232 ( .A1(n_1205), .A2(n_1221), .B1(n_1209), .B2(n_1204), .Y(n_1232) );
AOI21xp5_ASAP7_75t_L g1233 ( .A1(n_1213), .A2(n_1217), .B(n_1220), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1228), .B(n_1211), .Y(n_1234) );
AOI21xp33_ASAP7_75t_L g1235 ( .A1(n_1224), .A2(n_1210), .B(n_1216), .Y(n_1235) );
AOI22xp5_ASAP7_75t_SL g1236 ( .A1(n_1216), .A2(n_1226), .B1(n_1212), .B2(n_1230), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1215), .B(n_1217), .Y(n_1237) );
AOI22xp5_ASAP7_75t_L g1238 ( .A1(n_1199), .A2(n_1201), .B1(n_1208), .B2(n_1226), .Y(n_1238) );
AOI21xp5_ASAP7_75t_L g1239 ( .A1(n_1223), .A2(n_1227), .B(n_1199), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1203), .B(n_1206), .Y(n_1240) );
NOR2x1_ASAP7_75t_L g1241 ( .A(n_1232), .B(n_1199), .Y(n_1241) );
XNOR2xp5_ASAP7_75t_L g1242 ( .A(n_1236), .B(n_1207), .Y(n_1242) );
AOI22xp5_ASAP7_75t_SL g1243 ( .A1(n_1233), .A2(n_1189), .B1(n_1229), .B2(n_1227), .Y(n_1243) );
NAND4xp25_ASAP7_75t_L g1244 ( .A(n_1235), .B(n_1189), .C(n_1174), .D(n_1190), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1234), .B(n_1225), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1240), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1237), .B(n_1197), .Y(n_1247) );
AND2x4_ASAP7_75t_L g1248 ( .A(n_1246), .B(n_1239), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1245), .Y(n_1249) );
NAND4xp25_ASAP7_75t_L g1250 ( .A(n_1241), .B(n_1231), .C(n_1238), .D(n_1189), .Y(n_1250) );
NAND3xp33_ASAP7_75t_SL g1251 ( .A(n_1243), .B(n_1219), .C(n_1198), .Y(n_1251) );
NOR2x1p5_ASAP7_75t_L g1252 ( .A(n_1244), .B(n_1218), .Y(n_1252) );
NOR4xp25_ASAP7_75t_L g1253 ( .A(n_1250), .B(n_1247), .C(n_1242), .D(n_1222), .Y(n_1253) );
OAI22xp5_ASAP7_75t_L g1254 ( .A1(n_1252), .A2(n_1214), .B1(n_1196), .B2(n_1200), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1249), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1255), .Y(n_1256) );
OR3x1_ASAP7_75t_L g1257 ( .A(n_1253), .B(n_1251), .C(n_1248), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1254), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1256), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1258), .B(n_1190), .Y(n_1260) );
AOI21xp33_ASAP7_75t_SL g1261 ( .A1(n_1259), .A2(n_1257), .B(n_1180), .Y(n_1261) );
XNOR2xp5_ASAP7_75t_L g1262 ( .A(n_1260), .B(n_1257), .Y(n_1262) );
OAI31xp33_ASAP7_75t_L g1263 ( .A1(n_1262), .A2(n_1193), .A3(n_1186), .B(n_1194), .Y(n_1263) );
O2A1O1Ixp33_ASAP7_75t_L g1264 ( .A1(n_1263), .A2(n_1182), .B(n_1186), .C(n_1261), .Y(n_1264) );
endmodule