module fake_netlist_6_2859_n_1999 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1999);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1999;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_850;
wire n_690;
wire n_1886;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_145),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_147),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_29),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_55),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_17),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_63),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_180),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_85),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_47),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_12),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_199),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_43),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_18),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_18),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_74),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_166),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_91),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_95),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_65),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_72),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_59),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_137),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_40),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_57),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_171),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_44),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_44),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_114),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_115),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_200),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_161),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_41),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_80),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_126),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_128),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_69),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_73),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_61),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_158),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_109),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_172),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_136),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_96),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_54),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_194),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_174),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_150),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_117),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_185),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_50),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_21),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_132),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_101),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_135),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_197),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_40),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_84),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_157),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_50),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_100),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_204),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_8),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_1),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_38),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_2),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_59),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_167),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_62),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_71),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_202),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_144),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_83),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_24),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_183),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_121),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_148),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_175),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_151),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_107),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_43),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_75),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_159),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_26),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_98),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_37),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_14),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_82),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_203),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_76),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_116),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_165),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_118),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_39),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_112),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_48),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_113),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_169),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_97),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_49),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_92),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_10),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_51),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_170),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_5),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_26),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_53),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_81),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_47),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_106),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_28),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_102),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_8),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_37),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_41),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_68),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g329 ( 
.A(n_46),
.Y(n_329)
);

BUFx2_ASAP7_75t_SL g330 ( 
.A(n_52),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_162),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_54),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_20),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_57),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_49),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_52),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_142),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_138),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_45),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_87),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_35),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_154),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_20),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_108),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_39),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_173),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_13),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_181),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_168),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_104),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_2),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_149),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_58),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_64),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_205),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_120),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_55),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_68),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_156),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_193),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_9),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_23),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_67),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_79),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_64),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_179),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_99),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_70),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_9),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_53),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_7),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_62),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_89),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_36),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_25),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_0),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_34),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_133),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_111),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_69),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_7),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_143),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_103),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_127),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_124),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_14),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_35),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_45),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_123),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_34),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_28),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_21),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_29),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_10),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_12),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_19),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_94),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_24),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_131),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_23),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_17),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_19),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_146),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_22),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_31),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_176),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_71),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_48),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_51),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_206),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_0),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_272),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_244),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_334),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_266),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_257),
.B(n_1),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_301),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_207),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_211),
.B(n_3),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_334),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_213),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_272),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_214),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_217),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_334),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_408),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_305),
.B(n_259),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_216),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_221),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_316),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_216),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_223),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_224),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_220),
.B(n_3),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_225),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_228),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_229),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_233),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_305),
.B(n_4),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_368),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_271),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_210),
.B(n_4),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_208),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_271),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_259),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g457 ( 
.A(n_209),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_381),
.B(n_5),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_231),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_242),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_243),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_259),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_212),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_231),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_269),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_304),
.B(n_237),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_246),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_247),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_269),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_248),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_254),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_255),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_256),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_258),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_279),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_260),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_279),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_261),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_304),
.B(n_237),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_293),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_262),
.Y(n_481)
);

INVxp33_ASAP7_75t_SL g482 ( 
.A(n_215),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_268),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_210),
.B(n_6),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_236),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_293),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_296),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_218),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_219),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_296),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_270),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_274),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_280),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_283),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_327),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_327),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_284),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_222),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_333),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_304),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_287),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_227),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_333),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_R g504 ( 
.A(n_289),
.B(n_6),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_335),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_335),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_252),
.B(n_11),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_336),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_290),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_336),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_294),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_485),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_485),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_414),
.A2(n_263),
.B1(n_319),
.B2(n_245),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_462),
.B(n_295),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_410),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_415),
.B(n_421),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_485),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_485),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_415),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_458),
.B(n_226),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_421),
.B(n_427),
.Y(n_525)
);

BUFx8_ASAP7_75t_L g526 ( 
.A(n_458),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_427),
.B(n_252),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_456),
.B(n_226),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_430),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_455),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_500),
.B(n_300),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_422),
.B(n_355),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_422),
.B(n_355),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_485),
.B(n_230),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_428),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_466),
.B(n_230),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_454),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_431),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_456),
.B(n_232),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_434),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_434),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_459),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_459),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_464),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_507),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_464),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_465),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g551 ( 
.A(n_449),
.B(n_236),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_479),
.B(n_232),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_469),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_469),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_475),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_475),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_477),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_480),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_463),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_435),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_480),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_486),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_453),
.B(n_238),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_486),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_487),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_429),
.B(n_236),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_487),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_490),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_490),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_435),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_484),
.B(n_238),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_495),
.B(n_241),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_495),
.Y(n_574)
);

OA21x2_ASAP7_75t_L g575 ( 
.A1(n_496),
.A2(n_343),
.B(n_339),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_496),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_499),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_499),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_503),
.B(n_241),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_505),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_505),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_420),
.B(n_253),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_506),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_437),
.B(n_442),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_437),
.B(n_250),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_413),
.A2(n_386),
.B1(n_341),
.B2(n_345),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_506),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_508),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_510),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_510),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_442),
.B(n_302),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_447),
.B(n_250),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_524),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_547),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_547),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_533),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_553),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_547),
.B(n_236),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_520),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_583),
.B(n_428),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_561),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_533),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_561),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_528),
.B(n_447),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_583),
.B(n_411),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_517),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_564),
.A2(n_443),
.B1(n_439),
.B2(n_436),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_533),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_547),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_520),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_547),
.B(n_515),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_547),
.B(n_236),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_547),
.B(n_419),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_533),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_512),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_517),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_547),
.B(n_236),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_514),
.B(n_416),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_533),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_520),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_561),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_515),
.B(n_457),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_561),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_532),
.B(n_482),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_516),
.B(n_450),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_518),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_536),
.B(n_423),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_564),
.A2(n_572),
.B1(n_524),
.B2(n_552),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_572),
.A2(n_524),
.B1(n_552),
.B2(n_526),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_547),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_553),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_520),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_532),
.B(n_498),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_528),
.B(n_541),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_571),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_571),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_571),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_571),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_524),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_575),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_553),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_538),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_538),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_553),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_520),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_552),
.B(n_425),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_553),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_587),
.A2(n_417),
.B1(n_504),
.B2(n_412),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_553),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_572),
.B(n_426),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_520),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_552),
.B(n_432),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_536),
.B(n_438),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_553),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_575),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_552),
.B(n_440),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_552),
.A2(n_424),
.B1(n_299),
.B2(n_312),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_560),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_553),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_575),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_520),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_516),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_557),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_526),
.A2(n_299),
.B1(n_312),
.B2(n_281),
.Y(n_667)
);

XNOR2xp5_ASAP7_75t_L g668 ( 
.A(n_514),
.B(n_418),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_560),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_567),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_520),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_575),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_575),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_593),
.B(n_444),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_567),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_518),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_575),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_575),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_593),
.B(n_445),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_523),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_535),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_528),
.B(n_451),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_551),
.B(n_446),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_535),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_523),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_535),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_551),
.B(n_448),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_536),
.B(n_460),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_535),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_557),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_557),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_523),
.Y(n_692)
);

INVx6_ASAP7_75t_L g693 ( 
.A(n_526),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_529),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_537),
.B(n_461),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_535),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_551),
.B(n_467),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_SL g698 ( 
.A(n_587),
.B(n_478),
.C(n_472),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_529),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_529),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_530),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_530),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_567),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_526),
.A2(n_281),
.B1(n_489),
.B2(n_502),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_535),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_526),
.A2(n_489),
.B1(n_502),
.B2(n_351),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_520),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_537),
.A2(n_483),
.B1(n_501),
.B2(n_481),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_585),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_537),
.B(n_468),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_512),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_528),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_521),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_585),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_530),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_585),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_541),
.B(n_451),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_551),
.B(n_470),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_567),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_521),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_585),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_512),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_541),
.B(n_586),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_551),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_544),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_526),
.B(n_471),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_557),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_541),
.B(n_473),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_557),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_544),
.Y(n_730)
);

BUFx4f_ASAP7_75t_L g731 ( 
.A(n_567),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_521),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_587),
.B(n_474),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_514),
.A2(n_450),
.B1(n_433),
.B2(n_330),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_512),
.Y(n_735)
);

BUFx4f_ASAP7_75t_L g736 ( 
.A(n_567),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_586),
.B(n_476),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_539),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_SL g739 ( 
.A(n_531),
.B(n_491),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_573),
.B(n_330),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_544),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_551),
.A2(n_332),
.B1(n_398),
.B2(n_275),
.Y(n_742)
);

BUFx4f_ASAP7_75t_L g743 ( 
.A(n_567),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_653),
.B(n_551),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_695),
.B(n_493),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_631),
.A2(n_551),
.B1(n_567),
.B2(n_586),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_601),
.B(n_494),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_710),
.B(n_497),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_709),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_679),
.B(n_551),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_738),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_601),
.B(n_509),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_709),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_595),
.B(n_642),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_714),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_714),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_738),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_698),
.B(n_579),
.C(n_573),
.Y(n_758)
);

INVx8_ASAP7_75t_L g759 ( 
.A(n_740),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_609),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_645),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_625),
.B(n_511),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_595),
.B(n_551),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_601),
.B(n_406),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_620),
.A2(n_551),
.B1(n_567),
.B2(n_586),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_627),
.B(n_492),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_636),
.B(n_488),
.Y(n_767)
);

OR2x6_ASAP7_75t_L g768 ( 
.A(n_720),
.B(n_531),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_642),
.B(n_551),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_620),
.B(n_406),
.Y(n_770)
);

BUFx2_ASAP7_75t_SL g771 ( 
.A(n_645),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_712),
.B(n_562),
.Y(n_772)
);

BUFx6f_ASAP7_75t_SL g773 ( 
.A(n_661),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_610),
.B(n_594),
.C(n_235),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_712),
.B(n_562),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_728),
.B(n_273),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_649),
.B(n_366),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_665),
.Y(n_778)
);

AOI221xp5_ASAP7_75t_L g779 ( 
.A1(n_733),
.A2(n_343),
.B1(n_351),
.B2(n_357),
.C(n_339),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_655),
.B(n_379),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_620),
.A2(n_567),
.B1(n_594),
.B2(n_370),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_665),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_716),
.B(n_594),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_659),
.B(n_303),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_696),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_619),
.Y(n_786)
);

AND2x6_ASAP7_75t_L g787 ( 
.A(n_643),
.B(n_658),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_737),
.A2(n_567),
.B1(n_320),
.B2(n_324),
.Y(n_788)
);

O2A1O1Ixp5_ASAP7_75t_L g789 ( 
.A1(n_643),
.A2(n_527),
.B(n_534),
.C(n_562),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_674),
.B(n_562),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_L g791 ( 
.A(n_632),
.B(n_567),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_669),
.B(n_531),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_658),
.A2(n_573),
.B(n_579),
.C(n_527),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_614),
.B(n_562),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_723),
.B(n_562),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_713),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_716),
.A2(n_267),
.B1(n_285),
.B2(n_265),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_721),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_SL g799 ( 
.A(n_706),
.B(n_239),
.C(n_234),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_721),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_598),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_704),
.B(n_313),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_669),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_598),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_651),
.B(n_337),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_663),
.A2(n_579),
.B(n_527),
.C(n_534),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_663),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_732),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_723),
.B(n_578),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_731),
.B(n_406),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_637),
.B(n_578),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_651),
.B(n_342),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_672),
.A2(n_370),
.B1(n_387),
.B2(n_393),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_696),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_637),
.B(n_578),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_616),
.B(n_578),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_605),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_608),
.A2(n_344),
.B1(n_346),
.B2(n_348),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_725),
.B(n_578),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_628),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_646),
.B(n_329),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_607),
.B(n_548),
.Y(n_822)
);

AND2x6_ASAP7_75t_L g823 ( 
.A(n_672),
.B(n_265),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_708),
.B(n_350),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_667),
.B(n_352),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_L g826 ( 
.A(n_683),
.B(n_356),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_730),
.B(n_588),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_734),
.B(n_603),
.C(n_630),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_730),
.B(n_588),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_656),
.B(n_285),
.C(n_267),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_741),
.B(n_588),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_739),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_L g833 ( 
.A(n_697),
.B(n_360),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_726),
.B(n_548),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_741),
.B(n_588),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_607),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_742),
.B(n_367),
.Y(n_837)
);

BUFx12f_ASAP7_75t_L g838 ( 
.A(n_720),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_742),
.B(n_633),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_682),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_611),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_681),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_624),
.B(n_588),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_740),
.B(n_588),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_731),
.B(n_736),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_660),
.B(n_740),
.C(n_717),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_629),
.Y(n_847)
);

O2A1O1Ixp5_ASAP7_75t_L g848 ( 
.A1(n_673),
.A2(n_534),
.B(n_590),
.C(n_592),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_676),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_731),
.B(n_406),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_731),
.B(n_406),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_676),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_633),
.B(n_736),
.Y(n_853)
);

AND2x6_ASAP7_75t_L g854 ( 
.A(n_673),
.B(n_288),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_696),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_740),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_604),
.Y(n_857)
);

BUFx5_ASAP7_75t_L g858 ( 
.A(n_633),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_677),
.A2(n_407),
.B1(n_387),
.B2(n_338),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_604),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_633),
.B(n_373),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_624),
.B(n_590),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_611),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_736),
.B(n_385),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_677),
.A2(n_383),
.B1(n_291),
.B2(n_384),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_740),
.B(n_590),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_688),
.B(n_590),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_680),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_621),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_682),
.B(n_590),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_626),
.B(n_590),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_680),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_626),
.B(n_638),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_617),
.Y(n_874)
);

INVx5_ASAP7_75t_L g875 ( 
.A(n_615),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_638),
.B(n_592),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_622),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_717),
.B(n_329),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_685),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_736),
.B(n_389),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_681),
.A2(n_403),
.B1(n_399),
.B2(n_397),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_L g882 ( 
.A(n_718),
.B(n_292),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_743),
.B(n_557),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_639),
.B(n_592),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_L g885 ( 
.A(n_684),
.B(n_307),
.C(n_297),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_685),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_639),
.B(n_592),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_640),
.B(n_592),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_604),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_692),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_606),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_606),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_640),
.B(n_592),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_641),
.B(n_329),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_711),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_606),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_692),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_641),
.B(n_557),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_596),
.B(n_557),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_711),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_762),
.B(n_596),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_858),
.B(n_743),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_767),
.B(n_596),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_758),
.A2(n_678),
.B(n_687),
.C(n_686),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_801),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_780),
.B(n_597),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_767),
.A2(n_686),
.B1(n_689),
.B2(n_684),
.Y(n_907)
);

AOI21xp33_ASAP7_75t_L g908 ( 
.A1(n_766),
.A2(n_668),
.B(n_689),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_845),
.A2(n_612),
.B(n_597),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_845),
.A2(n_612),
.B(n_597),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_778),
.Y(n_911)
);

INVx5_ASAP7_75t_L g912 ( 
.A(n_787),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_853),
.A2(n_612),
.B(n_743),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_780),
.B(n_612),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_754),
.B(n_678),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_804),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_858),
.B(n_743),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_858),
.B(n_875),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_758),
.A2(n_705),
.B(n_699),
.C(n_700),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_790),
.B(n_705),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_860),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_858),
.B(n_724),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_771),
.B(n_621),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_794),
.A2(n_675),
.B(n_670),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_790),
.B(n_807),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_867),
.A2(n_735),
.B(n_618),
.C(n_722),
.Y(n_926)
);

NOR2x2_ASAP7_75t_L g927 ( 
.A(n_768),
.B(n_799),
.Y(n_927)
);

NOR2x1_ASAP7_75t_L g928 ( 
.A(n_846),
.B(n_670),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_807),
.B(n_749),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_785),
.Y(n_930)
);

AO21x1_ASAP7_75t_L g931 ( 
.A1(n_764),
.A2(n_307),
.B(n_297),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_867),
.A2(n_675),
.B1(n_670),
.B2(n_703),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_817),
.Y(n_933)
);

BUFx8_ASAP7_75t_SL g934 ( 
.A(n_838),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_816),
.A2(n_899),
.B(n_857),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_857),
.A2(n_675),
.B(n_670),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_753),
.B(n_711),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_900),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_789),
.A2(n_703),
.B(n_675),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_865),
.A2(n_615),
.B1(n_382),
.B2(n_384),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_900),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_755),
.B(n_711),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_883),
.A2(n_719),
.B(n_703),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_756),
.B(n_722),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_883),
.A2(n_719),
.B(n_703),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_865),
.A2(n_615),
.B1(n_383),
.B2(n_378),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_811),
.A2(n_719),
.B(n_613),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_860),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_858),
.B(n_724),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_798),
.B(n_722),
.Y(n_950)
);

NOR2x1_ASAP7_75t_L g951 ( 
.A(n_745),
.B(n_719),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_800),
.B(n_783),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_815),
.A2(n_613),
.B(n_724),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_795),
.A2(n_613),
.B(n_724),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_809),
.A2(n_613),
.B(n_602),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_783),
.B(n_822),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_841),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_785),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_822),
.B(n_722),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_803),
.B(n_329),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_870),
.B(n_694),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_870),
.B(n_694),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_836),
.B(n_699),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_808),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_840),
.B(n_548),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_785),
.B(n_554),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_750),
.A2(n_613),
.B(n_602),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_859),
.A2(n_615),
.B1(n_382),
.B2(n_378),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_863),
.B(n_700),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_782),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_874),
.B(n_877),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_781),
.B(n_701),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_781),
.B(n_859),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_792),
.B(n_554),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_858),
.B(n_613),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_787),
.B(n_701),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_768),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_760),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_791),
.A2(n_623),
.B(n_602),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_875),
.B(n_599),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_787),
.B(n_702),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_763),
.A2(n_769),
.B(n_839),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_787),
.B(n_702),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_787),
.B(n_715),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_747),
.A2(n_715),
.B(n_310),
.C(n_309),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_748),
.B(n_602),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_761),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_744),
.A2(n_775),
.B(n_772),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_746),
.A2(n_693),
.B1(n_349),
.B2(n_364),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_875),
.A2(n_635),
.B(n_623),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_848),
.A2(n_615),
.B(n_729),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_796),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_894),
.B(n_623),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_768),
.Y(n_994)
);

NOR2x1_ASAP7_75t_L g995 ( 
.A(n_747),
.B(n_309),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_813),
.A2(n_310),
.B(n_311),
.C(n_322),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_806),
.A2(n_615),
.B(n_729),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_878),
.B(n_623),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_813),
.B(n_635),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_832),
.B(n_599),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_860),
.B(n_889),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_844),
.A2(n_311),
.B(n_322),
.C(n_331),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_875),
.A2(n_648),
.B(n_635),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_873),
.A2(n_746),
.B(n_765),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_860),
.B(n_635),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_785),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_765),
.A2(n_693),
.B1(n_338),
.B2(n_340),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_820),
.B(n_766),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_821),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_805),
.B(n_648),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_793),
.A2(n_770),
.B(n_764),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_814),
.B(n_599),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_812),
.B(n_648),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_L g1014 ( 
.A(n_759),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_864),
.A2(n_664),
.B(n_654),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_880),
.A2(n_664),
.B(n_654),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_814),
.B(n_855),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_776),
.B(n_554),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_889),
.B(n_654),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_814),
.B(n_556),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_891),
.B(n_664),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_777),
.B(n_830),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_856),
.Y(n_1023)
);

OAI321xp33_ASAP7_75t_L g1024 ( 
.A1(n_779),
.A2(n_349),
.A3(n_331),
.B1(n_340),
.B2(n_359),
.C(n_364),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_786),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_843),
.A2(n_871),
.B(n_862),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_752),
.A2(n_359),
.B(n_574),
.C(n_565),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_891),
.B(n_664),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_876),
.A2(n_888),
.B(n_833),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_856),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_752),
.A2(n_574),
.B(n_580),
.C(n_576),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_844),
.A2(n_729),
.B(n_727),
.C(n_600),
.Y(n_1032)
);

AO21x1_ASAP7_75t_L g1033 ( 
.A1(n_770),
.A2(n_634),
.B(n_600),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_826),
.A2(n_850),
.B(n_810),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_891),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_810),
.A2(n_707),
.B(n_671),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_774),
.B(n_671),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_850),
.A2(n_707),
.B(n_671),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_851),
.A2(n_707),
.B(n_671),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_814),
.B(n_600),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_866),
.A2(n_727),
.B(n_634),
.C(n_691),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_891),
.B(n_707),
.Y(n_1042)
);

OAI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_828),
.A2(n_249),
.B(n_240),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_851),
.A2(n_882),
.B(n_895),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_855),
.B(n_634),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_855),
.Y(n_1046)
);

O2A1O1Ixp5_ASAP7_75t_L g1047 ( 
.A1(n_884),
.A2(n_727),
.B(n_644),
.C(n_691),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_824),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_847),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_855),
.B(n_556),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_898),
.A2(n_647),
.B(n_644),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_861),
.A2(n_647),
.B(n_644),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_819),
.A2(n_650),
.B(n_647),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_892),
.B(n_615),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_869),
.B(n_828),
.Y(n_1055)
);

BUFx4f_ASAP7_75t_L g1056 ( 
.A(n_759),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_892),
.Y(n_1057)
);

AND2x2_ASAP7_75t_SL g1058 ( 
.A(n_885),
.B(n_830),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_834),
.B(n_650),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_892),
.B(n_652),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_892),
.B(n_652),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_896),
.B(n_657),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_773),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_SL g1064 ( 
.A(n_773),
.B(n_693),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_827),
.A2(n_662),
.B(n_657),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_866),
.A2(n_662),
.B(n_657),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_896),
.A2(n_693),
.B1(n_759),
.B2(n_784),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_797),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_837),
.A2(n_842),
.B(n_885),
.C(n_802),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_849),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_829),
.A2(n_666),
.B(n_662),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_896),
.B(n_666),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_896),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_831),
.A2(n_563),
.B(n_570),
.C(n_574),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_825),
.B(n_556),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_884),
.B(n_666),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_975),
.A2(n_835),
.B(n_852),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_902),
.A2(n_893),
.B(n_887),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_903),
.A2(n_881),
.B1(n_788),
.B2(n_818),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_903),
.B(n_823),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_930),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_905),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_916),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_911),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_973),
.A2(n_946),
.B1(n_940),
.B2(n_968),
.Y(n_1085)
);

NAND2xp33_ASAP7_75t_SL g1086 ( 
.A(n_1022),
.B(n_868),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_933),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_1069),
.A2(n_893),
.B(n_887),
.C(n_890),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_902),
.A2(n_879),
.B(n_872),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_SL g1090 ( 
.A(n_908),
.B(n_264),
.C(n_251),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_957),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_977),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_996),
.A2(n_886),
.B(n_897),
.C(n_751),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_L g1094 ( 
.A(n_964),
.B(n_757),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1048),
.A2(n_854),
.B1(n_823),
.B2(n_691),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1068),
.A2(n_565),
.B(n_558),
.C(n_580),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_917),
.A2(n_690),
.B(n_522),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1008),
.B(n_823),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_917),
.A2(n_690),
.B(n_522),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_967),
.A2(n_690),
.B(n_525),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_940),
.A2(n_558),
.B1(n_563),
.B2(n_565),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_925),
.B(n_823),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_934),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_974),
.B(n_823),
.Y(n_1104)
);

NOR3xp33_ASAP7_75t_SL g1105 ( 
.A(n_1043),
.B(n_277),
.C(n_276),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_SL g1106 ( 
.A(n_1024),
.B(n_317),
.C(n_278),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1011),
.A2(n_568),
.B(n_580),
.C(n_576),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_930),
.Y(n_1108)
);

O2A1O1Ixp5_ASAP7_75t_SL g1109 ( 
.A1(n_1059),
.A2(n_558),
.B(n_576),
.C(n_570),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_1068),
.A2(n_563),
.B(n_568),
.C(n_570),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_965),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_L g1112 ( 
.A(n_1055),
.B(n_314),
.C(n_318),
.Y(n_1112)
);

BUFx4f_ASAP7_75t_L g1113 ( 
.A(n_930),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_964),
.B(n_1009),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1002),
.A2(n_568),
.B(n_591),
.C(n_589),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1004),
.B(n_854),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_911),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_992),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_956),
.A2(n_854),
.B1(n_253),
.B2(n_540),
.Y(n_1119)
);

OAI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_960),
.A2(n_306),
.B(n_308),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_901),
.B(n_854),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_996),
.A2(n_549),
.B(n_591),
.C(n_589),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_978),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_912),
.B(n_253),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_922),
.A2(n_512),
.B(n_522),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1037),
.A2(n_854),
.B(n_540),
.C(n_298),
.Y(n_1126)
);

OAI21xp33_ASAP7_75t_SL g1127 ( 
.A1(n_946),
.A2(n_519),
.B(n_525),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_963),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_922),
.A2(n_512),
.B(n_522),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_961),
.B(n_557),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_962),
.B(n_545),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_923),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_952),
.Y(n_1133)
);

NAND2x1p5_ASAP7_75t_L g1134 ( 
.A(n_912),
.B(n_958),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_920),
.B(n_545),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_949),
.A2(n_522),
.B(n_513),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_1063),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_970),
.B(n_282),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_929),
.B(n_545),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_971),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1037),
.A2(n_396),
.B(n_315),
.C(n_321),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1018),
.B(n_286),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1023),
.B(n_323),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1058),
.A2(n_995),
.B1(n_1020),
.B2(n_966),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_912),
.B(n_253),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_930),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_968),
.A2(n_401),
.B1(n_326),
.B2(n_328),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1058),
.A2(n_928),
.B1(n_1020),
.B2(n_966),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1030),
.B(n_325),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_904),
.A2(n_404),
.B(n_353),
.C(n_354),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1023),
.B(n_347),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_906),
.B(n_546),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_987),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_914),
.B(n_546),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1050),
.A2(n_591),
.B1(n_589),
.B2(n_584),
.Y(n_1155)
);

AO22x1_ASAP7_75t_L g1156 ( 
.A1(n_994),
.A2(n_400),
.B1(n_361),
.B2(n_362),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_949),
.A2(n_522),
.B(n_513),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1006),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_958),
.B(n_546),
.Y(n_1159)
);

INVx6_ASAP7_75t_L g1160 ( 
.A(n_1006),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1050),
.B(n_549),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1063),
.B(n_358),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_907),
.B(n_549),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_915),
.B(n_549),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_998),
.B(n_550),
.Y(n_1165)
);

OAI21xp33_ASAP7_75t_L g1166 ( 
.A1(n_1075),
.A2(n_365),
.B(n_369),
.Y(n_1166)
);

AOI21x1_ASAP7_75t_L g1167 ( 
.A1(n_975),
.A2(n_519),
.B(n_525),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1000),
.B(n_550),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1032),
.A2(n_591),
.B(n_589),
.C(n_584),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_918),
.A2(n_513),
.B(n_519),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1010),
.A2(n_409),
.B(n_375),
.C(n_376),
.Y(n_1171)
);

O2A1O1Ixp5_ASAP7_75t_L g1172 ( 
.A1(n_1034),
.A2(n_584),
.B(n_582),
.C(n_581),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_993),
.B(n_550),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1014),
.B(n_371),
.Y(n_1174)
);

O2A1O1Ixp5_ASAP7_75t_L g1175 ( 
.A1(n_931),
.A2(n_1033),
.B(n_997),
.C(n_1029),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_972),
.A2(n_377),
.B1(n_380),
.B2(n_388),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1010),
.A2(n_390),
.B(n_391),
.C(n_392),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_988),
.B(n_550),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_989),
.A2(n_394),
.B1(n_395),
.B2(n_402),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_918),
.A2(n_513),
.B(n_582),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1014),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_959),
.B(n_405),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_936),
.A2(n_584),
.B(n_582),
.Y(n_1183)
);

OR2x2_ASAP7_75t_SL g1184 ( 
.A(n_927),
.B(n_555),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_913),
.A2(n_582),
.B(n_581),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1006),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1006),
.Y(n_1187)
);

INVx8_ASAP7_75t_L g1188 ( 
.A(n_1057),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_982),
.B(n_581),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_999),
.A2(n_581),
.B1(n_577),
.B2(n_569),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_909),
.A2(n_577),
.B(n_569),
.Y(n_1191)
);

NAND2xp33_ASAP7_75t_L g1192 ( 
.A(n_1057),
.B(n_577),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_969),
.B(n_577),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_938),
.B(n_11),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1064),
.B(n_569),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1007),
.A2(n_569),
.B1(n_566),
.B2(n_559),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1057),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1056),
.B(n_566),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_L g1199 ( 
.A(n_1025),
.B(n_105),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_932),
.A2(n_566),
.B1(n_559),
.B2(n_555),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_941),
.B(n_566),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_986),
.B(n_13),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1049),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1076),
.B(n_559),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1056),
.A2(n_559),
.B1(n_555),
.B2(n_543),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1046),
.B(n_555),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1041),
.A2(n_543),
.B(n_542),
.C(n_539),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1057),
.Y(n_1208)
);

AND2x2_ASAP7_75t_SL g1209 ( 
.A(n_1046),
.B(n_543),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_910),
.A2(n_543),
.B(n_542),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1070),
.A2(n_539),
.B1(n_542),
.B2(n_22),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_921),
.Y(n_1212)
);

NAND3xp33_ASAP7_75t_SL g1213 ( 
.A(n_985),
.B(n_542),
.C(n_539),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1001),
.B(n_15),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_924),
.A2(n_90),
.B(n_198),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_976),
.B(n_15),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_921),
.B(n_16),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_981),
.A2(n_16),
.B1(n_25),
.B2(n_27),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_983),
.B(n_984),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_948),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1035),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_SL g1222 ( 
.A(n_1035),
.B(n_27),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_919),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1088),
.A2(n_1013),
.A3(n_935),
.B(n_926),
.Y(n_1224)
);

AOI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1176),
.A2(n_1027),
.B1(n_1031),
.B2(n_1074),
.C(n_1013),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1087),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1113),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1121),
.A2(n_939),
.B(n_954),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1079),
.A2(n_1044),
.B(n_951),
.C(n_1026),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1100),
.A2(n_1051),
.B(n_1052),
.Y(n_1230)
);

AOI221xp5_ASAP7_75t_L g1231 ( 
.A1(n_1176),
.A2(n_1067),
.B1(n_942),
.B2(n_937),
.C(n_950),
.Y(n_1231)
);

AO22x2_ASAP7_75t_L g1232 ( 
.A1(n_1218),
.A2(n_1017),
.B1(n_1066),
.B2(n_1059),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1118),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1191),
.A2(n_955),
.B(n_1015),
.Y(n_1234)
);

CKINVDCx6p67_ASAP7_75t_R g1235 ( 
.A(n_1103),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1133),
.B(n_1073),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1128),
.B(n_944),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1111),
.B(n_1017),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1117),
.B(n_1060),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1142),
.B(n_1061),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1178),
.A2(n_953),
.B(n_945),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_SL g1242 ( 
.A1(n_1150),
.A2(n_1126),
.B(n_1080),
.C(n_1116),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1185),
.A2(n_1016),
.B(n_1047),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1175),
.A2(n_1047),
.B(n_991),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_1112),
.B(n_1062),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1172),
.A2(n_1071),
.B(n_1065),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1182),
.B(n_1072),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1152),
.A2(n_1154),
.B(n_1078),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1116),
.A2(n_979),
.B(n_1053),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1098),
.A2(n_1054),
.B(n_1036),
.C(n_1038),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1181),
.B(n_1045),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1219),
.B(n_1005),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1107),
.A2(n_1039),
.B(n_1040),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1092),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1210),
.A2(n_947),
.B(n_1012),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1102),
.A2(n_943),
.B(n_1042),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1132),
.Y(n_1257)
);

AOI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1189),
.A2(n_1045),
.B(n_1040),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1189),
.A2(n_1028),
.B(n_1021),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1082),
.B(n_1019),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1109),
.A2(n_980),
.B(n_1003),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1083),
.B(n_980),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1200),
.A2(n_990),
.B(n_119),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1135),
.A2(n_110),
.B(n_196),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1089),
.A2(n_93),
.B(n_195),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1135),
.A2(n_1131),
.B(n_1164),
.Y(n_1266)
);

O2A1O1Ixp5_ASAP7_75t_L g1267 ( 
.A1(n_1086),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_SL g1268 ( 
.A(n_1085),
.B(n_33),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1141),
.A2(n_36),
.B(n_38),
.C(n_42),
.Y(n_1269)
);

AOI221x1_ASAP7_75t_L g1270 ( 
.A1(n_1218),
.A2(n_42),
.B1(n_46),
.B2(n_56),
.C(n_58),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1114),
.B(n_56),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1091),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1151),
.B(n_60),
.Y(n_1273)
);

AO32x2_ASAP7_75t_L g1274 ( 
.A1(n_1190),
.A2(n_60),
.A3(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1131),
.A2(n_140),
.B(n_192),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1077),
.A2(n_134),
.B(n_191),
.Y(n_1276)
);

NAND3xp33_ASAP7_75t_L g1277 ( 
.A(n_1090),
.B(n_66),
.C(n_67),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1094),
.B(n_66),
.Y(n_1278)
);

AOI221xp5_ASAP7_75t_L g1279 ( 
.A1(n_1179),
.A2(n_70),
.B1(n_77),
.B2(n_78),
.C(n_86),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1148),
.A2(n_88),
.B1(n_122),
.B2(n_125),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1084),
.B(n_129),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1204),
.A2(n_130),
.B(n_141),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1184),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1202),
.A2(n_152),
.B1(n_153),
.B2(n_160),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1137),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1216),
.B(n_163),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1105),
.A2(n_164),
.B(n_177),
.C(n_184),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1085),
.A2(n_187),
.B(n_201),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1144),
.A2(n_1194),
.B1(n_1166),
.B2(n_1120),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1190),
.A2(n_1200),
.A3(n_1130),
.B(n_1196),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1139),
.B(n_1123),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1204),
.A2(n_1165),
.B(n_1173),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1097),
.A2(n_1099),
.B(n_1136),
.Y(n_1293)
);

BUFx12f_ASAP7_75t_L g1294 ( 
.A(n_1149),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1153),
.Y(n_1295)
);

AO32x2_ASAP7_75t_L g1296 ( 
.A1(n_1101),
.A2(n_1179),
.A3(n_1205),
.B1(n_1147),
.B2(n_1108),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1220),
.B(n_1203),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1127),
.A2(n_1169),
.B(n_1207),
.Y(n_1298)
);

OAI22x1_ASAP7_75t_L g1299 ( 
.A1(n_1162),
.A2(n_1143),
.B1(n_1095),
.B2(n_1214),
.Y(n_1299)
);

INVx5_ASAP7_75t_L g1300 ( 
.A(n_1188),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1156),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1197),
.Y(n_1302)
);

AO21x1_ASAP7_75t_L g1303 ( 
.A1(n_1223),
.A2(n_1215),
.B(n_1104),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1193),
.A2(n_1209),
.B(n_1163),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1096),
.A2(n_1110),
.B(n_1115),
.Y(n_1305)
);

INVx5_ASAP7_75t_L g1306 ( 
.A(n_1188),
.Y(n_1306)
);

INVx5_ASAP7_75t_L g1307 ( 
.A(n_1188),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1208),
.Y(n_1308)
);

AOI221x1_ASAP7_75t_L g1309 ( 
.A1(n_1171),
.A2(n_1177),
.B1(n_1183),
.B2(n_1205),
.C(n_1213),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1157),
.A2(n_1129),
.B(n_1125),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1170),
.A2(n_1193),
.B(n_1168),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1101),
.A2(n_1180),
.A3(n_1201),
.B(n_1161),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1147),
.A2(n_1138),
.B1(n_1217),
.B2(n_1124),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1093),
.A2(n_1167),
.B(n_1206),
.Y(n_1314)
);

AND2x2_ASAP7_75t_SL g1315 ( 
.A(n_1113),
.B(n_1174),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1106),
.A2(n_1155),
.B(n_1122),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1160),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1192),
.A2(n_1198),
.B(n_1195),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1211),
.A2(n_1145),
.B1(n_1221),
.B2(n_1187),
.C(n_1186),
.Y(n_1319)
);

NOR2xp67_ASAP7_75t_SL g1320 ( 
.A(n_1212),
.B(n_1081),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1159),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1119),
.A2(n_1199),
.B(n_1159),
.Y(n_1322)
);

AOI221xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1081),
.A2(n_1187),
.B1(n_1146),
.B2(n_1186),
.C(n_1158),
.Y(n_1323)
);

OR2x6_ASAP7_75t_L g1324 ( 
.A(n_1134),
.B(n_1081),
.Y(n_1324)
);

AO21x1_ASAP7_75t_L g1325 ( 
.A1(n_1108),
.A2(n_1134),
.B(n_1222),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1158),
.A2(n_1160),
.B(n_1212),
.C(n_1186),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1146),
.B(n_1187),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_SL g1328 ( 
.A(n_1212),
.B(n_1146),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1160),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1212),
.A2(n_973),
.B1(n_946),
.B2(n_940),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1117),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1088),
.A2(n_1033),
.A3(n_1107),
.B(n_1126),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1121),
.A2(n_853),
.B(n_845),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1100),
.A2(n_1051),
.B(n_1191),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_SL g1335 ( 
.A1(n_1223),
.A2(n_1148),
.B(n_1033),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1092),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1088),
.A2(n_1033),
.A3(n_1107),
.B(n_1126),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1100),
.A2(n_1051),
.B(n_1191),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1100),
.A2(n_1051),
.B(n_1191),
.Y(n_1339)
);

BUFx2_ASAP7_75t_R g1340 ( 
.A(n_1103),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1087),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1117),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_L g1343 ( 
.A(n_1181),
.B(n_992),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1140),
.B(n_653),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1113),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1088),
.A2(n_1033),
.A3(n_1107),
.B(n_1126),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1085),
.A2(n_973),
.B1(n_946),
.B2(n_940),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1141),
.A2(n_767),
.B(n_766),
.C(n_762),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1100),
.A2(n_1051),
.B(n_1191),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1114),
.B(n_1008),
.Y(n_1350)
);

AO31x2_ASAP7_75t_L g1351 ( 
.A1(n_1088),
.A2(n_1033),
.A3(n_1107),
.B(n_1126),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1134),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1114),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1100),
.A2(n_1051),
.B(n_1191),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1088),
.A2(n_1033),
.A3(n_1107),
.B(n_1126),
.Y(n_1355)
);

OR2x6_ASAP7_75t_L g1356 ( 
.A(n_1188),
.B(n_1092),
.Y(n_1356)
);

NAND2x1p5_ASAP7_75t_L g1357 ( 
.A(n_1117),
.B(n_1113),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1107),
.A2(n_1011),
.B(n_1189),
.Y(n_1358)
);

INVxp67_ASAP7_75t_SL g1359 ( 
.A(n_1084),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1121),
.A2(n_853),
.B(n_845),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1100),
.A2(n_1051),
.B(n_1191),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1175),
.A2(n_1078),
.B(n_1088),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1140),
.B(n_653),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1140),
.B(n_653),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1079),
.A2(n_767),
.B(n_762),
.C(n_903),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1121),
.A2(n_853),
.B(n_845),
.Y(n_1366)
);

AO21x1_ASAP7_75t_L g1367 ( 
.A1(n_1086),
.A2(n_903),
.B(n_1080),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1087),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1121),
.A2(n_853),
.B(n_845),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1140),
.B(n_653),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1140),
.B(n_653),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1140),
.B(n_653),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_1084),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1121),
.A2(n_853),
.B(n_845),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1079),
.A2(n_767),
.B(n_762),
.C(n_903),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1140),
.B(n_653),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1087),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1100),
.A2(n_1051),
.B(n_1191),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_SL g1379 ( 
.A(n_1118),
.B(n_766),
.C(n_762),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1379),
.A2(n_1348),
.B(n_1365),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1268),
.A2(n_1299),
.B1(n_1313),
.B2(n_1277),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1324),
.Y(n_1382)
);

CKINVDCx11_ASAP7_75t_R g1383 ( 
.A(n_1235),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1344),
.B(n_1363),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1375),
.A2(n_1289),
.B(n_1271),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1362),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1268),
.A2(n_1347),
.B1(n_1330),
.B2(n_1277),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1226),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1364),
.A2(n_1370),
.B1(n_1371),
.B2(n_1372),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1295),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1376),
.A2(n_1279),
.B1(n_1289),
.B2(n_1347),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1300),
.Y(n_1392)
);

AND2x4_ASAP7_75t_SL g1393 ( 
.A(n_1227),
.B(n_1345),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1286),
.A2(n_1350),
.B1(n_1283),
.B2(n_1273),
.Y(n_1394)
);

BUFx4_ASAP7_75t_SL g1395 ( 
.A(n_1233),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1330),
.A2(n_1301),
.B1(n_1232),
.B2(n_1315),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1280),
.A2(n_1270),
.B(n_1269),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1294),
.A2(n_1240),
.B1(n_1353),
.B2(n_1257),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1232),
.A2(n_1225),
.B1(n_1263),
.B2(n_1280),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1331),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1272),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1227),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1237),
.B(n_1247),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1341),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1297),
.B(n_1342),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1278),
.A2(n_1252),
.B1(n_1238),
.B2(n_1368),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1377),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1263),
.A2(n_1284),
.B1(n_1335),
.B2(n_1245),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1274),
.A2(n_1328),
.B1(n_1298),
.B2(n_1316),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1245),
.A2(n_1281),
.B1(n_1303),
.B2(n_1251),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1300),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1251),
.A2(n_1297),
.B1(n_1316),
.B2(n_1305),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1321),
.A2(n_1231),
.B1(n_1343),
.B2(n_1322),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1322),
.A2(n_1367),
.B1(n_1308),
.B2(n_1302),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1274),
.A2(n_1328),
.B1(n_1298),
.B2(n_1362),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1274),
.A2(n_1359),
.B1(n_1373),
.B2(n_1285),
.Y(n_1416)
);

INVx4_ASAP7_75t_SL g1417 ( 
.A(n_1324),
.Y(n_1417)
);

INVxp33_ASAP7_75t_SL g1418 ( 
.A(n_1254),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1287),
.A2(n_1309),
.B(n_1264),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1357),
.A2(n_1236),
.B1(n_1304),
.B2(n_1260),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_1340),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1262),
.Y(n_1422)
);

BUFx8_ASAP7_75t_SL g1423 ( 
.A(n_1356),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1317),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1336),
.A2(n_1325),
.B1(n_1291),
.B2(n_1358),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1327),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1329),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1296),
.A2(n_1358),
.B1(n_1244),
.B2(n_1267),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1229),
.A2(n_1356),
.B1(n_1227),
.B2(n_1345),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1326),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1356),
.A2(n_1266),
.B1(n_1345),
.B2(n_1324),
.Y(n_1431)
);

NAND2x1_ASAP7_75t_L g1432 ( 
.A(n_1320),
.B(n_1352),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1282),
.A2(n_1275),
.B1(n_1311),
.B2(n_1249),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_SL g1434 ( 
.A(n_1300),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1311),
.A2(n_1249),
.B1(n_1292),
.B2(n_1244),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1258),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1296),
.A2(n_1288),
.B1(n_1319),
.B2(n_1307),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1306),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1318),
.A2(n_1306),
.B1(n_1307),
.B2(n_1374),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1312),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1296),
.A2(n_1319),
.B1(n_1306),
.B2(n_1307),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1248),
.A2(n_1333),
.B1(n_1369),
.B2(n_1366),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1323),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1360),
.A2(n_1228),
.B1(n_1259),
.B2(n_1253),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1276),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1261),
.A2(n_1241),
.B1(n_1256),
.B2(n_1253),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1265),
.Y(n_1447)
);

INVx6_ASAP7_75t_L g1448 ( 
.A(n_1323),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1332),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1314),
.A2(n_1261),
.B1(n_1255),
.B2(n_1246),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1314),
.A2(n_1242),
.B1(n_1346),
.B2(n_1332),
.Y(n_1451)
);

INVx6_ASAP7_75t_L g1452 ( 
.A(n_1250),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1293),
.A2(n_1243),
.B1(n_1310),
.B2(n_1338),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1332),
.B(n_1355),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1337),
.A2(n_1346),
.B1(n_1355),
.B2(n_1351),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1337),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1337),
.A2(n_1346),
.B1(n_1355),
.B2(n_1351),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1224),
.Y(n_1458)
);

BUFx12f_ASAP7_75t_L g1459 ( 
.A(n_1224),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1334),
.A2(n_1339),
.B1(n_1361),
.B2(n_1354),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1349),
.Y(n_1461)
);

CKINVDCx6p67_ASAP7_75t_R g1462 ( 
.A(n_1290),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1224),
.A2(n_1378),
.B1(n_1234),
.B2(n_1230),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1379),
.A2(n_767),
.B1(n_766),
.B2(n_762),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1233),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1226),
.Y(n_1466)
);

BUFx4_ASAP7_75t_R g1467 ( 
.A(n_1336),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1379),
.A2(n_767),
.B1(n_766),
.B2(n_762),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1365),
.A2(n_766),
.B1(n_1375),
.B2(n_767),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1379),
.A2(n_767),
.B1(n_766),
.B2(n_762),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1285),
.Y(n_1471)
);

OAI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1268),
.A2(n_1270),
.B1(n_1363),
.B2(n_1344),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1379),
.A2(n_767),
.B1(n_766),
.B2(n_762),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1226),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1379),
.A2(n_767),
.B1(n_766),
.B2(n_762),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1365),
.A2(n_766),
.B1(n_1375),
.B2(n_767),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1295),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1239),
.B(n_1350),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1226),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1268),
.A2(n_1270),
.B1(n_1363),
.B2(n_1344),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1268),
.A2(n_767),
.B1(n_1379),
.B2(n_766),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1233),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1379),
.A2(n_766),
.B1(n_762),
.B2(n_767),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1233),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1268),
.A2(n_767),
.B1(n_1379),
.B2(n_766),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1331),
.Y(n_1486)
);

INVx6_ASAP7_75t_L g1487 ( 
.A(n_1300),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1344),
.B(n_1363),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1233),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1233),
.Y(n_1490)
);

BUFx2_ASAP7_75t_SL g1491 ( 
.A(n_1295),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1300),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1268),
.A2(n_767),
.B1(n_1379),
.B2(n_766),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1331),
.Y(n_1494)
);

CKINVDCx11_ASAP7_75t_R g1495 ( 
.A(n_1235),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1226),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1379),
.A2(n_767),
.B1(n_766),
.B2(n_762),
.Y(n_1497)
);

INVx6_ASAP7_75t_L g1498 ( 
.A(n_1300),
.Y(n_1498)
);

BUFx10_ASAP7_75t_L g1499 ( 
.A(n_1233),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1268),
.A2(n_767),
.B1(n_766),
.B2(n_514),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1268),
.A2(n_767),
.B1(n_766),
.B2(n_514),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1268),
.A2(n_767),
.B1(n_1379),
.B2(n_766),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1300),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1331),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1362),
.Y(n_1505)
);

BUFx8_ASAP7_75t_L g1506 ( 
.A(n_1331),
.Y(n_1506)
);

OAI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1268),
.A2(n_1270),
.B1(n_1363),
.B2(n_1344),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1362),
.Y(n_1508)
);

BUFx8_ASAP7_75t_L g1509 ( 
.A(n_1331),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1233),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1226),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1365),
.A2(n_766),
.B1(n_1375),
.B2(n_767),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1226),
.Y(n_1513)
);

BUFx12f_ASAP7_75t_L g1514 ( 
.A(n_1285),
.Y(n_1514)
);

INVx6_ASAP7_75t_L g1515 ( 
.A(n_1300),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1379),
.A2(n_767),
.B1(n_766),
.B2(n_762),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1344),
.B(n_1363),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1268),
.A2(n_767),
.B1(n_1379),
.B2(n_766),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1379),
.A2(n_767),
.B1(n_766),
.B2(n_762),
.Y(n_1519)
);

BUFx10_ASAP7_75t_L g1520 ( 
.A(n_1233),
.Y(n_1520)
);

INVx6_ASAP7_75t_L g1521 ( 
.A(n_1300),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1405),
.Y(n_1522)
);

AO21x1_ASAP7_75t_L g1523 ( 
.A1(n_1469),
.A2(n_1512),
.B(n_1476),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1436),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1388),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1463),
.A2(n_1442),
.B(n_1446),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1459),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1407),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1456),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1404),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1396),
.B(n_1454),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1396),
.B(n_1449),
.Y(n_1532)
);

OAI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1483),
.A2(n_1385),
.B1(n_1397),
.B2(n_1380),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1466),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1474),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1479),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1478),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1496),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1426),
.Y(n_1539)
);

INVxp33_ASAP7_75t_L g1540 ( 
.A(n_1486),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1390),
.Y(n_1541)
);

AO32x2_ASAP7_75t_L g1542 ( 
.A1(n_1455),
.A2(n_1420),
.A3(n_1429),
.B1(n_1409),
.B2(n_1439),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1511),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1443),
.Y(n_1544)
);

BUFx10_ASAP7_75t_L g1545 ( 
.A(n_1465),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1460),
.A2(n_1453),
.B(n_1447),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1513),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1460),
.A2(n_1453),
.B(n_1447),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1462),
.B(n_1409),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1386),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1400),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1457),
.B(n_1399),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1386),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1443),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1505),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1508),
.Y(n_1556)
);

AO21x2_ASAP7_75t_L g1557 ( 
.A1(n_1463),
.A2(n_1442),
.B(n_1419),
.Y(n_1557)
);

OAI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1500),
.A2(n_1501),
.B1(n_1488),
.B2(n_1517),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1443),
.Y(n_1559)
);

AOI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1445),
.A2(n_1440),
.B(n_1458),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1448),
.Y(n_1561)
);

O2A1O1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1464),
.A2(n_1468),
.B(n_1497),
.C(n_1470),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1448),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1457),
.B(n_1399),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1448),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1452),
.B(n_1461),
.Y(n_1566)
);

CKINVDCx11_ASAP7_75t_R g1567 ( 
.A(n_1482),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1415),
.B(n_1387),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1506),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1389),
.B(n_1403),
.Y(n_1570)
);

INVx6_ASAP7_75t_L g1571 ( 
.A(n_1417),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1392),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1452),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1415),
.B(n_1387),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1494),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1384),
.B(n_1504),
.Y(n_1576)
);

AO21x1_ASAP7_75t_SL g1577 ( 
.A1(n_1408),
.A2(n_1381),
.B(n_1391),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1383),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1401),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1422),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1430),
.Y(n_1581)
);

INVx8_ASAP7_75t_L g1582 ( 
.A(n_1438),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1461),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1444),
.A2(n_1450),
.B(n_1433),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1450),
.A2(n_1444),
.B(n_1433),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1417),
.B(n_1382),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1506),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1392),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1452),
.Y(n_1589)
);

NAND2x1_ASAP7_75t_L g1590 ( 
.A(n_1413),
.B(n_1392),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1427),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1428),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1428),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1451),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1451),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1500),
.A2(n_1501),
.B1(n_1398),
.B2(n_1472),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1441),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1441),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1411),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1406),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1435),
.B(n_1414),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1411),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1432),
.Y(n_1603)
);

BUFx12f_ASAP7_75t_L g1604 ( 
.A(n_1495),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1435),
.A2(n_1391),
.B(n_1493),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1487),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1424),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1473),
.A2(n_1516),
.B(n_1475),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1431),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1416),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1434),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1477),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1481),
.B(n_1485),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1412),
.B(n_1425),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1472),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1490),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1480),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1498),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1519),
.B(n_1489),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1480),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1491),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1509),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1509),
.Y(n_1623)
);

AO21x1_ASAP7_75t_SL g1624 ( 
.A1(n_1410),
.A2(n_1481),
.B(n_1518),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1507),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1485),
.A2(n_1518),
.B(n_1502),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1493),
.B(n_1502),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1537),
.B(n_1394),
.Y(n_1628)
);

NAND4xp25_ASAP7_75t_L g1629 ( 
.A(n_1562),
.B(n_1437),
.C(n_1421),
.D(n_1418),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1522),
.B(n_1531),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1531),
.B(n_1437),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1591),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1607),
.Y(n_1633)
);

OAI211xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1558),
.A2(n_1608),
.B(n_1596),
.C(n_1533),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1605),
.A2(n_1492),
.B(n_1503),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1553),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1600),
.B(n_1402),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1581),
.Y(n_1638)
);

O2A1O1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1613),
.A2(n_1467),
.B(n_1510),
.C(n_1423),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1523),
.A2(n_1471),
.B1(n_1514),
.B2(n_1484),
.Y(n_1640)
);

INVx5_ASAP7_75t_L g1641 ( 
.A(n_1566),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1553),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1532),
.B(n_1499),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1530),
.Y(n_1644)
);

NAND2x1p5_ASAP7_75t_L g1645 ( 
.A(n_1581),
.B(n_1395),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1627),
.A2(n_1515),
.B1(n_1521),
.B2(n_1393),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1532),
.B(n_1499),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1527),
.B(n_1520),
.Y(n_1648)
);

AO21x2_ASAP7_75t_L g1649 ( 
.A1(n_1523),
.A2(n_1515),
.B(n_1395),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1570),
.A2(n_1515),
.B1(n_1520),
.B2(n_1619),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1527),
.B(n_1549),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1565),
.A2(n_1563),
.B1(n_1554),
.B2(n_1559),
.Y(n_1652)
);

BUFx4f_ASAP7_75t_L g1653 ( 
.A(n_1604),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1555),
.Y(n_1654)
);

BUFx4f_ASAP7_75t_SL g1655 ( 
.A(n_1541),
.Y(n_1655)
);

OA21x2_ASAP7_75t_L g1656 ( 
.A1(n_1584),
.A2(n_1548),
.B(n_1546),
.Y(n_1656)
);

O2A1O1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1615),
.A2(n_1617),
.B(n_1625),
.C(n_1620),
.Y(n_1657)
);

NAND4xp25_ASAP7_75t_SL g1658 ( 
.A(n_1568),
.B(n_1574),
.C(n_1552),
.D(n_1564),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1609),
.B(n_1568),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1626),
.A2(n_1590),
.B1(n_1609),
.B2(n_1574),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1565),
.A2(n_1563),
.B1(n_1554),
.B2(n_1561),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1586),
.B(n_1534),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1544),
.A2(n_1559),
.B1(n_1554),
.B2(n_1561),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1586),
.B(n_1535),
.Y(n_1664)
);

BUFx12f_ASAP7_75t_L g1665 ( 
.A(n_1567),
.Y(n_1665)
);

AO32x2_ASAP7_75t_L g1666 ( 
.A1(n_1572),
.A2(n_1588),
.A3(n_1599),
.B1(n_1618),
.B2(n_1606),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1535),
.B(n_1536),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1540),
.B(n_1576),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1526),
.A2(n_1585),
.B(n_1557),
.Y(n_1669)
);

OA21x2_ASAP7_75t_L g1670 ( 
.A1(n_1584),
.A2(n_1546),
.B(n_1548),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_1555),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1556),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1580),
.B(n_1524),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1538),
.B(n_1543),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1621),
.B(n_1612),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1583),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1551),
.B(n_1575),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1544),
.A2(n_1561),
.B1(n_1559),
.B2(n_1554),
.Y(n_1678)
);

AO21x2_ASAP7_75t_L g1679 ( 
.A1(n_1560),
.A2(n_1526),
.B(n_1557),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1552),
.B(n_1564),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1547),
.B(n_1525),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1567),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1626),
.A2(n_1590),
.B(n_1614),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1539),
.B(n_1528),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1579),
.B(n_1610),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1577),
.A2(n_1624),
.B1(n_1614),
.B2(n_1601),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1560),
.A2(n_1592),
.B(n_1593),
.Y(n_1687)
);

OAI211xp5_ASAP7_75t_L g1688 ( 
.A1(n_1601),
.A2(n_1598),
.B(n_1597),
.C(n_1593),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1598),
.A2(n_1592),
.B1(n_1594),
.B2(n_1595),
.C(n_1577),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1636),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1636),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1666),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1687),
.B(n_1550),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1630),
.B(n_1557),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1651),
.B(n_1687),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1638),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1683),
.B(n_1556),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1676),
.B(n_1550),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1634),
.A2(n_1561),
.B1(n_1559),
.B2(n_1573),
.C(n_1589),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1642),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1642),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1654),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1640),
.B(n_1561),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1634),
.A2(n_1623),
.B(n_1611),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1654),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1686),
.A2(n_1571),
.B1(n_1541),
.B2(n_1624),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1672),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_SL g1708 ( 
.A(n_1685),
.B(n_1603),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1650),
.A2(n_1589),
.B1(n_1573),
.B2(n_1569),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1671),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1649),
.B(n_1526),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1686),
.B(n_1589),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1674),
.B(n_1681),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1656),
.Y(n_1714)
);

BUFx12f_ASAP7_75t_L g1715 ( 
.A(n_1682),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1641),
.B(n_1529),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1644),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1684),
.B(n_1542),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1662),
.B(n_1542),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1662),
.B(n_1542),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1645),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1667),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1664),
.B(n_1542),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1664),
.B(n_1542),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1643),
.B(n_1585),
.Y(n_1725)
);

NAND4xp25_ASAP7_75t_L g1726 ( 
.A(n_1689),
.B(n_1587),
.C(n_1569),
.D(n_1622),
.Y(n_1726)
);

BUFx8_ASAP7_75t_SL g1727 ( 
.A(n_1665),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1673),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1714),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1692),
.B(n_1656),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1690),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1693),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1728),
.B(n_1680),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1692),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1692),
.B(n_1670),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1692),
.B(n_1679),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1692),
.Y(n_1737)
);

INVxp67_ASAP7_75t_SL g1738 ( 
.A(n_1693),
.Y(n_1738)
);

AOI211xp5_ASAP7_75t_L g1739 ( 
.A1(n_1704),
.A2(n_1658),
.B(n_1629),
.C(n_1639),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1727),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1704),
.A2(n_1658),
.B1(n_1689),
.B2(n_1680),
.C(n_1688),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1714),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1717),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1708),
.B(n_1679),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1695),
.B(n_1669),
.Y(n_1745)
);

INVxp67_ASAP7_75t_SL g1746 ( 
.A(n_1728),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1695),
.B(n_1633),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1690),
.Y(n_1748)
);

AOI31xp33_ASAP7_75t_L g1749 ( 
.A1(n_1703),
.A2(n_1645),
.A3(n_1660),
.B(n_1647),
.Y(n_1749)
);

BUFx3_ASAP7_75t_L g1750 ( 
.A(n_1716),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1697),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1716),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1708),
.B(n_1669),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1691),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1691),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1699),
.A2(n_1631),
.B1(n_1688),
.B2(n_1659),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1699),
.A2(n_1635),
.B(n_1657),
.Y(n_1757)
);

AOI33xp33_ASAP7_75t_L g1758 ( 
.A1(n_1697),
.A2(n_1657),
.A3(n_1632),
.B1(n_1639),
.B2(n_1709),
.B3(n_1718),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1716),
.B(n_1641),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_1710),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1708),
.B(n_1673),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1700),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1719),
.B(n_1666),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_R g1765 ( 
.A(n_1715),
.B(n_1578),
.Y(n_1765)
);

OAI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1726),
.A2(n_1628),
.B1(n_1653),
.B2(n_1668),
.C(n_1675),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1698),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1711),
.B(n_1677),
.C(n_1637),
.Y(n_1768)
);

AOI211xp5_ASAP7_75t_L g1769 ( 
.A1(n_1706),
.A2(n_1678),
.B(n_1663),
.C(n_1646),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1734),
.B(n_1719),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1754),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1733),
.B(n_1696),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1754),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1733),
.B(n_1722),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1755),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1736),
.B(n_1701),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1734),
.B(n_1720),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1746),
.B(n_1722),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1736),
.B(n_1732),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1755),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1734),
.B(n_1720),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1743),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1737),
.B(n_1759),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1763),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1763),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1737),
.B(n_1723),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1736),
.B(n_1702),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1743),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1746),
.B(n_1702),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1761),
.B(n_1738),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1768),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1737),
.B(n_1723),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1759),
.B(n_1724),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1729),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1761),
.B(n_1705),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1759),
.B(n_1724),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1731),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1738),
.B(n_1705),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1743),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1745),
.B(n_1725),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1745),
.B(n_1725),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1731),
.B(n_1707),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1764),
.B(n_1730),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1748),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1729),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1766),
.B(n_1726),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1730),
.B(n_1718),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1730),
.B(n_1713),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1735),
.B(n_1713),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1770),
.B(n_1750),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1797),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1770),
.B(n_1750),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1806),
.A2(n_1741),
.B1(n_1706),
.B2(n_1756),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1791),
.B(n_1758),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1782),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1797),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1804),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1791),
.B(n_1768),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1804),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1806),
.B(n_1758),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1772),
.B(n_1751),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1772),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1770),
.B(n_1750),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1771),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1782),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1771),
.Y(n_1826)
);

INVxp67_ASAP7_75t_L g1827 ( 
.A(n_1778),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1773),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1777),
.Y(n_1829)
);

NAND2x1p5_ASAP7_75t_L g1830 ( 
.A(n_1790),
.B(n_1711),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1777),
.B(n_1750),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1782),
.Y(n_1832)
);

AND2x4_ASAP7_75t_SL g1833 ( 
.A(n_1777),
.B(n_1760),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1773),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1774),
.B(n_1751),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1775),
.Y(n_1836)
);

INVx3_ASAP7_75t_SL g1837 ( 
.A(n_1783),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1782),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1775),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1781),
.B(n_1752),
.Y(n_1840)
);

INVx2_ASAP7_75t_SL g1841 ( 
.A(n_1781),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1774),
.B(n_1747),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1800),
.B(n_1747),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1780),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1781),
.B(n_1752),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1786),
.B(n_1752),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1780),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1784),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1784),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1785),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1783),
.B(n_1752),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1778),
.B(n_1762),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1785),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1800),
.B(n_1741),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1802),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1789),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1818),
.B(n_1790),
.Y(n_1857)
);

NOR2x1_ASAP7_75t_L g1858 ( 
.A(n_1818),
.B(n_1740),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1820),
.B(n_1808),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1814),
.B(n_1808),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1854),
.B(n_1740),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1837),
.B(n_1779),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1813),
.B(n_1808),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1822),
.B(n_1740),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1811),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1837),
.B(n_1833),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1837),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1811),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1829),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1841),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1827),
.B(n_1809),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1816),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1833),
.B(n_1783),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1856),
.B(n_1809),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1841),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1810),
.B(n_1803),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1810),
.B(n_1812),
.Y(n_1877)
);

NOR2xp67_ASAP7_75t_L g1878 ( 
.A(n_1851),
.B(n_1740),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1842),
.B(n_1779),
.Y(n_1879)
);

NOR2xp67_ASAP7_75t_SL g1880 ( 
.A(n_1852),
.B(n_1604),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1816),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1812),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1821),
.B(n_1779),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1823),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1834),
.B(n_1836),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1843),
.B(n_1715),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1851),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1847),
.B(n_1809),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1852),
.B(n_1776),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1819),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1823),
.B(n_1803),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1851),
.A2(n_1756),
.B1(n_1739),
.B2(n_1757),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1831),
.B(n_1803),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1869),
.Y(n_1894)
);

AOI321xp33_ASAP7_75t_SL g1895 ( 
.A1(n_1867),
.A2(n_1767),
.A3(n_1765),
.B1(n_1830),
.B2(n_1739),
.C(n_1792),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1858),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1863),
.B(n_1848),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1892),
.A2(n_1766),
.B1(n_1749),
.B2(n_1757),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1877),
.B(n_1831),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1861),
.B(n_1715),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1865),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1878),
.A2(n_1840),
.B1(n_1845),
.B2(n_1846),
.Y(n_1902)
);

AOI222xp33_ASAP7_75t_L g1903 ( 
.A1(n_1858),
.A2(n_1712),
.B1(n_1835),
.B2(n_1850),
.C1(n_1849),
.C2(n_1826),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1864),
.B(n_1840),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1865),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1862),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1877),
.B(n_1845),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1859),
.A2(n_1653),
.B(n_1749),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1886),
.B(n_1655),
.Y(n_1909)
);

OAI32xp33_ASAP7_75t_L g1910 ( 
.A1(n_1857),
.A2(n_1830),
.A3(n_1753),
.B1(n_1744),
.B2(n_1853),
.Y(n_1910)
);

NAND3xp33_ASAP7_75t_L g1911 ( 
.A(n_1880),
.B(n_1826),
.C(n_1824),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1862),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1873),
.Y(n_1913)
);

INVx2_ASAP7_75t_SL g1914 ( 
.A(n_1866),
.Y(n_1914)
);

AOI322xp5_ASAP7_75t_L g1915 ( 
.A1(n_1860),
.A2(n_1786),
.A3(n_1792),
.B1(n_1807),
.B2(n_1793),
.C1(n_1796),
.C2(n_1846),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1868),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1868),
.Y(n_1917)
);

NAND4xp25_ASAP7_75t_SL g1918 ( 
.A(n_1866),
.B(n_1769),
.C(n_1578),
.D(n_1753),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1876),
.B(n_1793),
.Y(n_1919)
);

NAND2xp33_ASAP7_75t_SL g1920 ( 
.A(n_1880),
.B(n_1765),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1896),
.Y(n_1921)
);

INVxp67_ASAP7_75t_SL g1922 ( 
.A(n_1906),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1894),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1914),
.B(n_1882),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1899),
.B(n_1907),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1898),
.A2(n_1887),
.B1(n_1884),
.B2(n_1882),
.Y(n_1926)
);

NOR3xp33_ASAP7_75t_L g1927 ( 
.A(n_1918),
.B(n_1857),
.C(n_1885),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1912),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1912),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1901),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1920),
.A2(n_1887),
.B1(n_1884),
.B2(n_1873),
.Y(n_1931)
);

OAI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1920),
.A2(n_1871),
.B1(n_1874),
.B2(n_1883),
.C(n_1830),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1901),
.Y(n_1933)
);

OAI21xp33_ASAP7_75t_L g1934 ( 
.A1(n_1903),
.A2(n_1888),
.B(n_1876),
.Y(n_1934)
);

AOI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1910),
.A2(n_1870),
.B1(n_1875),
.B2(n_1890),
.C(n_1872),
.Y(n_1935)
);

OAI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1902),
.A2(n_1753),
.B1(n_1875),
.B2(n_1870),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1900),
.B(n_1655),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1894),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1897),
.B(n_1883),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1908),
.A2(n_1893),
.B1(n_1891),
.B2(n_1879),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1922),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1927),
.A2(n_1911),
.B(n_1914),
.Y(n_1942)
);

AOI221xp5_ASAP7_75t_L g1943 ( 
.A1(n_1927),
.A2(n_1910),
.B1(n_1913),
.B2(n_1904),
.C(n_1895),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1926),
.A2(n_1913),
.B1(n_1899),
.B2(n_1907),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1925),
.B(n_1919),
.Y(n_1945)
);

OAI21xp33_ASAP7_75t_L g1946 ( 
.A1(n_1934),
.A2(n_1915),
.B(n_1905),
.Y(n_1946)
);

OAI322xp33_ASAP7_75t_L g1947 ( 
.A1(n_1923),
.A2(n_1916),
.A3(n_1917),
.B1(n_1881),
.B2(n_1872),
.C1(n_1890),
.C2(n_1889),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1928),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1931),
.B(n_1909),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1937),
.B(n_1919),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1929),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1924),
.B(n_1939),
.Y(n_1952)
);

NOR2x1_ASAP7_75t_L g1953 ( 
.A(n_1941),
.B(n_1938),
.Y(n_1953)
);

AOI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1942),
.A2(n_1932),
.B(n_1923),
.Y(n_1954)
);

NAND3xp33_ASAP7_75t_L g1955 ( 
.A(n_1943),
.B(n_1921),
.C(n_1935),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1946),
.B(n_1940),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1952),
.B(n_1936),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1946),
.A2(n_1933),
.B(n_1930),
.Y(n_1958)
);

O2A1O1Ixp33_ASAP7_75t_SL g1959 ( 
.A1(n_1944),
.A2(n_1881),
.B(n_1616),
.C(n_1889),
.Y(n_1959)
);

NOR4xp25_ASAP7_75t_L g1960 ( 
.A(n_1947),
.B(n_1839),
.C(n_1844),
.D(n_1828),
.Y(n_1960)
);

NAND4xp25_ASAP7_75t_L g1961 ( 
.A(n_1949),
.B(n_1622),
.C(n_1587),
.D(n_1769),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1950),
.B(n_1616),
.Y(n_1962)
);

AOI221xp5_ASAP7_75t_L g1963 ( 
.A1(n_1947),
.A2(n_1945),
.B1(n_1948),
.B2(n_1951),
.C(n_1893),
.Y(n_1963)
);

NAND3x1_ASAP7_75t_L g1964 ( 
.A(n_1953),
.B(n_1891),
.C(n_1828),
.Y(n_1964)
);

OAI221xp5_ASAP7_75t_SL g1965 ( 
.A1(n_1955),
.A2(n_1879),
.B1(n_1850),
.B2(n_1849),
.C(n_1853),
.Y(n_1965)
);

AOI211xp5_ASAP7_75t_SL g1966 ( 
.A1(n_1954),
.A2(n_1844),
.B(n_1839),
.C(n_1824),
.Y(n_1966)
);

NAND4xp75_ASAP7_75t_L g1967 ( 
.A(n_1958),
.B(n_1956),
.C(n_1963),
.D(n_1957),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_R g1968 ( 
.A(n_1962),
.B(n_1545),
.Y(n_1968)
);

AOI321xp33_ASAP7_75t_L g1969 ( 
.A1(n_1960),
.A2(n_1648),
.A3(n_1855),
.B1(n_1661),
.B2(n_1652),
.C(n_1819),
.Y(n_1969)
);

OAI221xp5_ASAP7_75t_SL g1970 ( 
.A1(n_1969),
.A2(n_1961),
.B1(n_1959),
.B2(n_1721),
.C(n_1855),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1967),
.A2(n_1817),
.B1(n_1721),
.B2(n_1786),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1965),
.A2(n_1787),
.B1(n_1776),
.B2(n_1789),
.Y(n_1972)
);

OAI211xp5_ASAP7_75t_SL g1973 ( 
.A1(n_1966),
.A2(n_1968),
.B(n_1964),
.C(n_1815),
.Y(n_1973)
);

OAI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1967),
.A2(n_1825),
.B(n_1815),
.Y(n_1974)
);

OAI211xp5_ASAP7_75t_L g1975 ( 
.A1(n_1965),
.A2(n_1582),
.B(n_1721),
.C(n_1838),
.Y(n_1975)
);

AOI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1965),
.A2(n_1582),
.B(n_1825),
.Y(n_1976)
);

NAND4xp75_ASAP7_75t_L g1977 ( 
.A(n_1974),
.B(n_1838),
.C(n_1832),
.D(n_1792),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1973),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1971),
.B(n_1807),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1976),
.B(n_1807),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1975),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1972),
.Y(n_1982)
);

OAI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1978),
.A2(n_1970),
.B1(n_1832),
.B2(n_1798),
.C(n_1795),
.Y(n_1983)
);

NOR3xp33_ASAP7_75t_SL g1984 ( 
.A(n_1981),
.B(n_1582),
.C(n_1545),
.Y(n_1984)
);

NAND3xp33_ASAP7_75t_L g1985 ( 
.A(n_1982),
.B(n_1798),
.C(n_1787),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1985),
.Y(n_1986)
);

INVx2_ASAP7_75t_SL g1987 ( 
.A(n_1986),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1987),
.A2(n_1980),
.B(n_1979),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1987),
.A2(n_1983),
.B1(n_1984),
.B2(n_1977),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1988),
.Y(n_1990)
);

XNOR2xp5_ASAP7_75t_L g1991 ( 
.A(n_1989),
.B(n_1545),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_SL g1992 ( 
.A1(n_1990),
.A2(n_1582),
.B1(n_1571),
.B2(n_1794),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1991),
.A2(n_1794),
.B1(n_1805),
.B2(n_1795),
.Y(n_1993)
);

NAND3xp33_ASAP7_75t_L g1994 ( 
.A(n_1993),
.B(n_1776),
.C(n_1787),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1992),
.A2(n_1805),
.B1(n_1794),
.B2(n_1742),
.Y(n_1995)
);

OAI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1994),
.A2(n_1800),
.B(n_1801),
.Y(n_1996)
);

CKINVDCx20_ASAP7_75t_R g1997 ( 
.A(n_1996),
.Y(n_1997)
);

AOI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1997),
.A2(n_1995),
.B1(n_1805),
.B2(n_1799),
.C(n_1788),
.Y(n_1998)
);

AOI211xp5_ASAP7_75t_L g1999 ( 
.A1(n_1998),
.A2(n_1602),
.B(n_1606),
.C(n_1618),
.Y(n_1999)
);


endmodule