module real_jpeg_23797_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_44),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_0),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_0),
.B(n_38),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_0),
.B(n_33),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_2),
.B(n_46),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_2),
.B(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_2),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_2),
.B(n_52),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_2),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_2),
.B(n_38),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_3),
.B(n_38),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_3),
.B(n_33),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_3),
.B(n_46),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_3),
.B(n_44),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_3),
.B(n_27),
.Y(n_313)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_7),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_7),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_7),
.B(n_27),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_7),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_7),
.B(n_38),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_7),
.B(n_33),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_7),
.Y(n_259)
);

INVx8_ASAP7_75t_SL g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_10),
.B(n_38),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_10),
.B(n_17),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_10),
.B(n_33),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_10),
.B(n_46),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_10),
.B(n_44),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_10),
.B(n_27),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_10),
.B(n_52),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_10),
.B(n_98),
.Y(n_300)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_12),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_12),
.B(n_38),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_12),
.B(n_33),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_12),
.B(n_46),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_12),
.B(n_44),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_12),
.B(n_27),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_12),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_12),
.B(n_98),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_13),
.B(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_13),
.B(n_27),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_14),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_14),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_14),
.B(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_14),
.B(n_204),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_14),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_14),
.B(n_33),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_15),
.B(n_46),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_15),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_15),
.B(n_38),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_15),
.B(n_44),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_15),
.B(n_27),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_15),
.B(n_52),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_16),
.B(n_33),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_16),
.B(n_38),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_16),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_16),
.B(n_46),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_44),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_16),
.B(n_27),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_16),
.B(n_52),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_16),
.B(n_56),
.Y(n_283)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_17),
.Y(n_134)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_17),
.Y(n_165)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_17),
.Y(n_196)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_104),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.C(n_88),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_22),
.A2(n_23),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_54),
.C(n_65),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_24),
.B(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_41),
.C(n_48),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_25),
.B(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_26),
.B(n_32),
.C(n_35),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_35),
.B2(n_40),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_31),
.A2(n_32),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_32),
.B(n_80),
.C(n_83),
.Y(n_95)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_33),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_68),
.C(n_71),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_35),
.A2(n_40),
.B1(n_68),
.B2(n_69),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_37),
.B(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_41),
.B(n_48),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.C(n_45),
.Y(n_41)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_42),
.B(n_43),
.CI(n_45),
.CON(n_327),
.SN(n_327)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_44),
.Y(n_294)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_48),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.CI(n_51),
.CON(n_48),
.SN(n_48)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_50),
.C(n_51),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_54),
.A2(n_65),
.B1(n_66),
.B2(n_364),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_54),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_61),
.C(n_64),
.Y(n_93)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_59),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_74),
.C(n_76),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_67),
.B(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_68),
.A2(n_69),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_68),
.B(n_304),
.C(n_305),
.Y(n_326)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_70),
.B(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_71),
.B(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_73),
.B(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_337),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_76),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_76),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_76),
.B(n_333),
.C(n_336),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_77),
.B(n_88),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_86),
.C(n_87),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_78),
.A2(n_79),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_81),
.B(n_84),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_85),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_101),
.C(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_84),
.B(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_86),
.B(n_87),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_95),
.C(n_96),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_107),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.CI(n_93),
.CON(n_90),
.SN(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_101),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_116),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_365),
.C(n_366),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_353),
.C(n_354),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_341),
.C(n_342),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_317),
.C(n_318),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_285),
.C(n_286),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_251),
.C(n_252),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_219),
.C(n_220),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_198),
.C(n_199),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_178),
.C(n_179),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_156),
.C(n_157),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.C(n_147),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_138),
.B2(n_139),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_140),
.C(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_132),
.Y(n_137)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.C(n_152),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_150),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_162),
.C(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_166),
.B(n_168),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_177),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_176),
.C(n_177),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_182),
.C(n_187),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_185),
.C(n_186),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_190),
.C(n_191),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_197),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_197),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_213),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_214),
.C(n_218),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_209),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_208),
.C(n_209),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_203),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_207),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_209),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.CI(n_212),
.CON(n_209),
.SN(n_209)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.CI(n_217),
.CON(n_214),
.SN(n_214)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_235),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_224),
.C(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_231),
.C(n_234),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g371 ( 
.A(n_226),
.Y(n_371)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.CI(n_229),
.CON(n_226),
.SN(n_226)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_228),
.C(n_229),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_242),
.C(n_249),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_242),
.B1(n_249),
.B2(n_250),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_238),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_241),
.B(n_276),
.C(n_277),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_242),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_247),
.C(n_248),
.Y(n_271)
);

INVx11_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_272),
.B2(n_284),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_273),
.C(n_274),
.Y(n_285)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_257),
.C(n_265),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_265),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_261),
.C(n_264),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_271),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_270),
.C(n_271),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_269),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_283),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_281),
.C(n_283),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_315),
.B2(n_316),
.Y(n_286)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_288),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_306),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_306),
.C(n_315),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_297),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_298),
.C(n_299),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_293),
.C(n_295),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_305),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_309),
.C(n_310),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_313),
.C(n_314),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_321),
.C(n_340),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_340),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_326),
.C(n_327),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g370 ( 
.A(n_327),
.Y(n_370)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_328),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_331),
.C(n_332),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_339),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_336),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_352),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_346),
.C(n_352),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_349),
.C(n_350),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_357),
.C(n_362),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_361),
.B2(n_362),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_367),
.Y(n_368)
);


endmodule