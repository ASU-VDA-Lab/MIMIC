module fake_jpeg_19320_n_155 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_76),
.Y(n_83)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_58),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_56),
.Y(n_79)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_69),
.B1(n_59),
.B2(n_50),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_88),
.B1(n_45),
.B2(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_90),
.Y(n_99)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_69),
.B1(n_44),
.B2(n_47),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_71),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_89),
.Y(n_91)
);

BUFx2_ASAP7_75t_SL g104 ( 
.A(n_91),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_90),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_101),
.Y(n_107)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_87),
.B1(n_80),
.B2(n_84),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_100),
.B1(n_0),
.B2(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_65),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_48),
.C(n_67),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_60),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_70),
.B1(n_66),
.B2(n_46),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_52),
.B1(n_51),
.B2(n_3),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_R g106 ( 
.A(n_103),
.B(n_61),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_119),
.B1(n_104),
.B2(n_117),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_99),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_117),
.B1(n_120),
.B2(n_0),
.Y(n_125)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_98),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_23),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_57),
.B1(n_49),
.B2(n_53),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_62),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_21),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_130),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_4),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_104),
.C(n_25),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_5),
.C(n_6),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_10),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_139),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_136),
.A2(n_123),
.B1(n_124),
.B2(n_121),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_142),
.A2(n_143),
.B(n_140),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_138),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_140),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_134),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_126),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_13),
.B(n_14),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_15),
.C(n_20),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_24),
.Y(n_155)
);


endmodule