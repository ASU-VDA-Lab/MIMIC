module fake_ariane_1495_n_3779 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_363, n_720, n_354, n_41, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_733, n_500, n_665, n_59, n_336, n_731, n_754, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_738, n_758, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_753, n_566, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_721, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_711, n_453, n_734, n_74, n_491, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_744, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_712, n_353, n_22, n_736, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_3779);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_363;
input n_720;
input n_354;
input n_41;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_733;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_736;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_3779;

wire n_2752;
wire n_3527;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_3619;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_2407;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_817;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_3765;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_3719;
wire n_2731;
wire n_3703;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_2278;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_3416;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_3145;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_813;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_829;
wire n_1062;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_2370;
wire n_1944;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_795;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_770;
wire n_3252;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_3315;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_3606;
wire n_786;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_868;
wire n_3474;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_823;
wire n_1900;
wire n_1074;
wire n_3230;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2391;
wire n_2332;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_1013;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3013;
wire n_3612;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3739;
wire n_1840;
wire n_1230;
wire n_2739;
wire n_3728;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_3271;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_2956;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_3458;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3472;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_772;
wire n_1216;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_3777;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_851;
wire n_1590;
wire n_3280;
wire n_1351;
wire n_3234;
wire n_3413;
wire n_3692;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_3698;
wire n_3716;
wire n_1179;
wire n_3284;
wire n_2703;
wire n_2926;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_1884;
wire n_912;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_3678;
wire n_2791;
wire n_762;
wire n_1468;
wire n_1661;
wire n_1253;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_2970;
wire n_3159;
wire n_966;
wire n_992;
wire n_955;
wire n_3549;
wire n_3624;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_3250;
wire n_3029;
wire n_2398;
wire n_3538;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_3530;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_3604;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3666;
wire n_3629;
wire n_3372;
wire n_990;
wire n_1623;
wire n_3559;
wire n_1903;
wire n_867;
wire n_2147;
wire n_3479;
wire n_2435;
wire n_2224;
wire n_1226;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3724;
wire n_1920;
wire n_2083;
wire n_815;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_3046;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_3741;
wire n_2388;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_3496;
wire n_3493;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3700;
wire n_3727;
wire n_976;
wire n_3567;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_1914;
wire n_965;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_2924;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1234;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_836;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3179;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_3262;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3699;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_776;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3615;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_2640;
wire n_1163;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_3642;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3498;
wire n_3513;
wire n_3682;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_3508;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_1304;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3599;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_3477;
wire n_3286;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_2075;
wire n_1726;
wire n_3263;
wire n_3542;
wire n_2523;
wire n_1945;
wire n_3569;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2496;
wire n_2031;
wire n_1258;
wire n_3260;
wire n_3349;
wire n_3761;
wire n_2118;
wire n_3222;
wire n_1740;
wire n_1602;
wire n_3139;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_777;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3653;
wire n_3035;
wire n_887;
wire n_3403;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_1202;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_3602;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2774;
wire n_2754;
wire n_2707;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_3611;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3501;
wire n_3492;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_3551;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_3766;
wire n_1711;
wire n_1219;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_3417;
wire n_2449;
wire n_890;
wire n_842;
wire n_3626;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_1373;
wire n_1975;
wire n_1081;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_3671;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_2623;
wire n_3392;
wire n_1800;
wire n_982;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_3367;
wire n_3669;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_3024;
wire n_2772;
wire n_3564;
wire n_1700;
wire n_862;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1714;
wire n_1044;
wire n_2696;
wire n_3340;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_3302;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_2489;
wire n_1161;
wire n_3685;
wire n_811;
wire n_3097;
wire n_3507;
wire n_791;
wire n_876;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_2622;
wire n_3447;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_854;
wire n_1318;
wire n_3452;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3422;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1873;
wire n_1137;
wire n_1733;
wire n_1856;
wire n_1476;
wire n_1524;
wire n_2723;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_1118;
wire n_943;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_3167;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3746;
wire n_961;
wire n_1807;
wire n_1046;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_1784;
wire n_3110;
wire n_771;
wire n_1321;
wire n_3050;
wire n_3157;
wire n_3753;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_3543;
wire n_3640;
wire n_1776;
wire n_3448;
wire n_2936;
wire n_1154;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_3718;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_3381;
wire n_807;
wire n_3455;
wire n_3736;
wire n_891;
wire n_3313;
wire n_1659;
wire n_885;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_3317;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_3560;
wire n_3345;
wire n_2170;
wire n_3605;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_3573;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_3291;
wire n_3654;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_3769;
wire n_825;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_3738;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_914;
wire n_1116;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_3462;
wire n_1197;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3731;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_3444;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_2343;
wire n_1048;
wire n_775;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3322;
wire n_2666;
wire n_3289;
wire n_1370;
wire n_1603;
wire n_2401;
wire n_2935;
wire n_889;
wire n_3255;
wire n_1549;
wire n_1066;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_3587;
wire n_3509;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1534;
wire n_1065;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_810;
wire n_3376;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_3770;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_3490;
wire n_2459;
wire n_962;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_1968;
wire n_918;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_2560;
wire n_1164;
wire n_3405;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1056;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1803;
wire n_1444;
wire n_1749;
wire n_820;
wire n_872;
wire n_1653;
wire n_3409;
wire n_3522;
wire n_3583;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3540;
wire n_3241;
wire n_1584;
wire n_1157;
wire n_848;
wire n_1664;
wire n_3481;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_3442;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3553;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_1175;
wire n_2299;
wire n_3751;
wire n_3402;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_2951;
wire n_3664;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_932;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_2503;
wire n_2270;
wire n_3470;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3259;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3676;
wire n_1564;
wire n_2010;
wire n_3677;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3558;
wire n_3576;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3658;
wire n_3091;
wire n_1024;
wire n_830;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_3521;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_956;
wire n_3360;
wire n_1930;
wire n_3687;
wire n_765;
wire n_1809;
wire n_2787;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_3575;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_3633;
wire n_857;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3379;
wire n_3111;
wire n_761;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_2569;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_816;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_3316;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2580;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_1792;
wire n_3351;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_3776;
wire n_2775;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_831;
wire n_3681;
wire n_778;
wire n_1619;
wire n_2351;
wire n_3303;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_3232;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_3445;
wire n_1409;
wire n_1588;
wire n_1684;
wire n_1148;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_904;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3285;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2705;
wire n_2664;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_3371;
wire n_1781;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3194;
wire n_3143;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_881;
wire n_1477;
wire n_1777;
wire n_1019;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_910;
wire n_3094;
wire n_1410;
wire n_939;
wire n_2297;
wire n_3441;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_2957;
wire n_1199;
wire n_865;
wire n_1983;
wire n_1273;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_1923;
wire n_3655;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_3763;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_3244;
wire n_3499;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_1821;
wire n_1168;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3593;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_3293;
wire n_2995;
wire n_3361;
wire n_1683;
wire n_2582;
wire n_1229;
wire n_3228;
wire n_3327;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_3707;
wire n_2052;
wire n_1091;
wire n_2485;
wire n_3149;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_2792;
wire n_1146;
wire n_3398;
wire n_3709;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3557;
wire n_3592;
wire n_3725;
wire n_2269;
wire n_1474;
wire n_2081;
wire n_937;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1722;
wire n_1001;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_3505;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_3547;
wire n_3771;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_773;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_3697;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_3427;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_3041;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1981;
wire n_1069;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx1_ASAP7_75t_L g761 ( 
.A(n_335),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_15),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_77),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_580),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_643),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_225),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_523),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_675),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_617),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_64),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_523),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_404),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_753),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_204),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_657),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_26),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_378),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_480),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_101),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_184),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_406),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_492),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_413),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_323),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_157),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_341),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_365),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_267),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_195),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_684),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_389),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_139),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_23),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_295),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_493),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_41),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_362),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_354),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_223),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_387),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_376),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_604),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_10),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_711),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_576),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_343),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_530),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_58),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_391),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_43),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_197),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_482),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_678),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_166),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_552),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_362),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_105),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_26),
.Y(n_818)
);

CKINVDCx14_ASAP7_75t_R g819 ( 
.A(n_695),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_574),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_483),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_411),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_132),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_526),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_101),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_320),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_252),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_98),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_709),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_662),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_107),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_554),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_699),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_456),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_164),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_567),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_229),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_710),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_498),
.Y(n_839)
);

CKINVDCx14_ASAP7_75t_R g840 ( 
.A(n_693),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_286),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_17),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_90),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_200),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_406),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_457),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_127),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_422),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_528),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_413),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_210),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_83),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_347),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_169),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_164),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_655),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_732),
.Y(n_857)
);

CKINVDCx14_ASAP7_75t_R g858 ( 
.A(n_514),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_161),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_196),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_748),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_268),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_731),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_579),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_746),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_392),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_680),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_719),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_374),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_569),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_292),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_83),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_493),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_365),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_734),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_702),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_192),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_206),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_5),
.Y(n_879)
);

BUFx2_ASAP7_75t_SL g880 ( 
.A(n_735),
.Y(n_880)
);

INVxp33_ASAP7_75t_SL g881 ( 
.A(n_482),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_742),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_205),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_574),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_259),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_213),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_698),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_418),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_368),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_615),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_194),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_708),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_747),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_681),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_278),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_522),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_313),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_96),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_730),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_676),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_521),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_541),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_389),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_575),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_348),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_569),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_407),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_602),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_455),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_260),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_300),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_564),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_240),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_740),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_84),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_215),
.Y(n_916)
);

BUFx5_ASAP7_75t_L g917 ( 
.A(n_469),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_419),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_200),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_435),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_477),
.Y(n_921)
);

CKINVDCx16_ASAP7_75t_R g922 ( 
.A(n_485),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_48),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_743),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_423),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_322),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_42),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_271),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_506),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_407),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_171),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_534),
.Y(n_932)
);

BUFx10_ASAP7_75t_L g933 ( 
.A(n_689),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_741),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_699),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_702),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_724),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_548),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_76),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_736),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_504),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_526),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_62),
.Y(n_943)
);

BUFx10_ASAP7_75t_L g944 ( 
.A(n_555),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_638),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_638),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_79),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_398),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_595),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_136),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_272),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_700),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_386),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_461),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_546),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_752),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_174),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_172),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_223),
.Y(n_959)
);

BUFx10_ASAP7_75t_L g960 ( 
.A(n_161),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_299),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_648),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_692),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_613),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_8),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_409),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_554),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_685),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_723),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_682),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_456),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_196),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_231),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_760),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_626),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_440),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_510),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_269),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_294),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_750),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_669),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_103),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_199),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_679),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_92),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_420),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_353),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_683),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_426),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_589),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_701),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_642),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_706),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_620),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_396),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_254),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_283),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_627),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_141),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_387),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_64),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_587),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_24),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_610),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_506),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_213),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_205),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_636),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_241),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_99),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_622),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_586),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_140),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_647),
.Y(n_1014)
);

BUFx10_ASAP7_75t_L g1015 ( 
.A(n_265),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_757),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_502),
.Y(n_1017)
);

BUFx10_ASAP7_75t_L g1018 ( 
.A(n_81),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_718),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_400),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_76),
.Y(n_1021)
);

CKINVDCx14_ASAP7_75t_R g1022 ( 
.A(n_374),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_4),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_621),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_183),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_486),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_514),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_505),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_221),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_613),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_339),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_58),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_225),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_48),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_332),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_501),
.Y(n_1036)
);

BUFx5_ASAP7_75t_L g1037 ( 
.A(n_172),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_729),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_135),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_250),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_241),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_479),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_758),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_508),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_369),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_744),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_355),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_292),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_180),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_166),
.Y(n_1050)
);

CKINVDCx16_ASAP7_75t_R g1051 ( 
.A(n_158),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_297),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_709),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_460),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_331),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_288),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_477),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_328),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_603),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_80),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_104),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_646),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_88),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_304),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_495),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_4),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_612),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_591),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_486),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_725),
.Y(n_1070)
);

CKINVDCx14_ASAP7_75t_R g1071 ( 
.A(n_326),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_691),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_534),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_565),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_519),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_490),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_532),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_467),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_547),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_188),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_521),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_687),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_402),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_351),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_209),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_14),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_212),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_141),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_322),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_745),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_516),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_635),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_273),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_693),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_749),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_21),
.Y(n_1096)
);

CKINVDCx16_ASAP7_75t_R g1097 ( 
.A(n_113),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_649),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_707),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_277),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_145),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_150),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_706),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_291),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_300),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_53),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_307),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_254),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_489),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_452),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_359),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_698),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_32),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_381),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_717),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_688),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_17),
.Y(n_1117)
);

BUFx8_ASAP7_75t_SL g1118 ( 
.A(n_553),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_639),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_599),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_382),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_686),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_595),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_230),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_364),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_507),
.Y(n_1126)
);

BUFx10_ASAP7_75t_L g1127 ( 
.A(n_688),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_739),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_520),
.Y(n_1129)
);

BUFx10_ASAP7_75t_L g1130 ( 
.A(n_256),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_567),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_566),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_694),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_754),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_606),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_359),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_142),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_63),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_707),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_547),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_266),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_47),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_738),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_169),
.Y(n_1144)
);

BUFx10_ASAP7_75t_L g1145 ( 
.A(n_32),
.Y(n_1145)
);

BUFx10_ASAP7_75t_L g1146 ( 
.A(n_690),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_107),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_184),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_561),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_357),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_703),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_561),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_331),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_323),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_216),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_188),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_261),
.Y(n_1157)
);

CKINVDCx14_ASAP7_75t_R g1158 ( 
.A(n_186),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_650),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_272),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_678),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_755),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_684),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_71),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_637),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_483),
.Y(n_1166)
);

BUFx5_ASAP7_75t_L g1167 ( 
.A(n_537),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_185),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_104),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_495),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_540),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_216),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_55),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_209),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_201),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_435),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_34),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_27),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_551),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_464),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_668),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_155),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_696),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_733),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_720),
.Y(n_1185)
);

CKINVDCx16_ASAP7_75t_R g1186 ( 
.A(n_634),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_669),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_404),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_346),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_680),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_140),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_704),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_751),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_253),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_108),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_294),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_659),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_737),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_472),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_491),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_690),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_123),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_116),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_587),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_75),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_697),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_462),
.Y(n_1207)
);

BUFx10_ASAP7_75t_L g1208 ( 
.A(n_73),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_385),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_360),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_605),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_471),
.Y(n_1212)
);

CKINVDCx16_ASAP7_75t_R g1213 ( 
.A(n_313),
.Y(n_1213)
);

CKINVDCx16_ASAP7_75t_R g1214 ( 
.A(n_673),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_74),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_437),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_302),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_298),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_524),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_756),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_537),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_396),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_625),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_202),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_436),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_267),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_545),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_496),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_705),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_446),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_511),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_582),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_318),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_386),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_327),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_210),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_393),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_255),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_137),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_353),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_463),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_298),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_155),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_558),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_401),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_243),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_611),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_376),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_94),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_285),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_438),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_466),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_395),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_545),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_301),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_356),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_453),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_375),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_759),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_49),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_123),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_621),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_452),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_532),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_642),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_130),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_91),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_403),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_314),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_84),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_151),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_617),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_393),
.Y(n_1273)
);

INVxp67_ASAP7_75t_SL g1274 ( 
.A(n_573),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_263),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_302),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_2),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_77),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_414),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_191),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_791),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_917),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_917),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_763),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_791),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_791),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_779),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_917),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_765),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_779),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_765),
.Y(n_1291)
);

CKINVDCx14_ASAP7_75t_R g1292 ( 
.A(n_819),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_919),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_919),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_984),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_984),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1003),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_917),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1003),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1005),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1118),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1005),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_766),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_766),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1073),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1118),
.Y(n_1306)
);

CKINVDCx14_ASAP7_75t_R g1307 ( 
.A(n_840),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1073),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1266),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1266),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_772),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_917),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_917),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_917),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1037),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_922),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1037),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1037),
.Y(n_1318)
);

INVxp67_ASAP7_75t_SL g1319 ( 
.A(n_786),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1037),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1037),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1037),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_786),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1037),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1167),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1167),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_786),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_772),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1167),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1051),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_851),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1167),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1167),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1167),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1167),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_761),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_764),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_770),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_774),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_778),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1097),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_785),
.Y(n_1342)
);

CKINVDCx16_ASAP7_75t_R g1343 ( 
.A(n_858),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_787),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_788),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_786),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_789),
.Y(n_1347)
);

CKINVDCx16_ASAP7_75t_R g1348 ( 
.A(n_1022),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1186),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_924),
.B(n_0),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_773),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_790),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_792),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_773),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_794),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_797),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_799),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_837),
.Y(n_1358)
);

CKINVDCx16_ASAP7_75t_R g1359 ( 
.A(n_1071),
.Y(n_1359)
);

INVxp33_ASAP7_75t_SL g1360 ( 
.A(n_1059),
.Y(n_1360)
);

INVxp33_ASAP7_75t_L g1361 ( 
.A(n_1243),
.Y(n_1361)
);

CKINVDCx16_ASAP7_75t_R g1362 ( 
.A(n_1158),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_860),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_809),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_811),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1213),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_860),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1214),
.Y(n_1368)
);

CKINVDCx14_ASAP7_75t_R g1369 ( 
.A(n_863),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_860),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_777),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_812),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_821),
.Y(n_1373)
);

CKINVDCx16_ASAP7_75t_R g1374 ( 
.A(n_933),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_901),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_762),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_828),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_829),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_860),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_903),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_831),
.Y(n_1381)
);

INVxp33_ASAP7_75t_SL g1382 ( 
.A(n_908),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_836),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_841),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_842),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_843),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_854),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_933),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_861),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_767),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_980),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_859),
.Y(n_1392)
);

CKINVDCx16_ASAP7_75t_R g1393 ( 
.A(n_933),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_768),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_771),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_775),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1038),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_873),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_903),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_874),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_883),
.Y(n_1401)
);

XNOR2x1_ASAP7_75t_L g1402 ( 
.A(n_793),
.B(n_0),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_888),
.Y(n_1403)
);

CKINVDCx16_ASAP7_75t_R g1404 ( 
.A(n_944),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1000),
.B(n_1),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_891),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_894),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_780),
.Y(n_1408)
);

INVxp33_ASAP7_75t_L g1409 ( 
.A(n_1139),
.Y(n_1409)
);

INVxp33_ASAP7_75t_SL g1410 ( 
.A(n_793),
.Y(n_1410)
);

INVxp33_ASAP7_75t_SL g1411 ( 
.A(n_795),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_895),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_896),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_897),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_L g1415 ( 
.A(n_769),
.B(n_803),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1090),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_769),
.Y(n_1417)
);

OAI22x1_ASAP7_75t_SL g1418 ( 
.A1(n_1289),
.A2(n_777),
.B1(n_830),
.B2(n_808),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1312),
.A2(n_914),
.B(n_857),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1319),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1351),
.B(n_803),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1375),
.Y(n_1422)
);

INVx5_ASAP7_75t_L g1423 ( 
.A(n_1282),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1363),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1323),
.B(n_1095),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1363),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1327),
.B(n_1115),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1346),
.B(n_1134),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1375),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1367),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1351),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1370),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1282),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1376),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1354),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1283),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1313),
.A2(n_914),
.B(n_857),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1354),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1316),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1283),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1314),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1292),
.B(n_944),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1370),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1288),
.Y(n_1444)
);

BUFx12f_ASAP7_75t_L g1445 ( 
.A(n_1301),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1390),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1369),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1360),
.A2(n_1033),
.B1(n_1132),
.B2(n_1025),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1399),
.B(n_1162),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1288),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1299),
.B(n_814),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1379),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1281),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1285),
.Y(n_1454)
);

BUFx12f_ASAP7_75t_L g1455 ( 
.A(n_1306),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1302),
.B(n_814),
.Y(n_1456)
);

INVx5_ASAP7_75t_L g1457 ( 
.A(n_1298),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1330),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1286),
.B(n_1185),
.Y(n_1459)
);

OA21x2_ASAP7_75t_L g1460 ( 
.A1(n_1315),
.A2(n_1128),
.B(n_1193),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1379),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1380),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1382),
.A2(n_931),
.B1(n_830),
.B2(n_872),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_SL g1464 ( 
.A(n_1343),
.B(n_1348),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1380),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1317),
.A2(n_1128),
.B(n_1198),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1292),
.B(n_1307),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1298),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1369),
.B(n_1070),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1318),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1329),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1329),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1389),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1361),
.A2(n_872),
.B1(n_887),
.B2(n_808),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1320),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1321),
.A2(n_1324),
.B(n_1322),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1402),
.A2(n_1236),
.B1(n_1129),
.B2(n_887),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1325),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1307),
.B(n_944),
.Y(n_1479)
);

INVx4_ASAP7_75t_L g1480 ( 
.A(n_1394),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1326),
.A2(n_1259),
.B(n_1070),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1359),
.B(n_960),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1332),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1333),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1334),
.B(n_865),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1395),
.Y(n_1486)
);

INVxp33_ASAP7_75t_SL g1487 ( 
.A(n_1341),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1335),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1389),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1336),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1287),
.A2(n_838),
.B(n_832),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1337),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1391),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1391),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1415),
.B(n_938),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1349),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1397),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1397),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1290),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1416),
.Y(n_1501)
);

BUFx8_ASAP7_75t_L g1502 ( 
.A(n_1358),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1416),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1362),
.B(n_960),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1338),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1293),
.A2(n_838),
.B(n_832),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1339),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1409),
.B(n_960),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1294),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1284),
.A2(n_1201),
.B1(n_1227),
.B2(n_1074),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1340),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1295),
.Y(n_1512)
);

CKINVDCx16_ASAP7_75t_R g1513 ( 
.A(n_1374),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1342),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1417),
.B(n_1296),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1344),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1297),
.B(n_938),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1300),
.B(n_1305),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1308),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1309),
.A2(n_921),
.B(n_902),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1350),
.B(n_903),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1345),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1361),
.A2(n_889),
.B1(n_970),
.B2(n_931),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1310),
.A2(n_921),
.B(n_902),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1347),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1352),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1353),
.Y(n_1527)
);

BUFx8_ASAP7_75t_L g1528 ( 
.A(n_1405),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1355),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1331),
.B(n_904),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1414),
.B(n_868),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1356),
.Y(n_1532)
);

INVx6_ASAP7_75t_L g1533 ( 
.A(n_1388),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1357),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1331),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1364),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1365),
.A2(n_990),
.B(n_936),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1372),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1350),
.B(n_1015),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1373),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_SL g1541 ( 
.A1(n_1289),
.A2(n_889),
.B1(n_1025),
.B2(n_970),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1377),
.Y(n_1542)
);

NAND2xp33_ASAP7_75t_SL g1543 ( 
.A(n_1447),
.B(n_1033),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1473),
.B(n_1396),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1535),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1472),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1509),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1508),
.B(n_1393),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1494),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1522),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1494),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1522),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1535),
.B(n_1404),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1439),
.B(n_1409),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1539),
.B(n_1408),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1450),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1450),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1534),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1534),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1536),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1539),
.B(n_1366),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1473),
.B(n_1378),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1536),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1458),
.B(n_1496),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1445),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1540),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1433),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1540),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1542),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1542),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1453),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1491),
.A2(n_1383),
.B(n_1381),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1436),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1454),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1472),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1440),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1444),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1468),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1500),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1506),
.A2(n_1385),
.B(n_1384),
.Y(n_1580)
);

NAND2xp33_ASAP7_75t_L g1581 ( 
.A(n_1447),
.B(n_1434),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1471),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1476),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1500),
.Y(n_1584)
);

CKINVDCx8_ASAP7_75t_R g1585 ( 
.A(n_1513),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1512),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1497),
.A2(n_881),
.B1(n_946),
.B2(n_864),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1431),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1493),
.B(n_1386),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1484),
.B(n_1368),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1512),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1476),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1493),
.B(n_1387),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1490),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1469),
.B(n_1392),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1431),
.B(n_1398),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1455),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1494),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1492),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1422),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1472),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1435),
.B(n_1420),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1516),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1529),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1469),
.B(n_1400),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1484),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1475),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1483),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1484),
.Y(n_1609)
);

AND2x6_ASAP7_75t_L g1610 ( 
.A(n_1467),
.B(n_1442),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1435),
.B(n_1401),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1488),
.B(n_875),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1479),
.B(n_1403),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1497),
.B(n_1406),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1498),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1498),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1422),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1532),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1488),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1441),
.B(n_1407),
.Y(n_1620)
);

INVx4_ASAP7_75t_L g1621 ( 
.A(n_1498),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1429),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1451),
.A2(n_881),
.B1(n_1050),
.B2(n_1040),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1488),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1499),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1519),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1519),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1520),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1438),
.B(n_1412),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1524),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1470),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1429),
.Y(n_1632)
);

INVx5_ASAP7_75t_L g1633 ( 
.A(n_1424),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1424),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1515),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1478),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1505),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1441),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1505),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1499),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1499),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1424),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1515),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1430),
.B(n_1489),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1419),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1505),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1451),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1507),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1503),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1507),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1507),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1482),
.B(n_1413),
.Y(n_1652)
);

INVx4_ASAP7_75t_L g1653 ( 
.A(n_1503),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1511),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1533),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1533),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1419),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1511),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1426),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1437),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1533),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1504),
.B(n_1015),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1511),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1437),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1438),
.B(n_994),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1489),
.B(n_882),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1446),
.B(n_1015),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1514),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_L g1669 ( 
.A(n_1485),
.B(n_903),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1514),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1514),
.Y(n_1671)
);

INVx2_ASAP7_75t_SL g1672 ( 
.A(n_1503),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1460),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1456),
.B(n_994),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1525),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1525),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1525),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1538),
.Y(n_1678)
);

AND2x6_ASAP7_75t_L g1679 ( 
.A(n_1673),
.B(n_1456),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1555),
.B(n_1487),
.Y(n_1680)
);

BUFx10_ASAP7_75t_L g1681 ( 
.A(n_1565),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1655),
.B(n_1446),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1546),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1580),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1647),
.A2(n_1521),
.B1(n_1460),
.B2(n_1466),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1631),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1656),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_L g1688 ( 
.A(n_1595),
.B(n_1485),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1631),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1555),
.B(n_1487),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1636),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1614),
.B(n_1480),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1548),
.B(n_1480),
.Y(n_1693)
);

INVx4_ASAP7_75t_L g1694 ( 
.A(n_1588),
.Y(n_1694)
);

OR2x6_ASAP7_75t_L g1695 ( 
.A(n_1661),
.B(n_1564),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1622),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1585),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1597),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1605),
.A2(n_1486),
.B1(n_1521),
.B2(n_1531),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1546),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1556),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1602),
.B(n_1486),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1602),
.B(n_1501),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1556),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1557),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1554),
.B(n_1464),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1632),
.B(n_1464),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1596),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1636),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1647),
.A2(n_1466),
.B1(n_1528),
.B2(n_1537),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1632),
.B(n_1448),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1546),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1613),
.B(n_1652),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1545),
.B(n_1448),
.Y(n_1714)
);

BUFx10_ASAP7_75t_L g1715 ( 
.A(n_1596),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_SL g1716 ( 
.A(n_1553),
.B(n_1474),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1557),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1667),
.B(n_1531),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_1545),
.Y(n_1719)
);

NAND2x1p5_ASAP7_75t_L g1720 ( 
.A(n_1588),
.B(n_1527),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1607),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1571),
.A2(n_1528),
.B1(n_1537),
.B2(n_1474),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1620),
.B(n_1501),
.Y(n_1723)
);

AND2x2_ASAP7_75t_SL g1724 ( 
.A(n_1623),
.B(n_1477),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1544),
.B(n_1527),
.Y(n_1725)
);

BUFx10_ASAP7_75t_L g1726 ( 
.A(n_1629),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1561),
.B(n_1530),
.Y(n_1727)
);

INVx4_ASAP7_75t_L g1728 ( 
.A(n_1621),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1594),
.B(n_1526),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1607),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1608),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1608),
.Y(n_1732)
);

INVx4_ASAP7_75t_L g1733 ( 
.A(n_1621),
.Y(n_1733)
);

INVx5_ASAP7_75t_L g1734 ( 
.A(n_1610),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1599),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1567),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1574),
.A2(n_1523),
.B1(n_1517),
.B2(n_1421),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1600),
.B(n_1463),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1635),
.B(n_1526),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1603),
.Y(n_1740)
);

INVxp33_ASAP7_75t_L g1741 ( 
.A(n_1600),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1617),
.B(n_1463),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1561),
.B(n_1425),
.Y(n_1743)
);

AND2x6_ASAP7_75t_L g1744 ( 
.A(n_1673),
.B(n_1421),
.Y(n_1744)
);

BUFx3_ASAP7_75t_L g1745 ( 
.A(n_1629),
.Y(n_1745)
);

CKINVDCx20_ASAP7_75t_R g1746 ( 
.A(n_1543),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1617),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1567),
.Y(n_1748)
);

BUFx10_ASAP7_75t_L g1749 ( 
.A(n_1674),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1604),
.B(n_1425),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1662),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1618),
.B(n_1427),
.Y(n_1752)
);

INVx4_ASAP7_75t_L g1753 ( 
.A(n_1653),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1546),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1638),
.B(n_1427),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1575),
.Y(n_1756)
);

AND2x2_ASAP7_75t_SL g1757 ( 
.A(n_1581),
.B(n_1477),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1635),
.B(n_1643),
.Y(n_1758)
);

NOR2x1p5_ASAP7_75t_L g1759 ( 
.A(n_1674),
.B(n_795),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1549),
.Y(n_1760)
);

INVx6_ASAP7_75t_L g1761 ( 
.A(n_1665),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1575),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1550),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1552),
.Y(n_1764)
);

BUFx3_ASAP7_75t_L g1765 ( 
.A(n_1549),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1573),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1558),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1643),
.B(n_1538),
.Y(n_1768)
);

BUFx10_ASAP7_75t_L g1769 ( 
.A(n_1665),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1653),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1551),
.B(n_1538),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1575),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1559),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1573),
.Y(n_1774)
);

BUFx3_ASAP7_75t_L g1775 ( 
.A(n_1551),
.Y(n_1775)
);

BUFx3_ASAP7_75t_L g1776 ( 
.A(n_1598),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1560),
.A2(n_1523),
.B1(n_1517),
.B2(n_1495),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1610),
.B(n_1495),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1598),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1638),
.B(n_1563),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1615),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1566),
.Y(n_1782)
);

OR2x6_ASAP7_75t_L g1783 ( 
.A(n_1590),
.B(n_1541),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1543),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1568),
.B(n_1428),
.Y(n_1785)
);

INVx3_ASAP7_75t_L g1786 ( 
.A(n_1615),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1616),
.B(n_1428),
.Y(n_1787)
);

INVx5_ASAP7_75t_L g1788 ( 
.A(n_1610),
.Y(n_1788)
);

INVx4_ASAP7_75t_L g1789 ( 
.A(n_1610),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1587),
.B(n_1040),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1576),
.Y(n_1791)
);

INVx5_ASAP7_75t_L g1792 ( 
.A(n_1610),
.Y(n_1792)
);

AND2x6_ASAP7_75t_L g1793 ( 
.A(n_1583),
.B(n_1518),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1569),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1616),
.B(n_1449),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1576),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1577),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1577),
.Y(n_1798)
);

AND2x6_ASAP7_75t_L g1799 ( 
.A(n_1583),
.B(n_1518),
.Y(n_1799)
);

AND2x6_ASAP7_75t_L g1800 ( 
.A(n_1592),
.B(n_1645),
.Y(n_1800)
);

INVx5_ASAP7_75t_L g1801 ( 
.A(n_1606),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1570),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1562),
.B(n_1510),
.Y(n_1803)
);

AND2x2_ASAP7_75t_SL g1804 ( 
.A(n_1581),
.B(n_1510),
.Y(n_1804)
);

AND2x6_ASAP7_75t_L g1805 ( 
.A(n_1592),
.B(n_1459),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1644),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1547),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1589),
.B(n_1449),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1625),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_1672),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1625),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1593),
.B(n_1541),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1572),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1626),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1611),
.B(n_1459),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1578),
.A2(n_1481),
.B1(n_1072),
.B2(n_1074),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1627),
.B(n_1481),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1578),
.Y(n_1818)
);

INVx4_ASAP7_75t_L g1819 ( 
.A(n_1606),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1579),
.A2(n_1086),
.B1(n_1274),
.B2(n_1047),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1582),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1582),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1584),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1601),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1575),
.Y(n_1825)
);

INVxp67_ASAP7_75t_SL g1826 ( 
.A(n_1606),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1645),
.A2(n_1072),
.B1(n_1126),
.B2(n_1050),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1637),
.B(n_1461),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1586),
.Y(n_1829)
);

AND2x6_ASAP7_75t_L g1830 ( 
.A(n_1657),
.B(n_936),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1590),
.B(n_1126),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1591),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1640),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1572),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1572),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1640),
.B(n_1129),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1657),
.A2(n_1201),
.B1(n_1203),
.B2(n_1132),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1639),
.B(n_1461),
.Y(n_1838)
);

AND2x6_ASAP7_75t_L g1839 ( 
.A(n_1660),
.B(n_990),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1711),
.B(n_1291),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1704),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1688),
.A2(n_1630),
.B(n_1628),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1724),
.A2(n_1303),
.B1(n_1304),
.B2(n_1291),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1682),
.B(n_1641),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1682),
.B(n_1641),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1702),
.B(n_1649),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1683),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1741),
.B(n_1303),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1704),
.Y(n_1849)
);

AOI22x1_ASAP7_75t_L g1850 ( 
.A1(n_1814),
.A2(n_1630),
.B1(n_1628),
.B2(n_1609),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1806),
.B(n_1660),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1735),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1701),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1815),
.B(n_1743),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1696),
.B(n_1649),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1705),
.Y(n_1856)
);

NAND3xp33_ASAP7_75t_L g1857 ( 
.A(n_1693),
.B(n_1669),
.C(n_1666),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1714),
.B(n_1304),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1740),
.Y(n_1859)
);

NOR3xp33_ASAP7_75t_L g1860 ( 
.A(n_1680),
.B(n_802),
.C(n_776),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1686),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1717),
.Y(n_1862)
);

INVx4_ASAP7_75t_L g1863 ( 
.A(n_1734),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1808),
.B(n_1646),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1736),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1748),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1766),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1687),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1689),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1719),
.B(n_1606),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1747),
.B(n_1619),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1793),
.B(n_1664),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1707),
.B(n_1619),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1690),
.B(n_1619),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1757),
.A2(n_1669),
.B1(n_1227),
.B2(n_1233),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1774),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1750),
.B(n_1752),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1713),
.B(n_1648),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1696),
.B(n_1311),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1691),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1791),
.Y(n_1881)
);

NAND2x1p5_ASAP7_75t_L g1882 ( 
.A(n_1697),
.B(n_1650),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1804),
.A2(n_1233),
.B1(n_1236),
.B2(n_1203),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1796),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_SL g1885 ( 
.A(n_1698),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1797),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1709),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1798),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1738),
.B(n_1311),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1778),
.B(n_1619),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1780),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1778),
.B(n_1651),
.Y(n_1892)
);

NAND2x1p5_ASAP7_75t_L g1893 ( 
.A(n_1734),
.B(n_1654),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1721),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1818),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1684),
.A2(n_1612),
.B(n_1664),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1679),
.B(n_1658),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1679),
.B(n_1663),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1821),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1679),
.B(n_1668),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1730),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1727),
.B(n_1670),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1822),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1749),
.B(n_1624),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1749),
.B(n_1624),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1783),
.A2(n_1371),
.B1(n_1328),
.B2(n_1671),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1793),
.B(n_1609),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1731),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1716),
.B(n_1328),
.Y(n_1909)
);

AND2x6_ASAP7_75t_L g1910 ( 
.A(n_1734),
.B(n_1601),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1695),
.B(n_1371),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1755),
.B(n_1675),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1785),
.B(n_1703),
.Y(n_1913)
);

BUFx3_ASAP7_75t_L g1914 ( 
.A(n_1681),
.Y(n_1914)
);

BUFx3_ASAP7_75t_L g1915 ( 
.A(n_1681),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1699),
.B(n_1718),
.Y(n_1916)
);

OAI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1783),
.A2(n_1280),
.B1(n_1246),
.B2(n_1065),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1742),
.B(n_1246),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1732),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1763),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1807),
.Y(n_1921)
);

NAND2xp33_ASAP7_75t_L g1922 ( 
.A(n_1788),
.B(n_1624),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1706),
.B(n_1280),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1764),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1767),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1788),
.B(n_1624),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1695),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1744),
.B(n_1676),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1744),
.B(n_1677),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1773),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1744),
.B(n_1678),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1782),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1794),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1793),
.B(n_1612),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1799),
.B(n_1634),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1799),
.B(n_1816),
.Y(n_1936)
);

NAND2xp33_ASAP7_75t_L g1937 ( 
.A(n_1788),
.B(n_1659),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1799),
.B(n_1642),
.Y(n_1938)
);

INVx5_ASAP7_75t_L g1939 ( 
.A(n_1769),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1792),
.B(n_1659),
.Y(n_1940)
);

INVxp33_ASAP7_75t_L g1941 ( 
.A(n_1836),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1805),
.B(n_1659),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1802),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1823),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1751),
.B(n_1418),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1683),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1829),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1824),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1832),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1792),
.B(n_1789),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1729),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1683),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1805),
.B(n_1659),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1805),
.B(n_1633),
.Y(n_1954)
);

INVx4_ASAP7_75t_L g1955 ( 
.A(n_1792),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1828),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1838),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1784),
.B(n_1502),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1723),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1800),
.B(n_1423),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1784),
.B(n_1502),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1803),
.B(n_1737),
.Y(n_1962)
);

INVx2_ASAP7_75t_SL g1963 ( 
.A(n_1769),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1708),
.Y(n_1964)
);

NOR2x1p5_ASAP7_75t_L g1965 ( 
.A(n_1745),
.B(n_796),
.Y(n_1965)
);

NAND2xp33_ASAP7_75t_L g1966 ( 
.A(n_1700),
.B(n_1633),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1789),
.B(n_1633),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1739),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1781),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1777),
.B(n_1633),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1786),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1758),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1800),
.B(n_1685),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1694),
.B(n_905),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1694),
.B(n_796),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1809),
.Y(n_1976)
);

INVxp67_ASAP7_75t_L g1977 ( 
.A(n_1831),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1710),
.B(n_1787),
.Y(n_1978)
);

A2O1A1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1790),
.A2(n_1065),
.B(n_1228),
.C(n_1004),
.Y(n_1979)
);

INVx8_ASAP7_75t_L g1980 ( 
.A(n_1830),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1795),
.B(n_1004),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1728),
.B(n_798),
.Y(n_1982)
);

NAND3x1_ASAP7_75t_L g1983 ( 
.A(n_1827),
.B(n_909),
.C(n_907),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1812),
.B(n_1228),
.Y(n_1984)
);

NAND2xp33_ASAP7_75t_L g1985 ( 
.A(n_1700),
.B(n_798),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1837),
.A2(n_898),
.B1(n_991),
.B2(n_850),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1728),
.B(n_1251),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1733),
.B(n_1251),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1817),
.A2(n_1109),
.B(n_1148),
.C(n_1108),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1759),
.B(n_1722),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1811),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1733),
.B(n_800),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1753),
.B(n_1152),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1768),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1753),
.B(n_1178),
.Y(n_1995)
);

OAI21xp33_ASAP7_75t_L g1996 ( 
.A1(n_1692),
.A2(n_911),
.B(n_910),
.Y(n_1996)
);

AOI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1746),
.A2(n_1195),
.B1(n_1200),
.B2(n_1188),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1833),
.Y(n_1998)
);

NOR2xp67_ASAP7_75t_L g1999 ( 
.A(n_1801),
.B(n_1465),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1770),
.B(n_1231),
.Y(n_2000)
);

A2O1A1Ixp33_ASAP7_75t_L g2001 ( 
.A1(n_1813),
.A2(n_1267),
.B(n_926),
.C(n_929),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1770),
.B(n_800),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1715),
.B(n_1726),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1761),
.B(n_801),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1771),
.Y(n_2005)
);

BUFx2_ASAP7_75t_L g2006 ( 
.A(n_1761),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1725),
.B(n_1720),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1800),
.B(n_1813),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_1715),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1852),
.Y(n_2010)
);

BUFx2_ASAP7_75t_L g2011 ( 
.A(n_1911),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1879),
.B(n_1726),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1885),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1877),
.B(n_1810),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1854),
.B(n_1760),
.Y(n_2015)
);

AO22x1_ASAP7_75t_L g2016 ( 
.A1(n_1909),
.A2(n_1839),
.B1(n_1830),
.B2(n_1775),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1859),
.Y(n_2017)
);

BUFx3_ASAP7_75t_L g2018 ( 
.A(n_1868),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1962),
.B(n_1765),
.Y(n_2019)
);

NOR3xp33_ASAP7_75t_SL g2020 ( 
.A(n_1982),
.B(n_804),
.C(n_801),
.Y(n_2020)
);

BUFx12f_ASAP7_75t_SL g2021 ( 
.A(n_1974),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1917),
.A2(n_1820),
.B1(n_1839),
.B2(n_1830),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1841),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1913),
.A2(n_1819),
.B1(n_1826),
.B2(n_1779),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1921),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1849),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1933),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1943),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1917),
.A2(n_1875),
.B1(n_1883),
.B2(n_1860),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1848),
.B(n_1883),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1959),
.B(n_1776),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1944),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1885),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1939),
.B(n_1801),
.Y(n_2034)
);

AOI21xp5_ASAP7_75t_L g2035 ( 
.A1(n_1842),
.A2(n_1835),
.B(n_1834),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1891),
.B(n_1839),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1947),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_1875),
.A2(n_782),
.B1(n_783),
.B2(n_781),
.Y(n_2038)
);

AND3x2_ASAP7_75t_SL g2039 ( 
.A(n_1949),
.B(n_1021),
.C(n_997),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1920),
.Y(n_2040)
);

NOR3xp33_ASAP7_75t_SL g2041 ( 
.A(n_1992),
.B(n_805),
.C(n_804),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1939),
.B(n_1801),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1924),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1925),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1951),
.B(n_1819),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1918),
.B(n_1700),
.Y(n_2046)
);

BUFx3_ASAP7_75t_L g2047 ( 
.A(n_1914),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1984),
.B(n_1712),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1923),
.A2(n_1117),
.B1(n_1127),
.B2(n_1018),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1930),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1864),
.B(n_1712),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1878),
.B(n_1712),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1932),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1916),
.A2(n_844),
.B1(n_845),
.B2(n_784),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1941),
.B(n_1754),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1861),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1902),
.B(n_1754),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1977),
.B(n_1754),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1983),
.A2(n_847),
.B1(n_848),
.B2(n_846),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_1840),
.A2(n_1117),
.B1(n_1127),
.B2(n_1018),
.Y(n_2060)
);

A2O1A1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_1934),
.A2(n_1021),
.B(n_1030),
.C(n_997),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1895),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1939),
.B(n_1756),
.Y(n_2063)
);

BUFx2_ASAP7_75t_L g2064 ( 
.A(n_1927),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1858),
.B(n_1018),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1892),
.B(n_1756),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1869),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1958),
.B(n_1756),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1896),
.A2(n_1772),
.B(n_1762),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1906),
.A2(n_1127),
.B1(n_1130),
.B2(n_1117),
.Y(n_2070)
);

AND2x4_ASAP7_75t_L g2071 ( 
.A(n_1892),
.B(n_1762),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_1863),
.Y(n_2072)
);

INVx1_ASAP7_75t_SL g2073 ( 
.A(n_2006),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1915),
.B(n_1762),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1880),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1889),
.B(n_1130),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1887),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_1855),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1894),
.Y(n_2079)
);

NOR2x1p5_ASAP7_75t_L g2080 ( 
.A(n_1993),
.B(n_805),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1901),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_R g2082 ( 
.A(n_1963),
.B(n_2009),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1961),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1964),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1899),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1847),
.Y(n_2086)
);

OAI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_1990),
.A2(n_807),
.B1(n_810),
.B2(n_806),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_1843),
.A2(n_1145),
.B1(n_1146),
.B2(n_1130),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_1972),
.B(n_1772),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1903),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1965),
.Y(n_2091)
);

OR2x6_ASAP7_75t_L g2092 ( 
.A(n_1980),
.B(n_1772),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1995),
.B(n_1825),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1851),
.B(n_1825),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_2000),
.B(n_1825),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1986),
.A2(n_1146),
.B1(n_1208),
.B2(n_1145),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_1974),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_R g2098 ( 
.A(n_1980),
.B(n_806),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1908),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1945),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2004),
.A2(n_852),
.B1(n_853),
.B2(n_849),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1919),
.Y(n_2102)
);

INVxp67_ASAP7_75t_SL g2103 ( 
.A(n_1937),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1851),
.B(n_807),
.Y(n_2104)
);

OR2x6_ASAP7_75t_L g2105 ( 
.A(n_1980),
.B(n_880),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1956),
.B(n_810),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1847),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1865),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1957),
.B(n_813),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_1936),
.A2(n_1146),
.B1(n_1208),
.B2(n_1145),
.Y(n_2110)
);

INVx2_ASAP7_75t_SL g2111 ( 
.A(n_1882),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1853),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1968),
.B(n_813),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1863),
.B(n_815),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1866),
.Y(n_2115)
);

BUFx4f_ASAP7_75t_L g2116 ( 
.A(n_1910),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1856),
.Y(n_2117)
);

INVx5_ASAP7_75t_L g2118 ( 
.A(n_1910),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1912),
.B(n_815),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1994),
.B(n_816),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1989),
.B(n_816),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1862),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1867),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1876),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1847),
.Y(n_2125)
);

BUFx3_ASAP7_75t_L g2126 ( 
.A(n_1969),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_SL g2127 ( 
.A(n_1955),
.B(n_817),
.Y(n_2127)
);

INVx2_ASAP7_75t_SL g2128 ( 
.A(n_2003),
.Y(n_2128)
);

HB1xp67_ASAP7_75t_L g2129 ( 
.A(n_1844),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1881),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1955),
.B(n_817),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1884),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_1910),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1886),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1997),
.B(n_1208),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1971),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1888),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_1845),
.Y(n_2138)
);

BUFx3_ASAP7_75t_L g2139 ( 
.A(n_1976),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1996),
.B(n_818),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1948),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1996),
.B(n_818),
.Y(n_2142)
);

INVxp67_ASAP7_75t_L g2143 ( 
.A(n_1991),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2005),
.Y(n_2144)
);

AND2x6_ASAP7_75t_SL g2145 ( 
.A(n_1987),
.B(n_913),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_1998),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1981),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1978),
.B(n_820),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1946),
.B(n_820),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1979),
.B(n_822),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2007),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1870),
.Y(n_2152)
);

AOI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_1890),
.A2(n_856),
.B1(n_862),
.B2(n_855),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1988),
.B(n_822),
.Y(n_2154)
);

INVx3_ASAP7_75t_L g2155 ( 
.A(n_1910),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_SL g2156 ( 
.A(n_1946),
.B(n_823),
.Y(n_2156)
);

AOI22xp5_ASAP7_75t_L g2157 ( 
.A1(n_1985),
.A2(n_867),
.B1(n_869),
.B2(n_866),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_1975),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2001),
.B(n_823),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1871),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1970),
.B(n_824),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_2083),
.B(n_1946),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_2068),
.B(n_1952),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_2116),
.B(n_1952),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_2116),
.B(n_2012),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_2030),
.B(n_1952),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2029),
.B(n_2002),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_2021),
.B(n_1904),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_2118),
.B(n_1857),
.Y(n_2169)
);

NAND2xp33_ASAP7_75t_SL g2170 ( 
.A(n_2098),
.B(n_824),
.Y(n_2170)
);

NAND2xp33_ASAP7_75t_SL g2171 ( 
.A(n_2020),
.B(n_825),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_2071),
.B(n_1905),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_2118),
.B(n_1857),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2029),
.B(n_1873),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_2118),
.B(n_1942),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_2089),
.B(n_1953),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_SL g2177 ( 
.A(n_2038),
.B(n_1954),
.Y(n_2177)
);

NAND2xp33_ASAP7_75t_SL g2178 ( 
.A(n_2041),
.B(n_825),
.Y(n_2178)
);

NAND2xp33_ASAP7_75t_SL g2179 ( 
.A(n_2082),
.B(n_826),
.Y(n_2179)
);

NAND2xp33_ASAP7_75t_SL g2180 ( 
.A(n_2015),
.B(n_826),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_2038),
.B(n_2008),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_2071),
.B(n_2008),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2065),
.B(n_827),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_2074),
.B(n_1999),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_2095),
.B(n_1907),
.Y(n_2185)
);

OR2x2_ASAP7_75t_L g2186 ( 
.A(n_2011),
.B(n_1872),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_2022),
.B(n_1907),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_2022),
.B(n_2019),
.Y(n_2188)
);

NAND2xp33_ASAP7_75t_SL g2189 ( 
.A(n_2091),
.B(n_2080),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_2066),
.B(n_1874),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_2046),
.B(n_1928),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_2084),
.B(n_2086),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_2086),
.B(n_1929),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_2086),
.B(n_1931),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2076),
.B(n_1935),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_2074),
.B(n_1999),
.Y(n_2196)
);

AND2x4_ASAP7_75t_L g2197 ( 
.A(n_2092),
.B(n_1926),
.Y(n_2197)
);

NAND2xp33_ASAP7_75t_SL g2198 ( 
.A(n_2106),
.B(n_827),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2078),
.B(n_833),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2097),
.B(n_833),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_2107),
.B(n_1938),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_SL g2202 ( 
.A(n_2107),
.B(n_1872),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_2107),
.B(n_1897),
.Y(n_2203)
);

NAND2xp33_ASAP7_75t_SL g2204 ( 
.A(n_2109),
.B(n_834),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2104),
.B(n_834),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_2125),
.B(n_1898),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2151),
.B(n_2148),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_2125),
.B(n_1900),
.Y(n_2208)
);

NAND2xp33_ASAP7_75t_SL g2209 ( 
.A(n_2154),
.B(n_2013),
.Y(n_2209)
);

NAND2xp33_ASAP7_75t_SL g2210 ( 
.A(n_2033),
.B(n_835),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_2125),
.B(n_1893),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_SL g2212 ( 
.A(n_2128),
.B(n_2158),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_2072),
.B(n_2055),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2073),
.B(n_835),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_2072),
.B(n_1940),
.Y(n_2215)
);

NAND2xp33_ASAP7_75t_SL g2216 ( 
.A(n_2114),
.B(n_839),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_2031),
.B(n_1960),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_2133),
.B(n_1960),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_2133),
.B(n_1973),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_SL g2220 ( 
.A(n_2155),
.B(n_1973),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_2155),
.B(n_1950),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2064),
.B(n_839),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_2024),
.B(n_1846),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2100),
.B(n_1068),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_SL g2225 ( 
.A(n_2018),
.B(n_1967),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_2045),
.B(n_1850),
.Y(n_2226)
);

NAND2xp33_ASAP7_75t_SL g2227 ( 
.A(n_2127),
.B(n_1068),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2054),
.B(n_1235),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_2136),
.B(n_1235),
.Y(n_2229)
);

NAND2xp33_ASAP7_75t_SL g2230 ( 
.A(n_2131),
.B(n_1237),
.Y(n_2230)
);

NAND2xp33_ASAP7_75t_SL g2231 ( 
.A(n_2119),
.B(n_1237),
.Y(n_2231)
);

AND2x2_ASAP7_75t_SL g2232 ( 
.A(n_2135),
.B(n_1922),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_2103),
.B(n_1238),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_2052),
.B(n_1238),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2010),
.B(n_1240),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2017),
.B(n_1240),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2032),
.B(n_1244),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2037),
.B(n_1244),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_2057),
.B(n_1247),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_2111),
.B(n_1247),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2040),
.B(n_1249),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2054),
.B(n_1249),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_2087),
.B(n_1250),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_SL g2244 ( 
.A(n_2058),
.B(n_1250),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2048),
.B(n_1252),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_SL g2246 ( 
.A(n_2051),
.B(n_1252),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_2146),
.B(n_1253),
.Y(n_2247)
);

NAND2xp33_ASAP7_75t_SL g2248 ( 
.A(n_2113),
.B(n_2120),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_2059),
.B(n_1253),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_2059),
.B(n_1254),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_2036),
.B(n_2043),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_2044),
.B(n_1254),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2050),
.B(n_1255),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2053),
.B(n_2147),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_2056),
.B(n_1255),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_2067),
.B(n_1256),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2075),
.B(n_1256),
.Y(n_2257)
);

NAND2xp33_ASAP7_75t_SL g2258 ( 
.A(n_2014),
.B(n_870),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_2077),
.B(n_1426),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_2079),
.B(n_1426),
.Y(n_2260)
);

NAND2xp33_ASAP7_75t_SL g2261 ( 
.A(n_2149),
.B(n_1273),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2081),
.B(n_2094),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2161),
.B(n_1432),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2047),
.B(n_1432),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2144),
.B(n_1432),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2027),
.B(n_871),
.Y(n_2266)
);

NAND2xp33_ASAP7_75t_SL g2267 ( 
.A(n_2156),
.B(n_1278),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_2129),
.B(n_1443),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2138),
.B(n_1443),
.Y(n_2269)
);

NAND2xp33_ASAP7_75t_SL g2270 ( 
.A(n_2034),
.B(n_1279),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2126),
.B(n_1443),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_2139),
.B(n_1452),
.Y(n_2272)
);

NAND2xp33_ASAP7_75t_SL g2273 ( 
.A(n_2042),
.B(n_876),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2025),
.B(n_1452),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_2028),
.B(n_1452),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_2140),
.B(n_1462),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_SL g2277 ( 
.A(n_2142),
.B(n_1462),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2063),
.B(n_1462),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2092),
.B(n_1465),
.Y(n_2279)
);

NAND2xp33_ASAP7_75t_SL g2280 ( 
.A(n_2150),
.B(n_877),
.Y(n_2280)
);

NAND2xp33_ASAP7_75t_SL g2281 ( 
.A(n_2152),
.B(n_878),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2088),
.B(n_879),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2085),
.B(n_884),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2090),
.B(n_885),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_2023),
.B(n_893),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2101),
.B(n_1263),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2026),
.B(n_899),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2102),
.B(n_886),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_2160),
.B(n_934),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2062),
.B(n_2099),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_2143),
.B(n_2093),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2157),
.B(n_937),
.Y(n_2292)
);

NAND2xp33_ASAP7_75t_SL g2293 ( 
.A(n_2159),
.B(n_1270),
.Y(n_2293)
);

NAND2xp33_ASAP7_75t_SL g2294 ( 
.A(n_2121),
.B(n_1271),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_2060),
.B(n_940),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_2108),
.B(n_956),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2115),
.B(n_969),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2070),
.B(n_890),
.Y(n_2298)
);

NAND2xp33_ASAP7_75t_SL g2299 ( 
.A(n_2096),
.B(n_892),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2124),
.B(n_974),
.Y(n_2300)
);

OR2x2_ASAP7_75t_L g2301 ( 
.A(n_2112),
.B(n_930),
.Y(n_2301)
);

NAND2xp33_ASAP7_75t_SL g2302 ( 
.A(n_2110),
.B(n_900),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2130),
.B(n_1016),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2134),
.B(n_1019),
.Y(n_2304)
);

NAND2xp33_ASAP7_75t_SL g2305 ( 
.A(n_2049),
.B(n_1261),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_2141),
.B(n_1043),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_2117),
.B(n_1046),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2122),
.B(n_1143),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_2123),
.B(n_1184),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_2132),
.B(n_2137),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2153),
.B(n_1272),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2016),
.B(n_906),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2061),
.B(n_1220),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_2069),
.B(n_912),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2105),
.B(n_915),
.Y(n_2315)
);

AND2x2_ASAP7_75t_SL g2316 ( 
.A(n_2232),
.B(n_2039),
.Y(n_2316)
);

AOI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2228),
.A2(n_2105),
.B1(n_2092),
.B2(n_918),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2242),
.B(n_939),
.Y(n_2318)
);

CKINVDCx12_ASAP7_75t_R g2319 ( 
.A(n_2301),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2207),
.B(n_2145),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2290),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2195),
.B(n_2105),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2183),
.B(n_941),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2195),
.B(n_949),
.Y(n_2324)
);

OAI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2167),
.A2(n_958),
.B1(n_959),
.B2(n_957),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2254),
.B(n_961),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2200),
.B(n_1268),
.Y(n_2327)
);

HB1xp67_ASAP7_75t_L g2328 ( 
.A(n_2186),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_2232),
.B(n_2035),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2310),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2262),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_2189),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2212),
.B(n_962),
.Y(n_2333)
);

AOI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_2281),
.A2(n_920),
.B1(n_923),
.B2(n_916),
.Y(n_2334)
);

INVx3_ASAP7_75t_L g2335 ( 
.A(n_2197),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2222),
.B(n_1275),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2188),
.B(n_968),
.Y(n_2337)
);

INVx3_ASAP7_75t_SL g2338 ( 
.A(n_2192),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2291),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2165),
.B(n_973),
.Y(n_2340)
);

BUFx6f_ASAP7_75t_L g2341 ( 
.A(n_2184),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2224),
.B(n_2315),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2190),
.Y(n_2343)
);

AND3x1_ASAP7_75t_SL g2344 ( 
.A(n_2209),
.B(n_981),
.C(n_979),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2251),
.Y(n_2345)
);

CKINVDCx20_ASAP7_75t_R g2346 ( 
.A(n_2210),
.Y(n_2346)
);

OAI21xp5_ASAP7_75t_L g2347 ( 
.A1(n_2248),
.A2(n_1966),
.B(n_986),
.Y(n_2347)
);

AOI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2249),
.A2(n_927),
.B1(n_928),
.B2(n_925),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2174),
.Y(n_2349)
);

OAI22xp5_ASAP7_75t_L g2350 ( 
.A1(n_2250),
.A2(n_988),
.B1(n_998),
.B2(n_983),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2166),
.B(n_1001),
.Y(n_2351)
);

AOI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2286),
.A2(n_2170),
.B1(n_2299),
.B2(n_2179),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2191),
.Y(n_2353)
);

AOI22xp5_ASAP7_75t_SL g2354 ( 
.A1(n_2168),
.A2(n_1008),
.B1(n_1017),
.B2(n_1006),
.Y(n_2354)
);

INVx1_ASAP7_75t_SL g2355 ( 
.A(n_2162),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2172),
.Y(n_2356)
);

BUFx3_ASAP7_75t_L g2357 ( 
.A(n_2184),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2235),
.B(n_1024),
.Y(n_2358)
);

INVx3_ASAP7_75t_SL g2359 ( 
.A(n_2229),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2236),
.B(n_1028),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2182),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2237),
.B(n_1035),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2238),
.B(n_1036),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2185),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2217),
.Y(n_2365)
);

AOI22xp5_ASAP7_75t_L g2366 ( 
.A1(n_2302),
.A2(n_935),
.B1(n_942),
.B2(n_932),
.Y(n_2366)
);

NAND2xp33_ASAP7_75t_SL g2367 ( 
.A(n_2233),
.B(n_943),
.Y(n_2367)
);

BUFx4f_ASAP7_75t_L g2368 ( 
.A(n_2197),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2311),
.B(n_1245),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2241),
.B(n_1039),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2201),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2172),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2202),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2187),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2253),
.B(n_2199),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2196),
.Y(n_2376)
);

AND2x2_ASAP7_75t_SL g2377 ( 
.A(n_2196),
.B(n_1030),
.Y(n_2377)
);

OAI22xp5_ASAP7_75t_SL g2378 ( 
.A1(n_2205),
.A2(n_1057),
.B1(n_1058),
.B2(n_1052),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_L g2379 ( 
.A(n_2214),
.B(n_945),
.Y(n_2379)
);

CKINVDCx11_ASAP7_75t_R g2380 ( 
.A(n_2279),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2219),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2220),
.Y(n_2382)
);

INVxp67_ASAP7_75t_L g2383 ( 
.A(n_2247),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2213),
.B(n_1060),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2193),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2194),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2203),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2279),
.B(n_1067),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2226),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2206),
.Y(n_2390)
);

INVx4_ASAP7_75t_L g2391 ( 
.A(n_2270),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2163),
.B(n_1076),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2208),
.Y(n_2393)
);

INVx3_ASAP7_75t_L g2394 ( 
.A(n_2312),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2283),
.B(n_1277),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2176),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2181),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2268),
.Y(n_2398)
);

OAI22xp5_ASAP7_75t_L g2399 ( 
.A1(n_2243),
.A2(n_2292),
.B1(n_2255),
.B2(n_2256),
.Y(n_2399)
);

AND2x4_ASAP7_75t_L g2400 ( 
.A(n_2164),
.B(n_1083),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2269),
.Y(n_2401)
);

BUFx8_ASAP7_75t_SL g2402 ( 
.A(n_2284),
.Y(n_2402)
);

BUFx12f_ASAP7_75t_L g2403 ( 
.A(n_2240),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_2225),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2265),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2275),
.Y(n_2406)
);

INVx2_ASAP7_75t_SL g2407 ( 
.A(n_2264),
.Y(n_2407)
);

INVx4_ASAP7_75t_L g2408 ( 
.A(n_2273),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2288),
.B(n_1088),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2274),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2239),
.B(n_1091),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_2177),
.B(n_947),
.Y(n_2412)
);

INVxp67_ASAP7_75t_L g2413 ( 
.A(n_2266),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2234),
.B(n_2246),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_2258),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_2211),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_L g2417 ( 
.A(n_2171),
.B(n_948),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2259),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2169),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2260),
.Y(n_2420)
);

CKINVDCx6p67_ASAP7_75t_R g2421 ( 
.A(n_2252),
.Y(n_2421)
);

INVx3_ASAP7_75t_SL g2422 ( 
.A(n_2257),
.Y(n_2422)
);

AOI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2305),
.A2(n_951),
.B1(n_952),
.B2(n_950),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2178),
.B(n_953),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2271),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2272),
.Y(n_2426)
);

AOI22x1_ASAP7_75t_L g2427 ( 
.A1(n_2231),
.A2(n_955),
.B1(n_963),
.B2(n_954),
.Y(n_2427)
);

BUFx2_ASAP7_75t_L g2428 ( 
.A(n_2180),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2263),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2245),
.B(n_1093),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2276),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2173),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_2198),
.Y(n_2433)
);

OAI21xp5_ASAP7_75t_L g2434 ( 
.A1(n_2223),
.A2(n_1099),
.B(n_1098),
.Y(n_2434)
);

HB1xp67_ASAP7_75t_L g2435 ( 
.A(n_2218),
.Y(n_2435)
);

BUFx12f_ASAP7_75t_L g2436 ( 
.A(n_2216),
.Y(n_2436)
);

AND3x1_ASAP7_75t_SL g2437 ( 
.A(n_2204),
.B(n_1276),
.C(n_1103),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_SL g2438 ( 
.A(n_2175),
.B(n_964),
.Y(n_2438)
);

A2O1A1Ixp33_ASAP7_75t_L g2439 ( 
.A1(n_2293),
.A2(n_1082),
.B(n_1092),
.C(n_1034),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2244),
.B(n_1101),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2277),
.Y(n_2441)
);

INVx1_ASAP7_75t_SL g2442 ( 
.A(n_2227),
.Y(n_2442)
);

AND3x1_ASAP7_75t_SL g2443 ( 
.A(n_2230),
.B(n_1110),
.C(n_1107),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2314),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2215),
.B(n_1114),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2298),
.B(n_1241),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2296),
.Y(n_2447)
);

AND3x1_ASAP7_75t_SL g2448 ( 
.A(n_2261),
.B(n_1269),
.C(n_1242),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2297),
.Y(n_2449)
);

CKINVDCx16_ASAP7_75t_R g2450 ( 
.A(n_2267),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2282),
.B(n_1116),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2295),
.B(n_1123),
.Y(n_2452)
);

BUFx2_ASAP7_75t_L g2453 ( 
.A(n_2280),
.Y(n_2453)
);

BUFx8_ASAP7_75t_L g2454 ( 
.A(n_2294),
.Y(n_2454)
);

AOI22xp33_ASAP7_75t_L g2455 ( 
.A1(n_2307),
.A2(n_1034),
.B1(n_1092),
.B2(n_1082),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2221),
.B(n_965),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_2289),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2278),
.Y(n_2458)
);

BUFx2_ASAP7_75t_L g2459 ( 
.A(n_2300),
.Y(n_2459)
);

INVx3_ASAP7_75t_L g2460 ( 
.A(n_2313),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2308),
.Y(n_2461)
);

BUFx3_ASAP7_75t_L g2462 ( 
.A(n_2380),
.Y(n_2462)
);

OAI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2434),
.A2(n_2325),
.B(n_2347),
.Y(n_2463)
);

BUFx3_ASAP7_75t_L g2464 ( 
.A(n_2357),
.Y(n_2464)
);

BUFx2_ASAP7_75t_L g2465 ( 
.A(n_2338),
.Y(n_2465)
);

NAND2x1p5_ASAP7_75t_L g2466 ( 
.A(n_2368),
.B(n_2285),
.Y(n_2466)
);

INVx3_ASAP7_75t_L g2467 ( 
.A(n_2404),
.Y(n_2467)
);

OAI21x1_ASAP7_75t_L g2468 ( 
.A1(n_2389),
.A2(n_2304),
.B(n_2303),
.Y(n_2468)
);

BUFx12f_ASAP7_75t_L g2469 ( 
.A(n_2433),
.Y(n_2469)
);

BUFx2_ASAP7_75t_SL g2470 ( 
.A(n_2346),
.Y(n_2470)
);

BUFx3_ASAP7_75t_L g2471 ( 
.A(n_2341),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2328),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2331),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2349),
.B(n_1124),
.Y(n_2474)
);

OR2x2_ASAP7_75t_L g2475 ( 
.A(n_2320),
.B(n_1135),
.Y(n_2475)
);

OAI21xp5_ASAP7_75t_L g2476 ( 
.A1(n_2337),
.A2(n_2309),
.B(n_2287),
.Y(n_2476)
);

BUFx2_ASAP7_75t_SL g2477 ( 
.A(n_2391),
.Y(n_2477)
);

OA21x2_ASAP7_75t_L g2478 ( 
.A1(n_2389),
.A2(n_2306),
.B(n_1140),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2321),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2402),
.Y(n_2480)
);

BUFx3_ASAP7_75t_L g2481 ( 
.A(n_2341),
.Y(n_2481)
);

INVx2_ASAP7_75t_SL g2482 ( 
.A(n_2341),
.Y(n_2482)
);

OAI21x1_ASAP7_75t_L g2483 ( 
.A1(n_2329),
.A2(n_1149),
.B(n_1137),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2335),
.B(n_1100),
.Y(n_2484)
);

OAI21x1_ASAP7_75t_L g2485 ( 
.A1(n_2441),
.A2(n_1151),
.B(n_1150),
.Y(n_2485)
);

OAI21x1_ASAP7_75t_L g2486 ( 
.A1(n_2441),
.A2(n_1168),
.B(n_1156),
.Y(n_2486)
);

OAI21x1_ASAP7_75t_L g2487 ( 
.A1(n_2431),
.A2(n_1182),
.B(n_1181),
.Y(n_2487)
);

HB1xp67_ASAP7_75t_L g2488 ( 
.A(n_2397),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2330),
.Y(n_2489)
);

BUFx2_ASAP7_75t_R g2490 ( 
.A(n_2332),
.Y(n_2490)
);

AOI21xp5_ASAP7_75t_L g2491 ( 
.A1(n_2412),
.A2(n_1121),
.B(n_1100),
.Y(n_2491)
);

INVx3_ASAP7_75t_L g2492 ( 
.A(n_2404),
.Y(n_2492)
);

AO21x2_ASAP7_75t_L g2493 ( 
.A1(n_2444),
.A2(n_1189),
.B(n_1187),
.Y(n_2493)
);

BUFx2_ASAP7_75t_R g2494 ( 
.A(n_2359),
.Y(n_2494)
);

OA21x2_ASAP7_75t_L g2495 ( 
.A1(n_2432),
.A2(n_1194),
.B(n_1190),
.Y(n_2495)
);

INVx1_ASAP7_75t_SL g2496 ( 
.A(n_2355),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_2404),
.Y(n_2497)
);

INVx4_ASAP7_75t_L g2498 ( 
.A(n_2391),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2335),
.B(n_1121),
.Y(n_2499)
);

BUFx3_ASAP7_75t_L g2500 ( 
.A(n_2376),
.Y(n_2500)
);

INVxp33_ASAP7_75t_SL g2501 ( 
.A(n_2415),
.Y(n_2501)
);

AOI21xp5_ASAP7_75t_L g2502 ( 
.A1(n_2374),
.A2(n_1205),
.B(n_1147),
.Y(n_2502)
);

OAI21x1_ASAP7_75t_SL g2503 ( 
.A1(n_2408),
.A2(n_1205),
.B(n_1147),
.Y(n_2503)
);

AO21x2_ASAP7_75t_L g2504 ( 
.A1(n_2444),
.A2(n_1204),
.B(n_1197),
.Y(n_2504)
);

OR2x2_ASAP7_75t_L g2505 ( 
.A(n_2322),
.B(n_1206),
.Y(n_2505)
);

BUFx2_ASAP7_75t_L g2506 ( 
.A(n_2396),
.Y(n_2506)
);

NAND3xp33_ASAP7_75t_L g2507 ( 
.A(n_2439),
.B(n_1211),
.C(n_1209),
.Y(n_2507)
);

BUFx2_ASAP7_75t_L g2508 ( 
.A(n_2339),
.Y(n_2508)
);

OAI21x1_ASAP7_75t_L g2509 ( 
.A1(n_2429),
.A2(n_1223),
.B(n_1217),
.Y(n_2509)
);

OAI21x1_ASAP7_75t_L g2510 ( 
.A1(n_2458),
.A2(n_1232),
.B(n_1224),
.Y(n_2510)
);

OAI21x1_ASAP7_75t_L g2511 ( 
.A1(n_2458),
.A2(n_1239),
.B(n_1219),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2345),
.Y(n_2512)
);

AO21x2_ASAP7_75t_L g2513 ( 
.A1(n_2398),
.A2(n_1219),
.B(n_1216),
.Y(n_2513)
);

BUFx3_ASAP7_75t_L g2514 ( 
.A(n_2368),
.Y(n_2514)
);

AO21x2_ASAP7_75t_L g2515 ( 
.A1(n_2401),
.A2(n_1248),
.B(n_1216),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2316),
.A2(n_1248),
.B1(n_1055),
.B2(n_1136),
.Y(n_2516)
);

AND2x4_ASAP7_75t_L g2517 ( 
.A(n_2356),
.B(n_977),
.Y(n_2517)
);

BUFx3_ASAP7_75t_L g2518 ( 
.A(n_2416),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2432),
.Y(n_2519)
);

OA21x2_ASAP7_75t_L g2520 ( 
.A1(n_2381),
.A2(n_967),
.B(n_966),
.Y(n_2520)
);

BUFx2_ASAP7_75t_L g2521 ( 
.A(n_2364),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2353),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2361),
.Y(n_2523)
);

AO21x2_ASAP7_75t_L g2524 ( 
.A1(n_2371),
.A2(n_1457),
.B(n_1423),
.Y(n_2524)
);

OAI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2324),
.A2(n_972),
.B(n_971),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2403),
.Y(n_2526)
);

BUFx4_ASAP7_75t_SL g2527 ( 
.A(n_2457),
.Y(n_2527)
);

AO21x2_ASAP7_75t_L g2528 ( 
.A1(n_2418),
.A2(n_1457),
.B(n_1423),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2365),
.Y(n_2529)
);

INVxp67_ASAP7_75t_L g2530 ( 
.A(n_2419),
.Y(n_2530)
);

INVx2_ASAP7_75t_SL g2531 ( 
.A(n_2342),
.Y(n_2531)
);

NAND2x1p5_ASAP7_75t_L g2532 ( 
.A(n_2416),
.B(n_977),
.Y(n_2532)
);

HB1xp67_ASAP7_75t_L g2533 ( 
.A(n_2382),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2390),
.Y(n_2534)
);

OAI21x1_ASAP7_75t_L g2535 ( 
.A1(n_2410),
.A2(n_2420),
.B(n_2406),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2373),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2372),
.Y(n_2537)
);

AOI22x1_ASAP7_75t_L g2538 ( 
.A1(n_2408),
.A2(n_976),
.B1(n_978),
.B2(n_975),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2385),
.Y(n_2539)
);

AOI22x1_ASAP7_75t_L g2540 ( 
.A1(n_2453),
.A2(n_982),
.B1(n_987),
.B2(n_985),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2386),
.Y(n_2541)
);

OAI21x1_ASAP7_75t_L g2542 ( 
.A1(n_2394),
.A2(n_713),
.B(n_712),
.Y(n_2542)
);

OA21x2_ASAP7_75t_L g2543 ( 
.A1(n_2387),
.A2(n_992),
.B(n_989),
.Y(n_2543)
);

AOI22x1_ASAP7_75t_L g2544 ( 
.A1(n_2428),
.A2(n_2450),
.B1(n_2442),
.B2(n_2436),
.Y(n_2544)
);

OAI21x1_ASAP7_75t_L g2545 ( 
.A1(n_2394),
.A2(n_715),
.B(n_714),
.Y(n_2545)
);

OR2x2_ASAP7_75t_L g2546 ( 
.A(n_2318),
.B(n_977),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2421),
.Y(n_2547)
);

NAND2x1p5_ASAP7_75t_L g2548 ( 
.A(n_2416),
.B(n_977),
.Y(n_2548)
);

BUFx3_ASAP7_75t_L g2549 ( 
.A(n_2459),
.Y(n_2549)
);

AOI22xp33_ASAP7_75t_L g2550 ( 
.A1(n_2369),
.A2(n_1136),
.B1(n_1166),
.B2(n_1055),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2393),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2435),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2343),
.B(n_1055),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2392),
.Y(n_2554)
);

BUFx3_ASAP7_75t_L g2555 ( 
.A(n_2454),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_2454),
.Y(n_2556)
);

OAI21x1_ASAP7_75t_L g2557 ( 
.A1(n_2405),
.A2(n_721),
.B(n_716),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2351),
.Y(n_2558)
);

BUFx3_ASAP7_75t_L g2559 ( 
.A(n_2447),
.Y(n_2559)
);

BUFx4f_ASAP7_75t_SL g2560 ( 
.A(n_2422),
.Y(n_2560)
);

OAI21x1_ASAP7_75t_L g2561 ( 
.A1(n_2426),
.A2(n_726),
.B(n_722),
.Y(n_2561)
);

AOI21x1_ASAP7_75t_L g2562 ( 
.A1(n_2326),
.A2(n_1136),
.B(n_1055),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2449),
.Y(n_2563)
);

BUFx8_ASAP7_75t_SL g2564 ( 
.A(n_2375),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2425),
.Y(n_2565)
);

OAI21x1_ASAP7_75t_L g2566 ( 
.A1(n_2460),
.A2(n_728),
.B(n_727),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2384),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2425),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2413),
.B(n_2445),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2489),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2516),
.A2(n_2377),
.B1(n_2352),
.B2(n_2378),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2549),
.Y(n_2572)
);

INVx3_ASAP7_75t_L g2573 ( 
.A(n_2498),
.Y(n_2573)
);

OAI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2516),
.A2(n_2317),
.B1(n_2399),
.B2(n_2366),
.Y(n_2574)
);

INVx1_ASAP7_75t_SL g2575 ( 
.A(n_2494),
.Y(n_2575)
);

BUFx12f_ASAP7_75t_L g2576 ( 
.A(n_2480),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2533),
.Y(n_2577)
);

BUFx12f_ASAP7_75t_L g2578 ( 
.A(n_2547),
.Y(n_2578)
);

INVx6_ASAP7_75t_L g2579 ( 
.A(n_2469),
.Y(n_2579)
);

CKINVDCx20_ASAP7_75t_R g2580 ( 
.A(n_2564),
.Y(n_2580)
);

INVx1_ASAP7_75t_SL g2581 ( 
.A(n_2494),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2523),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2533),
.Y(n_2583)
);

OAI22xp5_ASAP7_75t_L g2584 ( 
.A1(n_2463),
.A2(n_2354),
.B1(n_2423),
.B2(n_2334),
.Y(n_2584)
);

BUFx4f_ASAP7_75t_SL g2585 ( 
.A(n_2555),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2496),
.B(n_2336),
.Y(n_2586)
);

AOI22xp33_ASAP7_75t_L g2587 ( 
.A1(n_2520),
.A2(n_2327),
.B1(n_2323),
.B2(n_2395),
.Y(n_2587)
);

CKINVDCx11_ASAP7_75t_R g2588 ( 
.A(n_2462),
.Y(n_2588)
);

BUFx8_ASAP7_75t_L g2589 ( 
.A(n_2555),
.Y(n_2589)
);

BUFx2_ASAP7_75t_SL g2590 ( 
.A(n_2556),
.Y(n_2590)
);

AOI22xp33_ASAP7_75t_SL g2591 ( 
.A1(n_2520),
.A2(n_2451),
.B1(n_2446),
.B2(n_2452),
.Y(n_2591)
);

BUFx2_ASAP7_75t_L g2592 ( 
.A(n_2549),
.Y(n_2592)
);

AOI22xp33_ASAP7_75t_SL g2593 ( 
.A1(n_2520),
.A2(n_2417),
.B1(n_2424),
.B2(n_2460),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_2498),
.Y(n_2594)
);

CKINVDCx6p67_ASAP7_75t_R g2595 ( 
.A(n_2556),
.Y(n_2595)
);

BUFx12f_ASAP7_75t_L g2596 ( 
.A(n_2526),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_SL g2597 ( 
.A1(n_2493),
.A2(n_2461),
.B1(n_2350),
.B2(n_2400),
.Y(n_2597)
);

INVx4_ASAP7_75t_L g2598 ( 
.A(n_2465),
.Y(n_2598)
);

CKINVDCx11_ASAP7_75t_R g2599 ( 
.A(n_2462),
.Y(n_2599)
);

OAI22xp5_ASAP7_75t_L g2600 ( 
.A1(n_2463),
.A2(n_2550),
.B1(n_2560),
.B2(n_2531),
.Y(n_2600)
);

AOI22xp33_ASAP7_75t_L g2601 ( 
.A1(n_2543),
.A2(n_2440),
.B1(n_2409),
.B2(n_2383),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2550),
.A2(n_2340),
.B1(n_2348),
.B2(n_2414),
.Y(n_2602)
);

INVx1_ASAP7_75t_SL g2603 ( 
.A(n_2560),
.Y(n_2603)
);

OAI21xp33_ASAP7_75t_L g2604 ( 
.A1(n_2488),
.A2(n_2379),
.B(n_2360),
.Y(n_2604)
);

INVx3_ASAP7_75t_L g2605 ( 
.A(n_2464),
.Y(n_2605)
);

BUFx8_ASAP7_75t_L g2606 ( 
.A(n_2475),
.Y(n_2606)
);

OAI21xp33_ASAP7_75t_L g2607 ( 
.A1(n_2488),
.A2(n_2362),
.B(n_2358),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2473),
.Y(n_2608)
);

AOI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2543),
.A2(n_2400),
.B1(n_2363),
.B2(n_2370),
.Y(n_2609)
);

INVx6_ASAP7_75t_L g2610 ( 
.A(n_2464),
.Y(n_2610)
);

CKINVDCx11_ASAP7_75t_R g2611 ( 
.A(n_2496),
.Y(n_2611)
);

AOI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_2569),
.A2(n_2344),
.B1(n_2448),
.B2(n_2443),
.Y(n_2612)
);

INVx1_ASAP7_75t_SL g2613 ( 
.A(n_2564),
.Y(n_2613)
);

AOI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_2559),
.A2(n_2445),
.B1(n_2411),
.B2(n_2430),
.Y(n_2614)
);

AOI22xp33_ASAP7_75t_L g2615 ( 
.A1(n_2559),
.A2(n_2388),
.B1(n_2425),
.B2(n_2455),
.Y(n_2615)
);

CKINVDCx11_ASAP7_75t_R g2616 ( 
.A(n_2497),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2512),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2522),
.Y(n_2618)
);

CKINVDCx8_ASAP7_75t_R g2619 ( 
.A(n_2470),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2529),
.Y(n_2620)
);

BUFx3_ASAP7_75t_L g2621 ( 
.A(n_2501),
.Y(n_2621)
);

INVxp67_ASAP7_75t_SL g2622 ( 
.A(n_2530),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_SL g2623 ( 
.A1(n_2493),
.A2(n_2427),
.B1(n_2407),
.B2(n_2333),
.Y(n_2623)
);

INVx1_ASAP7_75t_SL g2624 ( 
.A(n_2527),
.Y(n_2624)
);

NAND2x1p5_ASAP7_75t_L g2625 ( 
.A(n_2514),
.B(n_2438),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_2527),
.Y(n_2626)
);

INVx6_ASAP7_75t_L g2627 ( 
.A(n_2497),
.Y(n_2627)
);

INVx1_ASAP7_75t_SL g2628 ( 
.A(n_2501),
.Y(n_2628)
);

INVx8_ASAP7_75t_L g2629 ( 
.A(n_2484),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2536),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2539),
.Y(n_2631)
);

AOI22xp33_ASAP7_75t_L g2632 ( 
.A1(n_2563),
.A2(n_2456),
.B1(n_2367),
.B2(n_1166),
.Y(n_2632)
);

AOI22xp33_ASAP7_75t_L g2633 ( 
.A1(n_2504),
.A2(n_2500),
.B1(n_2567),
.B2(n_2478),
.Y(n_2633)
);

OAI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2569),
.A2(n_2437),
.B1(n_2319),
.B2(n_1210),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_SL g2635 ( 
.A1(n_2477),
.A2(n_995),
.B1(n_996),
.B2(n_993),
.Y(n_2635)
);

OAI21xp5_ASAP7_75t_SL g2636 ( 
.A1(n_2525),
.A2(n_1166),
.B(n_1136),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2541),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2551),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2519),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_2504),
.A2(n_1169),
.B1(n_1210),
.B2(n_1166),
.Y(n_2640)
);

AO22x1_ASAP7_75t_L g2641 ( 
.A1(n_2554),
.A2(n_1002),
.B1(n_1007),
.B2(n_999),
.Y(n_2641)
);

BUFx6f_ASAP7_75t_L g2642 ( 
.A(n_2514),
.Y(n_2642)
);

BUFx2_ASAP7_75t_L g2643 ( 
.A(n_2508),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2479),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2521),
.B(n_1169),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2472),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2534),
.Y(n_2647)
);

BUFx8_ASAP7_75t_SL g2648 ( 
.A(n_2506),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2544),
.A2(n_1210),
.B1(n_1230),
.B2(n_1169),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2500),
.A2(n_1210),
.B1(n_1230),
.B2(n_1169),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2537),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2608),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2622),
.B(n_2552),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2643),
.B(n_2530),
.Y(n_2654)
);

OAI21x1_ASAP7_75t_L g2655 ( 
.A1(n_2633),
.A2(n_2562),
.B(n_2535),
.Y(n_2655)
);

OA21x2_ASAP7_75t_L g2656 ( 
.A1(n_2607),
.A2(n_2553),
.B(n_2502),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2577),
.B(n_2553),
.Y(n_2657)
);

BUFx3_ASAP7_75t_L g2658 ( 
.A(n_2589),
.Y(n_2658)
);

AO31x2_ASAP7_75t_L g2659 ( 
.A1(n_2570),
.A2(n_2568),
.A3(n_2565),
.B(n_2502),
.Y(n_2659)
);

OAI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2571),
.A2(n_2525),
.B1(n_2546),
.B2(n_2507),
.Y(n_2660)
);

BUFx8_ASAP7_75t_L g2661 ( 
.A(n_2576),
.Y(n_2661)
);

OAI21x1_ASAP7_75t_L g2662 ( 
.A1(n_2645),
.A2(n_2495),
.B(n_2542),
.Y(n_2662)
);

OA21x2_ASAP7_75t_L g2663 ( 
.A1(n_2583),
.A2(n_2474),
.B(n_2558),
.Y(n_2663)
);

OAI21x1_ASAP7_75t_L g2664 ( 
.A1(n_2600),
.A2(n_2495),
.B(n_2545),
.Y(n_2664)
);

OR2x2_ASAP7_75t_L g2665 ( 
.A(n_2646),
.B(n_2505),
.Y(n_2665)
);

AOI21xp5_ASAP7_75t_L g2666 ( 
.A1(n_2636),
.A2(n_2478),
.B(n_2495),
.Y(n_2666)
);

OR2x2_ASAP7_75t_L g2667 ( 
.A(n_2617),
.B(n_2474),
.Y(n_2667)
);

OAI21x1_ASAP7_75t_L g2668 ( 
.A1(n_2573),
.A2(n_2468),
.B(n_2511),
.Y(n_2668)
);

BUFx2_ASAP7_75t_L g2669 ( 
.A(n_2648),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2582),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2618),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2620),
.B(n_2467),
.Y(n_2672)
);

BUFx3_ASAP7_75t_L g2673 ( 
.A(n_2589),
.Y(n_2673)
);

INVxp67_ASAP7_75t_L g2674 ( 
.A(n_2572),
.Y(n_2674)
);

INVx8_ASAP7_75t_L g2675 ( 
.A(n_2596),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2630),
.Y(n_2676)
);

HB1xp67_ASAP7_75t_L g2677 ( 
.A(n_2631),
.Y(n_2677)
);

AOI21xp5_ASAP7_75t_L g2678 ( 
.A1(n_2584),
.A2(n_2478),
.B(n_2476),
.Y(n_2678)
);

AOI21xp5_ASAP7_75t_L g2679 ( 
.A1(n_2574),
.A2(n_2476),
.B(n_2503),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2637),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2638),
.B(n_2467),
.Y(n_2681)
);

INVx4_ASAP7_75t_SL g2682 ( 
.A(n_2585),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2592),
.B(n_2492),
.Y(n_2683)
);

HB1xp67_ASAP7_75t_L g2684 ( 
.A(n_2639),
.Y(n_2684)
);

OAI21xp5_ASAP7_75t_L g2685 ( 
.A1(n_2604),
.A2(n_2491),
.B(n_2487),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2644),
.Y(n_2686)
);

AOI21xp5_ASAP7_75t_L g2687 ( 
.A1(n_2649),
.A2(n_2524),
.B(n_2483),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2647),
.Y(n_2688)
);

BUFx3_ASAP7_75t_L g2689 ( 
.A(n_2621),
.Y(n_2689)
);

AOI21xp5_ASAP7_75t_L g2690 ( 
.A1(n_2602),
.A2(n_2524),
.B(n_2528),
.Y(n_2690)
);

OAI22xp5_ASAP7_75t_L g2691 ( 
.A1(n_2587),
.A2(n_2591),
.B1(n_2612),
.B2(n_2593),
.Y(n_2691)
);

CKINVDCx20_ASAP7_75t_R g2692 ( 
.A(n_2580),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_2588),
.Y(n_2693)
);

HB1xp67_ASAP7_75t_L g2694 ( 
.A(n_2605),
.Y(n_2694)
);

INVx3_ASAP7_75t_L g2695 ( 
.A(n_2610),
.Y(n_2695)
);

AOI22xp33_ASAP7_75t_L g2696 ( 
.A1(n_2601),
.A2(n_2515),
.B1(n_2513),
.B2(n_2517),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2634),
.A2(n_2528),
.B(n_2566),
.Y(n_2697)
);

AO21x2_ASAP7_75t_L g2698 ( 
.A1(n_2586),
.A2(n_2515),
.B(n_2513),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2651),
.Y(n_2699)
);

OA21x2_ASAP7_75t_L g2700 ( 
.A1(n_2609),
.A2(n_2491),
.B(n_2486),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2605),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2627),
.Y(n_2702)
);

BUFx4f_ASAP7_75t_SL g2703 ( 
.A(n_2578),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2598),
.B(n_2492),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2627),
.Y(n_2705)
);

INVx3_ASAP7_75t_L g2706 ( 
.A(n_2610),
.Y(n_2706)
);

OAI21x1_ASAP7_75t_L g2707 ( 
.A1(n_2573),
.A2(n_2485),
.B(n_2510),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2598),
.Y(n_2708)
);

OAI221xp5_ASAP7_75t_L g2709 ( 
.A1(n_2623),
.A2(n_2540),
.B1(n_2538),
.B2(n_2466),
.C(n_1056),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2611),
.B(n_2594),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2594),
.B(n_2518),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2642),
.Y(n_2712)
);

OAI21xp5_ASAP7_75t_L g2713 ( 
.A1(n_2597),
.A2(n_2640),
.B(n_2650),
.Y(n_2713)
);

INVx3_ASAP7_75t_L g2714 ( 
.A(n_2642),
.Y(n_2714)
);

OA21x2_ASAP7_75t_L g2715 ( 
.A1(n_2614),
.A2(n_2561),
.B(n_2557),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2641),
.A2(n_2548),
.B(n_2532),
.Y(n_2716)
);

BUFx3_ASAP7_75t_L g2717 ( 
.A(n_2626),
.Y(n_2717)
);

HB1xp67_ASAP7_75t_L g2718 ( 
.A(n_2642),
.Y(n_2718)
);

A2O1A1Ixp33_ASAP7_75t_L g2719 ( 
.A1(n_2632),
.A2(n_2499),
.B(n_2484),
.C(n_2518),
.Y(n_2719)
);

INVxp33_ASAP7_75t_L g2720 ( 
.A(n_2599),
.Y(n_2720)
);

NOR2x1_ASAP7_75t_SL g2721 ( 
.A(n_2590),
.B(n_2471),
.Y(n_2721)
);

A2O1A1Ixp33_ASAP7_75t_L g2722 ( 
.A1(n_2575),
.A2(n_2499),
.B(n_2509),
.C(n_2481),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2616),
.B(n_2471),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2629),
.Y(n_2724)
);

AOI21xp5_ASAP7_75t_L g2725 ( 
.A1(n_2629),
.A2(n_2548),
.B(n_2532),
.Y(n_2725)
);

A2O1A1Ixp33_ASAP7_75t_L g2726 ( 
.A1(n_2581),
.A2(n_2481),
.B(n_2517),
.C(n_1041),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2606),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2628),
.B(n_2490),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2606),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2663),
.Y(n_2730)
);

OAI221xp5_ASAP7_75t_L g2731 ( 
.A1(n_2691),
.A2(n_2625),
.B1(n_2635),
.B2(n_2615),
.C(n_2466),
.Y(n_2731)
);

INVx3_ASAP7_75t_SL g2732 ( 
.A(n_2693),
.Y(n_2732)
);

OAI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2679),
.A2(n_2619),
.B1(n_2613),
.B2(n_2624),
.Y(n_2733)
);

AOI22xp33_ASAP7_75t_SL g2734 ( 
.A1(n_2691),
.A2(n_2579),
.B1(n_2482),
.B2(n_2603),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_2692),
.Y(n_2735)
);

AND2x4_ASAP7_75t_L g2736 ( 
.A(n_2721),
.B(n_2595),
.Y(n_2736)
);

AOI22xp33_ASAP7_75t_SL g2737 ( 
.A1(n_2678),
.A2(n_2579),
.B1(n_1230),
.B2(n_1042),
.Y(n_2737)
);

AOI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2660),
.A2(n_1225),
.B1(n_1226),
.B2(n_1222),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2677),
.B(n_1230),
.Y(n_2739)
);

AND2x4_ASAP7_75t_L g2740 ( 
.A(n_2702),
.B(n_1),
.Y(n_2740)
);

INVx3_ASAP7_75t_L g2741 ( 
.A(n_2695),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2694),
.B(n_2490),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2684),
.B(n_1009),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2653),
.B(n_2657),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_L g2745 ( 
.A1(n_2713),
.A2(n_1257),
.B1(n_1011),
.B2(n_1012),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2674),
.B(n_2),
.Y(n_2746)
);

OAI21x1_ASAP7_75t_L g2747 ( 
.A1(n_2655),
.A2(n_3),
.B(n_5),
.Y(n_2747)
);

AOI211xp5_ASAP7_75t_L g2748 ( 
.A1(n_2660),
.A2(n_1013),
.B(n_1014),
.C(n_1010),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2695),
.B(n_3),
.Y(n_2749)
);

OAI221xp5_ASAP7_75t_L g2750 ( 
.A1(n_2709),
.A2(n_1026),
.B1(n_1027),
.B2(n_1023),
.C(n_1020),
.Y(n_2750)
);

OR2x6_ASAP7_75t_L g2751 ( 
.A(n_2675),
.B(n_6),
.Y(n_2751)
);

AOI22xp33_ASAP7_75t_SL g2752 ( 
.A1(n_2656),
.A2(n_1031),
.B1(n_1078),
.B2(n_1061),
.Y(n_2752)
);

OAI22xp5_ASAP7_75t_L g2753 ( 
.A1(n_2706),
.A2(n_1032),
.B1(n_1044),
.B2(n_1029),
.Y(n_2753)
);

OAI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_2706),
.A2(n_1048),
.B1(n_1049),
.B2(n_1045),
.Y(n_2754)
);

OAI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2654),
.A2(n_1054),
.B1(n_1062),
.B2(n_1053),
.Y(n_2755)
);

BUFx2_ASAP7_75t_L g2756 ( 
.A(n_2718),
.Y(n_2756)
);

HB1xp67_ASAP7_75t_L g2757 ( 
.A(n_2657),
.Y(n_2757)
);

AOI21xp33_ASAP7_75t_L g2758 ( 
.A1(n_2663),
.A2(n_1064),
.B(n_1063),
.Y(n_2758)
);

INVxp67_ASAP7_75t_L g2759 ( 
.A(n_2708),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2705),
.B(n_6),
.Y(n_2760)
);

OAI22xp33_ASAP7_75t_L g2761 ( 
.A1(n_2713),
.A2(n_1069),
.B1(n_1077),
.B2(n_1066),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_SL g2762 ( 
.A(n_2689),
.B(n_1075),
.Y(n_2762)
);

AOI22xp33_ASAP7_75t_L g2763 ( 
.A1(n_2696),
.A2(n_1234),
.B1(n_1080),
.B2(n_1081),
.Y(n_2763)
);

OAI22xp33_ASAP7_75t_L g2764 ( 
.A1(n_2685),
.A2(n_1084),
.B1(n_1087),
.B2(n_1079),
.Y(n_2764)
);

OAI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2727),
.A2(n_1089),
.B1(n_1094),
.B2(n_1085),
.Y(n_2765)
);

AND2x2_ASAP7_75t_L g2766 ( 
.A(n_2701),
.B(n_7),
.Y(n_2766)
);

AND2x4_ASAP7_75t_L g2767 ( 
.A(n_2712),
.B(n_7),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2683),
.B(n_8),
.Y(n_2768)
);

AND2x2_ASAP7_75t_SL g2769 ( 
.A(n_2669),
.B(n_9),
.Y(n_2769)
);

OAI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2685),
.A2(n_1102),
.B1(n_1104),
.B2(n_1096),
.Y(n_2770)
);

INVx3_ASAP7_75t_L g2771 ( 
.A(n_2714),
.Y(n_2771)
);

AOI22xp33_ASAP7_75t_L g2772 ( 
.A1(n_2700),
.A2(n_1218),
.B1(n_1106),
.B2(n_1111),
.Y(n_2772)
);

AOI222xp33_ASAP7_75t_L g2773 ( 
.A1(n_2664),
.A2(n_1119),
.B1(n_1112),
.B2(n_1120),
.C1(n_1113),
.C2(n_1105),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2670),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2667),
.B(n_1122),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_SL g2776 ( 
.A1(n_2656),
.A2(n_1160),
.B1(n_1173),
.B2(n_1141),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2741),
.B(n_2756),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2730),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2741),
.B(n_2714),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2757),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2739),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2742),
.B(n_2728),
.Y(n_2782)
);

HB1xp67_ASAP7_75t_L g2783 ( 
.A(n_2759),
.Y(n_2783)
);

NOR2x1_ASAP7_75t_SL g2784 ( 
.A(n_2751),
.B(n_2658),
.Y(n_2784)
);

BUFx6f_ASAP7_75t_L g2785 ( 
.A(n_2747),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2771),
.B(n_2710),
.Y(n_2786)
);

HB1xp67_ASAP7_75t_L g2787 ( 
.A(n_2744),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2774),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2743),
.B(n_2652),
.Y(n_2789)
);

BUFx4f_ASAP7_75t_SL g2790 ( 
.A(n_2732),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2771),
.B(n_2704),
.Y(n_2791)
);

AND2x4_ASAP7_75t_L g2792 ( 
.A(n_2736),
.B(n_2682),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_2736),
.B(n_2720),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2768),
.B(n_2671),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2766),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2738),
.B(n_2676),
.Y(n_2796)
);

OR2x2_ASAP7_75t_L g2797 ( 
.A(n_2775),
.B(n_2665),
.Y(n_2797)
);

BUFx3_ASAP7_75t_L g2798 ( 
.A(n_2735),
.Y(n_2798)
);

OA21x2_ASAP7_75t_L g2799 ( 
.A1(n_2772),
.A2(n_2690),
.B(n_2662),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2767),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2767),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2746),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2749),
.Y(n_2803)
);

INVx2_ASAP7_75t_SL g2804 ( 
.A(n_2740),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2738),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2760),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2740),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2769),
.B(n_2680),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2734),
.B(n_2672),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2752),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2751),
.B(n_2711),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2751),
.Y(n_2812)
);

AOI22xp33_ASAP7_75t_L g2813 ( 
.A1(n_2761),
.A2(n_2698),
.B1(n_2700),
.B2(n_2666),
.Y(n_2813)
);

HB1xp67_ASAP7_75t_L g2814 ( 
.A(n_2733),
.Y(n_2814)
);

BUFx2_ASAP7_75t_L g2815 ( 
.A(n_2792),
.Y(n_2815)
);

AOI21xp33_ASAP7_75t_L g2816 ( 
.A1(n_2799),
.A2(n_2748),
.B(n_2773),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2785),
.Y(n_2817)
);

AO21x2_ASAP7_75t_L g2818 ( 
.A1(n_2778),
.A2(n_2758),
.B(n_2764),
.Y(n_2818)
);

OAI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_2814),
.A2(n_2748),
.B1(n_2737),
.B2(n_2745),
.Y(n_2819)
);

AOI22xp33_ASAP7_75t_L g2820 ( 
.A1(n_2805),
.A2(n_2731),
.B1(n_2770),
.B2(n_2776),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2785),
.Y(n_2821)
);

OAI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2809),
.A2(n_2729),
.B1(n_2723),
.B2(n_2724),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2785),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2780),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2780),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2797),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2778),
.Y(n_2827)
);

AOI21xp5_ASAP7_75t_L g2828 ( 
.A1(n_2784),
.A2(n_2793),
.B(n_2805),
.Y(n_2828)
);

OAI21xp33_ASAP7_75t_SL g2829 ( 
.A1(n_2782),
.A2(n_2681),
.B(n_2762),
.Y(n_2829)
);

OAI21xp33_ASAP7_75t_L g2830 ( 
.A1(n_2787),
.A2(n_2755),
.B(n_2765),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2785),
.Y(n_2831)
);

CKINVDCx14_ASAP7_75t_R g2832 ( 
.A(n_2792),
.Y(n_2832)
);

AND2x4_ASAP7_75t_SL g2833 ( 
.A(n_2792),
.B(n_2682),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2785),
.Y(n_2834)
);

OAI211xp5_ASAP7_75t_SL g2835 ( 
.A1(n_2796),
.A2(n_2750),
.B(n_2754),
.C(n_2753),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2797),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2786),
.B(n_2673),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2812),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2803),
.Y(n_2839)
);

INVx3_ASAP7_75t_L g2840 ( 
.A(n_2792),
.Y(n_2840)
);

AOI22xp33_ASAP7_75t_SL g2841 ( 
.A1(n_2784),
.A2(n_2715),
.B1(n_2698),
.B2(n_2697),
.Y(n_2841)
);

CKINVDCx20_ASAP7_75t_R g2842 ( 
.A(n_2790),
.Y(n_2842)
);

OAI22xp33_ASAP7_75t_L g2843 ( 
.A1(n_2812),
.A2(n_2715),
.B1(n_2703),
.B2(n_2687),
.Y(n_2843)
);

AND2x4_ASAP7_75t_L g2844 ( 
.A(n_2804),
.B(n_2717),
.Y(n_2844)
);

BUFx6f_ASAP7_75t_L g2845 ( 
.A(n_2798),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2781),
.Y(n_2846)
);

A2O1A1Ixp33_ASAP7_75t_L g2847 ( 
.A1(n_2810),
.A2(n_2726),
.B(n_2763),
.C(n_2722),
.Y(n_2847)
);

OAI21x1_ASAP7_75t_L g2848 ( 
.A1(n_2777),
.A2(n_2668),
.B(n_2686),
.Y(n_2848)
);

OAI21x1_ASAP7_75t_L g2849 ( 
.A1(n_2777),
.A2(n_2699),
.B(n_2688),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2803),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2783),
.B(n_2707),
.Y(n_2851)
);

AND2x4_ASAP7_75t_SL g2852 ( 
.A(n_2782),
.B(n_2807),
.Y(n_2852)
);

AND2x4_ASAP7_75t_L g2853 ( 
.A(n_2804),
.B(n_2659),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2803),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2826),
.B(n_2781),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2818),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2832),
.B(n_2786),
.Y(n_2857)
);

HB1xp67_ASAP7_75t_L g2858 ( 
.A(n_2824),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2832),
.B(n_2811),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2836),
.B(n_2794),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2816),
.B(n_2794),
.Y(n_2861)
);

NAND3xp33_ASAP7_75t_SL g2862 ( 
.A(n_2828),
.B(n_2813),
.C(n_2810),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2846),
.Y(n_2863)
);

AOI221xp5_ASAP7_75t_L g2864 ( 
.A1(n_2843),
.A2(n_2808),
.B1(n_2789),
.B2(n_2795),
.C(n_2802),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2852),
.B(n_2811),
.Y(n_2865)
);

BUFx3_ASAP7_75t_L g2866 ( 
.A(n_2842),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2852),
.B(n_2791),
.Y(n_2867)
);

OAI31xp33_ASAP7_75t_L g2868 ( 
.A1(n_2843),
.A2(n_2808),
.A3(n_2806),
.B(n_2795),
.Y(n_2868)
);

OR2x2_ASAP7_75t_L g2869 ( 
.A(n_2825),
.B(n_2802),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2839),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2815),
.B(n_2791),
.Y(n_2871)
);

OR2x2_ASAP7_75t_L g2872 ( 
.A(n_2854),
.B(n_2806),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2839),
.Y(n_2873)
);

OR2x2_ASAP7_75t_L g2874 ( 
.A(n_2850),
.B(n_2800),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_2842),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2850),
.Y(n_2876)
);

OR2x2_ASAP7_75t_L g2877 ( 
.A(n_2854),
.B(n_2800),
.Y(n_2877)
);

NOR2x1_ASAP7_75t_R g2878 ( 
.A(n_2845),
.B(n_2798),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2840),
.B(n_2779),
.Y(n_2879)
);

INVx3_ASAP7_75t_L g2880 ( 
.A(n_2833),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2838),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2827),
.Y(n_2882)
);

INVx3_ASAP7_75t_L g2883 ( 
.A(n_2833),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2840),
.B(n_2837),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2829),
.B(n_2801),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2818),
.Y(n_2886)
);

INVx3_ASAP7_75t_L g2887 ( 
.A(n_2845),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2827),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2853),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2853),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2858),
.Y(n_2891)
);

INVx2_ASAP7_75t_SL g2892 ( 
.A(n_2866),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2861),
.B(n_2845),
.Y(n_2893)
);

OR2x2_ASAP7_75t_L g2894 ( 
.A(n_2860),
.B(n_2845),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2856),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2857),
.B(n_2830),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2856),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2886),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2857),
.B(n_2819),
.Y(n_2899)
);

AND2x4_ASAP7_75t_L g2900 ( 
.A(n_2880),
.B(n_2844),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2866),
.B(n_2798),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2869),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2869),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2871),
.B(n_2820),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2886),
.Y(n_2905)
);

OR2x2_ASAP7_75t_L g2906 ( 
.A(n_2855),
.B(n_2822),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2859),
.B(n_2844),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2871),
.Y(n_2908)
);

NOR2x1_ASAP7_75t_L g2909 ( 
.A(n_2875),
.B(n_2835),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2859),
.B(n_2779),
.Y(n_2910)
);

OR2x2_ASAP7_75t_L g2911 ( 
.A(n_2872),
.B(n_2817),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2889),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2889),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2880),
.B(n_2801),
.Y(n_2914)
);

NAND2x1p5_ASAP7_75t_L g2915 ( 
.A(n_2880),
.B(n_2834),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2872),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2883),
.B(n_2821),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2883),
.B(n_2823),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2863),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2883),
.B(n_2831),
.Y(n_2920)
);

INVx2_ASAP7_75t_SL g2921 ( 
.A(n_2875),
.Y(n_2921)
);

NAND4xp25_ASAP7_75t_L g2922 ( 
.A(n_2884),
.B(n_2820),
.C(n_2851),
.D(n_2847),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2874),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2884),
.B(n_2834),
.Y(n_2924)
);

HB1xp67_ASAP7_75t_L g2925 ( 
.A(n_2887),
.Y(n_2925)
);

OR2x2_ASAP7_75t_L g2926 ( 
.A(n_2885),
.B(n_2799),
.Y(n_2926)
);

AOI21xp5_ASAP7_75t_L g2927 ( 
.A1(n_2862),
.A2(n_2847),
.B(n_2835),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2867),
.B(n_2865),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2887),
.B(n_2841),
.Y(n_2929)
);

INVxp33_ASAP7_75t_L g2930 ( 
.A(n_2878),
.Y(n_2930)
);

HB1xp67_ASAP7_75t_L g2931 ( 
.A(n_2887),
.Y(n_2931)
);

AND2x4_ASAP7_75t_SL g2932 ( 
.A(n_2865),
.B(n_2661),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2867),
.B(n_2848),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2890),
.Y(n_2934)
);

OR2x2_ASAP7_75t_L g2935 ( 
.A(n_2874),
.B(n_2799),
.Y(n_2935)
);

NOR2x1p5_ASAP7_75t_L g2936 ( 
.A(n_2879),
.B(n_2661),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2879),
.B(n_2675),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2932),
.B(n_2675),
.Y(n_2938)
);

AOI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2927),
.A2(n_2864),
.B1(n_2841),
.B2(n_2799),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2932),
.B(n_2868),
.Y(n_2940)
);

INVxp67_ASAP7_75t_L g2941 ( 
.A(n_2901),
.Y(n_2941)
);

NAND3xp33_ASAP7_75t_L g2942 ( 
.A(n_2909),
.B(n_2890),
.C(n_2873),
.Y(n_2942)
);

INVx5_ASAP7_75t_L g2943 ( 
.A(n_2892),
.Y(n_2943)
);

XNOR2xp5_ASAP7_75t_L g2944 ( 
.A(n_2936),
.B(n_2881),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2912),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2912),
.Y(n_2946)
);

NOR2xp33_ASAP7_75t_L g2947 ( 
.A(n_2892),
.B(n_2877),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2907),
.B(n_2877),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2921),
.B(n_2870),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2915),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2901),
.B(n_2876),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2908),
.B(n_2882),
.Y(n_2952)
);

XNOR2x1_ASAP7_75t_L g2953 ( 
.A(n_2904),
.B(n_2888),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2908),
.B(n_2923),
.Y(n_2954)
);

NAND3xp33_ASAP7_75t_SL g2955 ( 
.A(n_2927),
.B(n_2926),
.C(n_2929),
.Y(n_2955)
);

AND2x4_ASAP7_75t_L g2956 ( 
.A(n_2900),
.B(n_2937),
.Y(n_2956)
);

AOI22xp5_ASAP7_75t_L g2957 ( 
.A1(n_2922),
.A2(n_2849),
.B1(n_2788),
.B2(n_2716),
.Y(n_2957)
);

XNOR2xp5_ASAP7_75t_L g2958 ( 
.A(n_2928),
.B(n_2725),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2900),
.B(n_2910),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2900),
.B(n_2788),
.Y(n_2960)
);

INVx2_ASAP7_75t_SL g2961 ( 
.A(n_2914),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2915),
.Y(n_2962)
);

BUFx2_ASAP7_75t_L g2963 ( 
.A(n_2917),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2930),
.B(n_1125),
.Y(n_2964)
);

NAND4xp75_ASAP7_75t_L g2965 ( 
.A(n_2899),
.B(n_2719),
.C(n_11),
.D(n_9),
.Y(n_2965)
);

XNOR2x2_ASAP7_75t_L g2966 ( 
.A(n_2896),
.B(n_10),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2902),
.Y(n_2967)
);

XNOR2xp5_ASAP7_75t_L g2968 ( 
.A(n_2930),
.B(n_11),
.Y(n_2968)
);

XNOR2xp5_ASAP7_75t_L g2969 ( 
.A(n_2893),
.B(n_12),
.Y(n_2969)
);

INVxp67_ASAP7_75t_L g2970 ( 
.A(n_2918),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2925),
.Y(n_2971)
);

HB1xp67_ASAP7_75t_L g2972 ( 
.A(n_2925),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2903),
.B(n_1131),
.Y(n_2973)
);

NAND4xp75_ASAP7_75t_L g2974 ( 
.A(n_2920),
.B(n_14),
.C(n_12),
.D(n_13),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2933),
.B(n_2894),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2913),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2913),
.Y(n_2977)
);

NOR3xp33_ASAP7_75t_L g2978 ( 
.A(n_2924),
.B(n_1138),
.C(n_1133),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2934),
.Y(n_2979)
);

NAND4xp75_ASAP7_75t_L g2980 ( 
.A(n_2934),
.B(n_16),
.C(n_13),
.D(n_15),
.Y(n_2980)
);

AO22x2_ASAP7_75t_L g2981 ( 
.A1(n_2895),
.A2(n_2659),
.B1(n_19),
.B2(n_16),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2931),
.Y(n_2982)
);

NAND4xp75_ASAP7_75t_L g2983 ( 
.A(n_2895),
.B(n_20),
.C(n_18),
.D(n_19),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2931),
.B(n_18),
.Y(n_2984)
);

INVx2_ASAP7_75t_SL g2985 ( 
.A(n_2911),
.Y(n_2985)
);

INVx2_ASAP7_75t_SL g2986 ( 
.A(n_2891),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2916),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2897),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2897),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2906),
.B(n_1142),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2919),
.B(n_1144),
.Y(n_2991)
);

NAND4xp75_ASAP7_75t_L g2992 ( 
.A(n_2898),
.B(n_2905),
.C(n_2935),
.D(n_22),
.Y(n_2992)
);

XOR2x2_ASAP7_75t_L g2993 ( 
.A(n_2898),
.B(n_20),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2905),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2892),
.B(n_1153),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2927),
.A2(n_1212),
.B1(n_1215),
.B2(n_1207),
.Y(n_2996)
);

BUFx2_ASAP7_75t_L g2997 ( 
.A(n_2900),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2923),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2912),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2892),
.B(n_1154),
.Y(n_3000)
);

AND2x4_ASAP7_75t_L g3001 ( 
.A(n_2932),
.B(n_21),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2892),
.B(n_1155),
.Y(n_3002)
);

NAND4xp75_ASAP7_75t_L g3003 ( 
.A(n_2927),
.B(n_24),
.C(n_22),
.D(n_23),
.Y(n_3003)
);

NOR2x1p5_ASAP7_75t_L g3004 ( 
.A(n_2896),
.B(n_1157),
.Y(n_3004)
);

NAND3xp33_ASAP7_75t_L g3005 ( 
.A(n_2909),
.B(n_1161),
.C(n_1159),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2984),
.B(n_1163),
.Y(n_3006)
);

AND2x2_ASAP7_75t_SL g3007 ( 
.A(n_2997),
.B(n_25),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2963),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2972),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2943),
.B(n_2948),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_3001),
.Y(n_3011)
);

A2O1A1O1Ixp25_ASAP7_75t_L g3012 ( 
.A1(n_2966),
.A2(n_1170),
.B(n_1171),
.C(n_1165),
.D(n_1164),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2971),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2982),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2943),
.B(n_2947),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2945),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2943),
.B(n_2996),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_2959),
.B(n_1172),
.Y(n_3018)
);

AND2x2_ASAP7_75t_L g3019 ( 
.A(n_2956),
.B(n_1174),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2946),
.Y(n_3020)
);

AND2x4_ASAP7_75t_L g3021 ( 
.A(n_2956),
.B(n_25),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2975),
.B(n_1175),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2961),
.B(n_1176),
.Y(n_3023)
);

NOR2x1_ASAP7_75t_L g3024 ( 
.A(n_3005),
.B(n_27),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2976),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2977),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2970),
.B(n_1177),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2979),
.Y(n_3028)
);

NAND2x1_ASAP7_75t_L g3029 ( 
.A(n_2950),
.B(n_2962),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2941),
.B(n_2985),
.Y(n_3030)
);

INVx1_ASAP7_75t_SL g3031 ( 
.A(n_3001),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2938),
.B(n_1179),
.Y(n_3032)
);

INVxp67_ASAP7_75t_SL g3033 ( 
.A(n_2968),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2992),
.B(n_1180),
.Y(n_3034)
);

HB1xp67_ASAP7_75t_L g3035 ( 
.A(n_2969),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2999),
.Y(n_3036)
);

AND2x2_ASAP7_75t_L g3037 ( 
.A(n_2940),
.B(n_1183),
.Y(n_3037)
);

OR2x2_ASAP7_75t_L g3038 ( 
.A(n_2955),
.B(n_28),
.Y(n_3038)
);

OR2x2_ASAP7_75t_L g3039 ( 
.A(n_2954),
.B(n_28),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_2951),
.B(n_1191),
.Y(n_3040)
);

AND2x2_ASAP7_75t_L g3041 ( 
.A(n_2964),
.B(n_1192),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2995),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_3000),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_3002),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2981),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2978),
.B(n_1196),
.Y(n_3046)
);

AOI21x1_ASAP7_75t_L g3047 ( 
.A1(n_2993),
.A2(n_38),
.B(n_29),
.Y(n_3047)
);

AOI22xp5_ASAP7_75t_L g3048 ( 
.A1(n_2939),
.A2(n_1202),
.B1(n_1221),
.B2(n_1199),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_3003),
.B(n_1229),
.Y(n_3049)
);

INVx2_ASAP7_75t_SL g3050 ( 
.A(n_2944),
.Y(n_3050)
);

INVx2_ASAP7_75t_SL g3051 ( 
.A(n_2958),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2998),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2952),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2990),
.B(n_1258),
.Y(n_3054)
);

OAI21xp33_ASAP7_75t_L g3055 ( 
.A1(n_2949),
.A2(n_1262),
.B(n_1260),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2998),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2967),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2942),
.B(n_1264),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2981),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2967),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2960),
.B(n_1265),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2991),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2973),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2987),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2974),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2986),
.Y(n_3066)
);

AND2x4_ASAP7_75t_SL g3067 ( 
.A(n_2988),
.B(n_29),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_SL g3068 ( 
.A(n_2980),
.B(n_30),
.Y(n_3068)
);

NAND2xp33_ASAP7_75t_L g3069 ( 
.A(n_3004),
.B(n_30),
.Y(n_3069)
);

AND2x4_ASAP7_75t_L g3070 ( 
.A(n_2989),
.B(n_31),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2953),
.B(n_31),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2983),
.B(n_33),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2965),
.B(n_2957),
.Y(n_3073)
);

NOR2xp67_ASAP7_75t_L g3074 ( 
.A(n_2994),
.B(n_33),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2972),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_2959),
.B(n_34),
.Y(n_3076)
);

OR2x2_ASAP7_75t_L g3077 ( 
.A(n_2985),
.B(n_35),
.Y(n_3077)
);

INVx2_ASAP7_75t_SL g3078 ( 
.A(n_2943),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2997),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2984),
.B(n_35),
.Y(n_3080)
);

OR2x2_ASAP7_75t_L g3081 ( 
.A(n_2985),
.B(n_36),
.Y(n_3081)
);

INVx2_ASAP7_75t_SL g3082 ( 
.A(n_2943),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2984),
.B(n_36),
.Y(n_3083)
);

INVxp67_ASAP7_75t_L g3084 ( 
.A(n_2997),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2984),
.B(n_37),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2972),
.Y(n_3086)
);

INVx4_ASAP7_75t_L g3087 ( 
.A(n_3001),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2984),
.B(n_37),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2959),
.B(n_38),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2972),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2972),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_2959),
.B(n_39),
.Y(n_3092)
);

INVxp67_ASAP7_75t_L g3093 ( 
.A(n_2997),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2972),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2972),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2984),
.B(n_39),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2972),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_2959),
.B(n_40),
.Y(n_3098)
);

NAND3xp33_ASAP7_75t_L g3099 ( 
.A(n_3012),
.B(n_40),
.C(n_41),
.Y(n_3099)
);

OR2x2_ASAP7_75t_L g3100 ( 
.A(n_3079),
.B(n_42),
.Y(n_3100)
);

NAND3xp33_ASAP7_75t_L g3101 ( 
.A(n_3038),
.B(n_43),
.C(n_44),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_3007),
.B(n_44),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3008),
.Y(n_3103)
);

XOR2x2_ASAP7_75t_L g3104 ( 
.A(n_3050),
.B(n_46),
.Y(n_3104)
);

OAI21xp33_ASAP7_75t_L g3105 ( 
.A1(n_3048),
.A2(n_45),
.B(n_46),
.Y(n_3105)
);

OAI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_3071),
.A2(n_45),
.B(n_47),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_3039),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_3033),
.Y(n_3108)
);

OAI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_3068),
.A2(n_2659),
.B1(n_51),
.B2(n_49),
.Y(n_3109)
);

AOI22xp5_ASAP7_75t_L g3110 ( 
.A1(n_3073),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_3110)
);

A2O1A1Ixp33_ASAP7_75t_L g3111 ( 
.A1(n_3058),
.A2(n_53),
.B(n_50),
.C(n_52),
.Y(n_3111)
);

NOR3xp33_ASAP7_75t_L g3112 ( 
.A(n_3035),
.B(n_54),
.C(n_55),
.Y(n_3112)
);

INVxp67_ASAP7_75t_L g3113 ( 
.A(n_3076),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_3045),
.A2(n_1457),
.B1(n_1423),
.B2(n_57),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_3080),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_3083),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_3085),
.Y(n_3117)
);

NAND3xp33_ASAP7_75t_L g3118 ( 
.A(n_3084),
.B(n_54),
.C(n_56),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_3088),
.Y(n_3119)
);

OAI21xp5_ASAP7_75t_SL g3120 ( 
.A1(n_3093),
.A2(n_56),
.B(n_57),
.Y(n_3120)
);

AOI21xp33_ASAP7_75t_SL g3121 ( 
.A1(n_3011),
.A2(n_59),
.B(n_60),
.Y(n_3121)
);

AO21x1_ASAP7_75t_SL g3122 ( 
.A1(n_3010),
.A2(n_68),
.B(n_59),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_3087),
.B(n_60),
.Y(n_3123)
);

XNOR2xp5_ASAP7_75t_L g3124 ( 
.A(n_3047),
.B(n_61),
.Y(n_3124)
);

INVx2_ASAP7_75t_SL g3125 ( 
.A(n_3021),
.Y(n_3125)
);

INVxp67_ASAP7_75t_L g3126 ( 
.A(n_3089),
.Y(n_3126)
);

AOI22xp33_ASAP7_75t_L g3127 ( 
.A1(n_3059),
.A2(n_1457),
.B1(n_63),
.B2(n_61),
.Y(n_3127)
);

OAI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_3031),
.A2(n_66),
.B1(n_62),
.B2(n_65),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_3034),
.A2(n_65),
.B(n_66),
.Y(n_3129)
);

AOI211xp5_ASAP7_75t_L g3130 ( 
.A1(n_3017),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_3130)
);

OR4x1_ASAP7_75t_L g3131 ( 
.A(n_3078),
.B(n_70),
.C(n_67),
.D(n_69),
.Y(n_3131)
);

OAI22xp33_ASAP7_75t_SL g3132 ( 
.A1(n_3029),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_3096),
.Y(n_3133)
);

OAI31xp33_ASAP7_75t_L g3134 ( 
.A1(n_3064),
.A2(n_3037),
.A3(n_3065),
.B(n_3052),
.Y(n_3134)
);

OAI21xp5_ASAP7_75t_L g3135 ( 
.A1(n_3015),
.A2(n_72),
.B(n_73),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3009),
.Y(n_3136)
);

OAI31xp33_ASAP7_75t_L g3137 ( 
.A1(n_3052),
.A2(n_78),
.A3(n_74),
.B(n_75),
.Y(n_3137)
);

NAND3xp33_ASAP7_75t_L g3138 ( 
.A(n_3087),
.B(n_78),
.C(n_79),
.Y(n_3138)
);

INVxp67_ASAP7_75t_SL g3139 ( 
.A(n_3006),
.Y(n_3139)
);

NAND2x1_ASAP7_75t_L g3140 ( 
.A(n_3082),
.B(n_80),
.Y(n_3140)
);

OAI22xp5_ASAP7_75t_L g3141 ( 
.A1(n_3030),
.A2(n_85),
.B1(n_81),
.B2(n_82),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3009),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3095),
.Y(n_3143)
);

INVxp67_ASAP7_75t_SL g3144 ( 
.A(n_3022),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_3021),
.Y(n_3145)
);

XOR2x2_ASAP7_75t_L g3146 ( 
.A(n_3024),
.B(n_85),
.Y(n_3146)
);

OAI21xp33_ASAP7_75t_L g3147 ( 
.A1(n_3066),
.A2(n_82),
.B(n_86),
.Y(n_3147)
);

INVx3_ASAP7_75t_L g3148 ( 
.A(n_3092),
.Y(n_3148)
);

AOI22xp5_ASAP7_75t_L g3149 ( 
.A1(n_3069),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_3095),
.Y(n_3150)
);

OAI221xp5_ASAP7_75t_L g3151 ( 
.A1(n_3077),
.A2(n_3081),
.B1(n_3063),
.B2(n_3062),
.C(n_3044),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_3042),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3097),
.Y(n_3153)
);

AND2x4_ASAP7_75t_L g3154 ( 
.A(n_3098),
.B(n_3013),
.Y(n_3154)
);

AO22x1_ASAP7_75t_L g3155 ( 
.A1(n_3018),
.A2(n_98),
.B1(n_109),
.B2(n_89),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3097),
.Y(n_3156)
);

AOI21xp33_ASAP7_75t_L g3157 ( 
.A1(n_3053),
.A2(n_91),
.B(n_92),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_3072),
.A2(n_93),
.B(n_94),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_3070),
.Y(n_3159)
);

AOI22xp5_ASAP7_75t_L g3160 ( 
.A1(n_3043),
.A2(n_96),
.B1(n_93),
.B2(n_95),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_3070),
.Y(n_3161)
);

AOI22xp5_ASAP7_75t_SL g3162 ( 
.A1(n_3019),
.A2(n_99),
.B1(n_95),
.B2(n_97),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_3075),
.Y(n_3163)
);

NOR3xp33_ASAP7_75t_L g3164 ( 
.A(n_3055),
.B(n_97),
.C(n_100),
.Y(n_3164)
);

OAI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_3014),
.A2(n_3051),
.B(n_3040),
.Y(n_3165)
);

OAI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_3086),
.A2(n_100),
.B(n_102),
.Y(n_3166)
);

AOI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_3049),
.A2(n_102),
.B(n_103),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_3027),
.A2(n_105),
.B(n_106),
.Y(n_3168)
);

AOI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_3061),
.A2(n_106),
.B(n_108),
.Y(n_3169)
);

INVxp33_ASAP7_75t_L g3170 ( 
.A(n_3032),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3090),
.Y(n_3171)
);

OAI22xp5_ASAP7_75t_L g3172 ( 
.A1(n_3091),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_3172)
);

AOI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_3041),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_3173)
);

XNOR2x1_ASAP7_75t_L g3174 ( 
.A(n_3074),
.B(n_113),
.Y(n_3174)
);

NAND2xp33_ASAP7_75t_L g3175 ( 
.A(n_3023),
.B(n_112),
.Y(n_3175)
);

AOI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_3054),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_3067),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_3056),
.A2(n_3060),
.B(n_3057),
.Y(n_3178)
);

INVx1_ASAP7_75t_SL g3179 ( 
.A(n_3046),
.Y(n_3179)
);

NOR3xp33_ASAP7_75t_L g3180 ( 
.A(n_3016),
.B(n_114),
.C(n_115),
.Y(n_3180)
);

AOI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_3020),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_3181)
);

O2A1O1Ixp33_ASAP7_75t_L g3182 ( 
.A1(n_3094),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_3182)
);

AOI22xp5_ASAP7_75t_L g3183 ( 
.A1(n_3025),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_3026),
.Y(n_3184)
);

OAI211xp5_ASAP7_75t_L g3185 ( 
.A1(n_3028),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_3185)
);

NAND3xp33_ASAP7_75t_SL g3186 ( 
.A(n_3036),
.B(n_124),
.C(n_125),
.Y(n_3186)
);

AO22x1_ASAP7_75t_L g3187 ( 
.A1(n_3011),
.A2(n_132),
.B1(n_142),
.B2(n_124),
.Y(n_3187)
);

INVxp67_ASAP7_75t_L g3188 ( 
.A(n_3068),
.Y(n_3188)
);

INVxp67_ASAP7_75t_L g3189 ( 
.A(n_3068),
.Y(n_3189)
);

XOR2x2_ASAP7_75t_L g3190 ( 
.A(n_3050),
.B(n_126),
.Y(n_3190)
);

INVx1_ASAP7_75t_SL g3191 ( 
.A(n_3011),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3079),
.Y(n_3192)
);

OAI31xp33_ASAP7_75t_L g3193 ( 
.A1(n_3073),
.A2(n_127),
.A3(n_125),
.B(n_126),
.Y(n_3193)
);

NOR3xp33_ASAP7_75t_L g3194 ( 
.A(n_3050),
.B(n_128),
.C(n_129),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_3079),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_3007),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3079),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_3076),
.B(n_128),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3079),
.Y(n_3199)
);

OAI31xp33_ASAP7_75t_L g3200 ( 
.A1(n_3073),
.A2(n_131),
.A3(n_129),
.B(n_130),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_3079),
.Y(n_3201)
);

OR2x2_ASAP7_75t_L g3202 ( 
.A(n_3079),
.B(n_131),
.Y(n_3202)
);

OAI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_3012),
.A2(n_133),
.B(n_134),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3079),
.Y(n_3204)
);

OAI221xp5_ASAP7_75t_L g3205 ( 
.A1(n_3048),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.C(n_136),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3079),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3079),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3007),
.B(n_137),
.Y(n_3208)
);

XNOR2xp5_ASAP7_75t_L g3209 ( 
.A(n_3011),
.B(n_138),
.Y(n_3209)
);

CKINVDCx5p33_ASAP7_75t_R g3210 ( 
.A(n_3011),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_3071),
.A2(n_138),
.B(n_139),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3079),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3079),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3079),
.Y(n_3214)
);

INVx2_ASAP7_75t_SL g3215 ( 
.A(n_3011),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3079),
.Y(n_3216)
);

OAI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_3012),
.A2(n_143),
.B(n_144),
.Y(n_3217)
);

INVx2_ASAP7_75t_SL g3218 ( 
.A(n_3011),
.Y(n_3218)
);

NAND4xp25_ASAP7_75t_L g3219 ( 
.A(n_3030),
.B(n_145),
.C(n_143),
.D(n_144),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3079),
.Y(n_3220)
);

INVx3_ASAP7_75t_L g3221 ( 
.A(n_3087),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_SL g3222 ( 
.A(n_3011),
.B(n_146),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_3076),
.B(n_146),
.Y(n_3223)
);

INVx3_ASAP7_75t_L g3224 ( 
.A(n_3087),
.Y(n_3224)
);

OAI21xp33_ASAP7_75t_SL g3225 ( 
.A1(n_3048),
.A2(n_147),
.B(n_148),
.Y(n_3225)
);

OAI22xp5_ASAP7_75t_SL g3226 ( 
.A1(n_3011),
.A2(n_156),
.B1(n_167),
.B2(n_147),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3007),
.B(n_148),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3079),
.Y(n_3228)
);

OAI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_3048),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_3229)
);

INVxp67_ASAP7_75t_SL g3230 ( 
.A(n_3050),
.Y(n_3230)
);

NAND3xp33_ASAP7_75t_SL g3231 ( 
.A(n_3048),
.B(n_149),
.C(n_152),
.Y(n_3231)
);

OAI21xp33_ASAP7_75t_L g3232 ( 
.A1(n_3050),
.A2(n_152),
.B(n_153),
.Y(n_3232)
);

OR2x2_ASAP7_75t_L g3233 ( 
.A(n_3079),
.B(n_153),
.Y(n_3233)
);

INVx1_ASAP7_75t_SL g3234 ( 
.A(n_3011),
.Y(n_3234)
);

NOR2xp33_ASAP7_75t_L g3235 ( 
.A(n_3087),
.B(n_154),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3079),
.Y(n_3236)
);

AO22x1_ASAP7_75t_L g3237 ( 
.A1(n_3011),
.A2(n_165),
.B1(n_176),
.B2(n_154),
.Y(n_3237)
);

OAI21xp33_ASAP7_75t_L g3238 ( 
.A1(n_3050),
.A2(n_156),
.B(n_157),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3079),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3079),
.Y(n_3240)
);

XOR2x2_ASAP7_75t_L g3241 ( 
.A(n_3050),
.B(n_159),
.Y(n_3241)
);

OAI22xp5_ASAP7_75t_L g3242 ( 
.A1(n_3011),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_3242)
);

NAND3xp33_ASAP7_75t_SL g3243 ( 
.A(n_3048),
.B(n_160),
.C(n_162),
.Y(n_3243)
);

AOI21xp33_ASAP7_75t_L g3244 ( 
.A1(n_3029),
.A2(n_162),
.B(n_163),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3079),
.Y(n_3245)
);

NOR3xp33_ASAP7_75t_L g3246 ( 
.A(n_3050),
.B(n_163),
.C(n_165),
.Y(n_3246)
);

OAI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_3012),
.A2(n_167),
.B(n_168),
.Y(n_3247)
);

NAND3xp33_ASAP7_75t_SL g3248 ( 
.A(n_3048),
.B(n_168),
.C(n_170),
.Y(n_3248)
);

OAI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_3012),
.A2(n_170),
.B(n_171),
.Y(n_3249)
);

INVxp67_ASAP7_75t_L g3250 ( 
.A(n_3068),
.Y(n_3250)
);

AOI21xp33_ASAP7_75t_L g3251 ( 
.A1(n_3029),
.A2(n_173),
.B(n_174),
.Y(n_3251)
);

OAI211xp5_ASAP7_75t_L g3252 ( 
.A1(n_3048),
.A2(n_176),
.B(n_173),
.C(n_175),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3079),
.Y(n_3253)
);

INVx1_ASAP7_75t_SL g3254 ( 
.A(n_3210),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3187),
.B(n_175),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_3131),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_3148),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3230),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3209),
.Y(n_3259)
);

AOI22xp5_ASAP7_75t_L g3260 ( 
.A1(n_3144),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_3260)
);

OR2x2_ASAP7_75t_L g3261 ( 
.A(n_3191),
.B(n_177),
.Y(n_3261)
);

OAI221xp5_ASAP7_75t_L g3262 ( 
.A1(n_3134),
.A2(n_3196),
.B1(n_3244),
.B2(n_3251),
.C(n_3151),
.Y(n_3262)
);

NAND3xp33_ASAP7_75t_L g3263 ( 
.A(n_3188),
.B(n_178),
.C(n_179),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_3148),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3234),
.B(n_180),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3198),
.Y(n_3266)
);

OAI22xp33_ASAP7_75t_L g3267 ( 
.A1(n_3170),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3223),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_3215),
.B(n_181),
.Y(n_3269)
);

OAI221xp5_ASAP7_75t_L g3270 ( 
.A1(n_3113),
.A2(n_3126),
.B1(n_3250),
.B2(n_3189),
.C(n_3139),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_3237),
.B(n_3155),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_SL g3272 ( 
.A(n_3132),
.B(n_182),
.Y(n_3272)
);

OAI21xp33_ASAP7_75t_L g3273 ( 
.A1(n_3218),
.A2(n_185),
.B(n_186),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3124),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_3221),
.B(n_187),
.Y(n_3275)
);

INVx1_ASAP7_75t_SL g3276 ( 
.A(n_3104),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3221),
.B(n_3224),
.Y(n_3277)
);

INVx1_ASAP7_75t_SL g3278 ( 
.A(n_3190),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3140),
.Y(n_3279)
);

NOR2xp33_ASAP7_75t_L g3280 ( 
.A(n_3121),
.B(n_187),
.Y(n_3280)
);

AOI22xp5_ASAP7_75t_L g3281 ( 
.A1(n_3146),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_3281)
);

OAI322xp33_ASAP7_75t_L g3282 ( 
.A1(n_3136),
.A2(n_195),
.A3(n_194),
.B1(n_192),
.B2(n_189),
.C1(n_190),
.C2(n_193),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3241),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3154),
.B(n_193),
.Y(n_3284)
);

AOI21xp33_ASAP7_75t_SL g3285 ( 
.A1(n_3123),
.A2(n_197),
.B(n_198),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3154),
.B(n_3125),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3162),
.B(n_3145),
.Y(n_3287)
);

OAI32xp33_ASAP7_75t_L g3288 ( 
.A1(n_3192),
.A2(n_201),
.A3(n_198),
.B1(n_199),
.B2(n_202),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3226),
.Y(n_3289)
);

O2A1O1Ixp33_ASAP7_75t_L g3290 ( 
.A1(n_3120),
.A2(n_206),
.B(n_203),
.C(n_204),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3174),
.Y(n_3291)
);

OAI21xp33_ASAP7_75t_SL g3292 ( 
.A1(n_3142),
.A2(n_203),
.B(n_207),
.Y(n_3292)
);

NOR3xp33_ASAP7_75t_L g3293 ( 
.A(n_3165),
.B(n_207),
.C(n_208),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3159),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3161),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3107),
.Y(n_3296)
);

AOI22xp33_ASAP7_75t_L g3297 ( 
.A1(n_3179),
.A2(n_212),
.B1(n_208),
.B2(n_211),
.Y(n_3297)
);

AOI22xp5_ASAP7_75t_L g3298 ( 
.A1(n_3225),
.A2(n_215),
.B1(n_211),
.B2(n_214),
.Y(n_3298)
);

O2A1O1Ixp33_ASAP7_75t_SL g3299 ( 
.A1(n_3195),
.A2(n_218),
.B(n_214),
.C(n_217),
.Y(n_3299)
);

AOI221xp5_ASAP7_75t_L g3300 ( 
.A1(n_3158),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.C(n_220),
.Y(n_3300)
);

NAND3xp33_ASAP7_75t_L g3301 ( 
.A(n_3194),
.B(n_219),
.C(n_220),
.Y(n_3301)
);

O2A1O1Ixp5_ASAP7_75t_L g3302 ( 
.A1(n_3224),
.A2(n_224),
.B(n_221),
.C(n_222),
.Y(n_3302)
);

OAI221xp5_ASAP7_75t_L g3303 ( 
.A1(n_3101),
.A2(n_226),
.B1(n_222),
.B2(n_224),
.C(n_227),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3100),
.Y(n_3304)
);

OAI21xp33_ASAP7_75t_L g3305 ( 
.A1(n_3108),
.A2(n_226),
.B(n_227),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3202),
.Y(n_3306)
);

OAI22xp33_ASAP7_75t_L g3307 ( 
.A1(n_3110),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_3307)
);

OAI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_3178),
.A2(n_228),
.B(n_231),
.Y(n_3308)
);

OAI32xp33_ASAP7_75t_L g3309 ( 
.A1(n_3197),
.A2(n_234),
.A3(n_232),
.B1(n_233),
.B2(n_235),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3233),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3246),
.B(n_232),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3102),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3208),
.Y(n_3313)
);

INVxp67_ASAP7_75t_SL g3314 ( 
.A(n_3222),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_3199),
.B(n_233),
.Y(n_3315)
);

INVxp67_ASAP7_75t_SL g3316 ( 
.A(n_3227),
.Y(n_3316)
);

AOI33xp33_ASAP7_75t_L g3317 ( 
.A1(n_3201),
.A2(n_236),
.A3(n_238),
.B1(n_234),
.B2(n_235),
.B3(n_237),
.Y(n_3317)
);

OAI22xp33_ASAP7_75t_L g3318 ( 
.A1(n_3149),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_3318)
);

BUFx2_ASAP7_75t_L g3319 ( 
.A(n_3135),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3099),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3204),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3177),
.Y(n_3322)
);

OAI22xp5_ASAP7_75t_L g3323 ( 
.A1(n_3206),
.A2(n_242),
.B1(n_239),
.B2(n_240),
.Y(n_3323)
);

AOI21xp33_ASAP7_75t_L g3324 ( 
.A1(n_3115),
.A2(n_239),
.B(n_242),
.Y(n_3324)
);

AOI211xp5_ASAP7_75t_L g3325 ( 
.A1(n_3207),
.A2(n_245),
.B(n_243),
.C(n_244),
.Y(n_3325)
);

INVxp33_ASAP7_75t_L g3326 ( 
.A(n_3219),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3212),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3116),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3211),
.B(n_244),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3213),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3214),
.Y(n_3331)
);

AOI21xp5_ASAP7_75t_L g3332 ( 
.A1(n_3186),
.A2(n_245),
.B(n_246),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3216),
.B(n_246),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3220),
.Y(n_3334)
);

NOR2xp33_ASAP7_75t_L g3335 ( 
.A(n_3232),
.B(n_247),
.Y(n_3335)
);

INVx3_ASAP7_75t_L g3336 ( 
.A(n_3228),
.Y(n_3336)
);

AOI222xp33_ASAP7_75t_L g3337 ( 
.A1(n_3143),
.A2(n_3153),
.B1(n_3156),
.B2(n_3150),
.C1(n_3184),
.C2(n_3133),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3175),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3236),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3239),
.Y(n_3340)
);

NOR2x1_ASAP7_75t_L g3341 ( 
.A(n_3138),
.B(n_248),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3240),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3245),
.Y(n_3343)
);

OAI21xp5_ASAP7_75t_SL g3344 ( 
.A1(n_3253),
.A2(n_249),
.B(n_250),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3235),
.B(n_251),
.Y(n_3345)
);

AOI221xp5_ASAP7_75t_L g3346 ( 
.A1(n_3117),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.C(n_255),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3119),
.Y(n_3347)
);

OAI21xp33_ASAP7_75t_L g3348 ( 
.A1(n_3103),
.A2(n_256),
.B(n_257),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3130),
.B(n_257),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3203),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3217),
.Y(n_3351)
);

OAI32xp33_ASAP7_75t_L g3352 ( 
.A1(n_3180),
.A2(n_260),
.A3(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_3352)
);

AOI22xp5_ASAP7_75t_L g3353 ( 
.A1(n_3231),
.A2(n_263),
.B1(n_258),
.B2(n_262),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3247),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3249),
.Y(n_3355)
);

AOI22xp5_ASAP7_75t_L g3356 ( 
.A1(n_3243),
.A2(n_265),
.B1(n_262),
.B2(n_264),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3185),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3128),
.Y(n_3358)
);

AOI22xp5_ASAP7_75t_L g3359 ( 
.A1(n_3248),
.A2(n_268),
.B1(n_264),
.B2(n_266),
.Y(n_3359)
);

INVxp67_ASAP7_75t_L g3360 ( 
.A(n_3122),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3182),
.Y(n_3361)
);

CKINVDCx6p67_ASAP7_75t_R g3362 ( 
.A(n_3163),
.Y(n_3362)
);

AOI221xp5_ASAP7_75t_L g3363 ( 
.A1(n_3114),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.C(n_273),
.Y(n_3363)
);

AOI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_3168),
.A2(n_270),
.B(n_274),
.Y(n_3364)
);

OAI221xp5_ASAP7_75t_L g3365 ( 
.A1(n_3127),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_3365)
);

INVx1_ASAP7_75t_SL g3366 ( 
.A(n_3169),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3112),
.B(n_275),
.Y(n_3367)
);

AND2x4_ASAP7_75t_L g3368 ( 
.A(n_3171),
.B(n_276),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_3118),
.Y(n_3369)
);

OAI222xp33_ASAP7_75t_L g3370 ( 
.A1(n_3109),
.A2(n_280),
.B1(n_282),
.B2(n_278),
.C1(n_279),
.C2(n_281),
.Y(n_3370)
);

AOI222xp33_ASAP7_75t_L g3371 ( 
.A1(n_3106),
.A2(n_281),
.B1(n_283),
.B2(n_279),
.C1(n_280),
.C2(n_282),
.Y(n_3371)
);

AOI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_3238),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3193),
.B(n_284),
.Y(n_3373)
);

OAI221xp5_ASAP7_75t_L g3374 ( 
.A1(n_3200),
.A2(n_3129),
.B1(n_3167),
.B2(n_3137),
.C(n_3166),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3160),
.Y(n_3375)
);

O2A1O1Ixp5_ASAP7_75t_L g3376 ( 
.A1(n_3157),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_3376)
);

OAI22xp5_ASAP7_75t_L g3377 ( 
.A1(n_3360),
.A2(n_3147),
.B1(n_3183),
.B2(n_3181),
.Y(n_3377)
);

NOR2x1_ASAP7_75t_L g3378 ( 
.A(n_3286),
.B(n_3141),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3254),
.B(n_3164),
.Y(n_3379)
);

OAI31xp33_ASAP7_75t_L g3380 ( 
.A1(n_3262),
.A2(n_3252),
.A3(n_3111),
.B(n_3172),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3317),
.Y(n_3381)
);

NOR2x1_ASAP7_75t_L g3382 ( 
.A(n_3336),
.B(n_3242),
.Y(n_3382)
);

OAI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3256),
.A2(n_3152),
.B1(n_3173),
.B2(n_3176),
.Y(n_3383)
);

NAND2x1_ASAP7_75t_L g3384 ( 
.A(n_3279),
.B(n_3105),
.Y(n_3384)
);

OR2x2_ASAP7_75t_L g3385 ( 
.A(n_3257),
.B(n_3205),
.Y(n_3385)
);

INVxp67_ASAP7_75t_SL g3386 ( 
.A(n_3336),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3261),
.Y(n_3387)
);

AOI222xp33_ASAP7_75t_L g3388 ( 
.A1(n_3366),
.A2(n_3229),
.B1(n_290),
.B2(n_293),
.C1(n_287),
.C2(n_289),
.Y(n_3388)
);

OR2x2_ASAP7_75t_L g3389 ( 
.A(n_3264),
.B(n_290),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3266),
.Y(n_3390)
);

AOI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3350),
.A2(n_295),
.B1(n_291),
.B2(n_293),
.Y(n_3391)
);

OR2x2_ASAP7_75t_L g3392 ( 
.A(n_3258),
.B(n_296),
.Y(n_3392)
);

OAI31xp33_ASAP7_75t_L g3393 ( 
.A1(n_3274),
.A2(n_299),
.A3(n_296),
.B(n_297),
.Y(n_3393)
);

AOI22xp5_ASAP7_75t_L g3394 ( 
.A1(n_3351),
.A2(n_304),
.B1(n_301),
.B2(n_303),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3276),
.B(n_303),
.Y(n_3395)
);

AOI221xp5_ASAP7_75t_L g3396 ( 
.A1(n_3354),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.C(n_308),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3268),
.Y(n_3397)
);

AOI22xp5_ASAP7_75t_L g3398 ( 
.A1(n_3355),
.A2(n_308),
.B1(n_305),
.B2(n_306),
.Y(n_3398)
);

INVxp67_ASAP7_75t_L g3399 ( 
.A(n_3277),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_3315),
.Y(n_3400)
);

AOI22xp5_ASAP7_75t_L g3401 ( 
.A1(n_3316),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3278),
.B(n_309),
.Y(n_3402)
);

OAI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3292),
.A2(n_310),
.B(n_311),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_L g3404 ( 
.A(n_3285),
.B(n_312),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3333),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3368),
.B(n_312),
.Y(n_3406)
);

OAI22xp5_ASAP7_75t_L g3407 ( 
.A1(n_3314),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3368),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3265),
.Y(n_3409)
);

OAI21xp33_ASAP7_75t_L g3410 ( 
.A1(n_3326),
.A2(n_3320),
.B(n_3322),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3285),
.B(n_315),
.Y(n_3411)
);

OAI32xp33_ASAP7_75t_L g3412 ( 
.A1(n_3357),
.A2(n_318),
.A3(n_316),
.B1(n_317),
.B2(n_319),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3284),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3362),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3291),
.Y(n_3415)
);

OAI211xp5_ASAP7_75t_L g3416 ( 
.A1(n_3337),
.A2(n_320),
.B(n_317),
.C(n_319),
.Y(n_3416)
);

OAI221xp5_ASAP7_75t_SL g3417 ( 
.A1(n_3283),
.A2(n_325),
.B1(n_321),
.B2(n_324),
.C(n_326),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3275),
.B(n_321),
.Y(n_3418)
);

OAI21xp33_ASAP7_75t_SL g3419 ( 
.A1(n_3321),
.A2(n_324),
.B(n_325),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3302),
.Y(n_3420)
);

AOI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3312),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_3421)
);

OR2x2_ASAP7_75t_L g3422 ( 
.A(n_3327),
.B(n_329),
.Y(n_3422)
);

OAI21xp5_ASAP7_75t_L g3423 ( 
.A1(n_3341),
.A2(n_330),
.B(n_332),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3329),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3319),
.Y(n_3425)
);

HB1xp67_ASAP7_75t_L g3426 ( 
.A(n_3255),
.Y(n_3426)
);

INVx2_ASAP7_75t_SL g3427 ( 
.A(n_3269),
.Y(n_3427)
);

INVx1_ASAP7_75t_SL g3428 ( 
.A(n_3271),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3296),
.B(n_330),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3304),
.Y(n_3430)
);

AOI31xp33_ASAP7_75t_L g3431 ( 
.A1(n_3330),
.A2(n_335),
.A3(n_333),
.B(n_334),
.Y(n_3431)
);

OAI221xp5_ASAP7_75t_SL g3432 ( 
.A1(n_3270),
.A2(n_336),
.B1(n_333),
.B2(n_334),
.C(n_337),
.Y(n_3432)
);

HB1xp67_ASAP7_75t_L g3433 ( 
.A(n_3259),
.Y(n_3433)
);

INVxp67_ASAP7_75t_SL g3434 ( 
.A(n_3290),
.Y(n_3434)
);

OAI221xp5_ASAP7_75t_L g3435 ( 
.A1(n_3374),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.C(n_339),
.Y(n_3435)
);

OAI21xp33_ASAP7_75t_L g3436 ( 
.A1(n_3358),
.A2(n_338),
.B(n_340),
.Y(n_3436)
);

NAND3xp33_ASAP7_75t_L g3437 ( 
.A(n_3293),
.B(n_340),
.C(n_341),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3344),
.B(n_342),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3306),
.Y(n_3439)
);

INVxp67_ASAP7_75t_L g3440 ( 
.A(n_3280),
.Y(n_3440)
);

NAND2xp33_ASAP7_75t_SL g3441 ( 
.A(n_3331),
.B(n_342),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3310),
.Y(n_3442)
);

OAI31xp33_ASAP7_75t_L g3443 ( 
.A1(n_3361),
.A2(n_345),
.A3(n_343),
.B(n_344),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3287),
.Y(n_3444)
);

OR2x2_ASAP7_75t_L g3445 ( 
.A(n_3334),
.B(n_344),
.Y(n_3445)
);

OAI221xp5_ASAP7_75t_L g3446 ( 
.A1(n_3308),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.C(n_348),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3349),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3313),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3311),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3364),
.B(n_349),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3339),
.B(n_350),
.Y(n_3451)
);

INVx1_ASAP7_75t_SL g3452 ( 
.A(n_3345),
.Y(n_3452)
);

OAI21xp5_ASAP7_75t_SL g3453 ( 
.A1(n_3340),
.A2(n_352),
.B(n_354),
.Y(n_3453)
);

NOR2xp33_ASAP7_75t_L g3454 ( 
.A(n_3299),
.B(n_352),
.Y(n_3454)
);

O2A1O1Ixp5_ASAP7_75t_L g3455 ( 
.A1(n_3342),
.A2(n_357),
.B(n_355),
.C(n_356),
.Y(n_3455)
);

OAI22xp5_ASAP7_75t_L g3456 ( 
.A1(n_3343),
.A2(n_361),
.B1(n_358),
.B2(n_360),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3367),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3376),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3282),
.Y(n_3459)
);

AOI222xp33_ASAP7_75t_L g3460 ( 
.A1(n_3289),
.A2(n_363),
.B1(n_366),
.B2(n_358),
.C1(n_361),
.C2(n_364),
.Y(n_3460)
);

NAND3xp33_ASAP7_75t_L g3461 ( 
.A(n_3325),
.B(n_363),
.C(n_366),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_SL g3462 ( 
.A1(n_3294),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3295),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3373),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3338),
.B(n_367),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3281),
.B(n_3371),
.Y(n_3466)
);

OAI221xp5_ASAP7_75t_SL g3467 ( 
.A1(n_3328),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.C(n_373),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3347),
.Y(n_3468)
);

INVxp67_ASAP7_75t_L g3469 ( 
.A(n_3272),
.Y(n_3469)
);

BUFx2_ASAP7_75t_L g3470 ( 
.A(n_3369),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3260),
.Y(n_3471)
);

OAI221xp5_ASAP7_75t_L g3472 ( 
.A1(n_3332),
.A2(n_3301),
.B1(n_3375),
.B2(n_3300),
.C(n_3348),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3263),
.Y(n_3473)
);

AOI222xp33_ASAP7_75t_L g3474 ( 
.A1(n_3370),
.A2(n_372),
.B1(n_375),
.B2(n_370),
.C1(n_371),
.C2(n_373),
.Y(n_3474)
);

OAI22xp5_ASAP7_75t_L g3475 ( 
.A1(n_3372),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_3475)
);

AOI221xp5_ASAP7_75t_L g3476 ( 
.A1(n_3352),
.A2(n_380),
.B1(n_377),
.B2(n_379),
.C(n_381),
.Y(n_3476)
);

AOI21xp33_ASAP7_75t_L g3477 ( 
.A1(n_3298),
.A2(n_380),
.B(n_382),
.Y(n_3477)
);

INVxp67_ASAP7_75t_L g3478 ( 
.A(n_3335),
.Y(n_3478)
);

NOR3xp33_ASAP7_75t_L g3479 ( 
.A(n_3324),
.B(n_383),
.C(n_384),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3323),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3353),
.B(n_383),
.Y(n_3481)
);

INVxp67_ASAP7_75t_L g3482 ( 
.A(n_3303),
.Y(n_3482)
);

NOR3xp33_ASAP7_75t_L g3483 ( 
.A(n_3305),
.B(n_384),
.C(n_385),
.Y(n_3483)
);

NOR4xp25_ASAP7_75t_SL g3484 ( 
.A(n_3273),
.B(n_391),
.C(n_388),
.D(n_390),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_3356),
.Y(n_3485)
);

NOR2xp33_ASAP7_75t_L g3486 ( 
.A(n_3288),
.B(n_388),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3309),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3359),
.B(n_390),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3267),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3365),
.Y(n_3490)
);

OR2x2_ASAP7_75t_L g3491 ( 
.A(n_3297),
.B(n_392),
.Y(n_3491)
);

A2O1A1Ixp33_ASAP7_75t_L g3492 ( 
.A1(n_3363),
.A2(n_397),
.B(n_394),
.C(n_395),
.Y(n_3492)
);

AND2x2_ASAP7_75t_L g3493 ( 
.A(n_3346),
.B(n_394),
.Y(n_3493)
);

OAI221xp5_ASAP7_75t_L g3494 ( 
.A1(n_3307),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.C(n_400),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3318),
.B(n_399),
.Y(n_3495)
);

HB1xp67_ASAP7_75t_L g3496 ( 
.A(n_3360),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3276),
.B(n_401),
.Y(n_3497)
);

NAND3xp33_ASAP7_75t_L g3498 ( 
.A(n_3337),
.B(n_402),
.C(n_403),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3276),
.B(n_405),
.Y(n_3499)
);

AOI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_3350),
.A2(n_409),
.B1(n_405),
.B2(n_408),
.Y(n_3500)
);

NOR2xp33_ASAP7_75t_L g3501 ( 
.A(n_3360),
.B(n_408),
.Y(n_3501)
);

AOI221xp5_ASAP7_75t_L g3502 ( 
.A1(n_3262),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.C(n_414),
.Y(n_3502)
);

INVxp67_ASAP7_75t_L g3503 ( 
.A(n_3286),
.Y(n_3503)
);

AO21x1_ASAP7_75t_L g3504 ( 
.A1(n_3286),
.A2(n_410),
.B(n_412),
.Y(n_3504)
);

AOI22xp33_ASAP7_75t_SL g3505 ( 
.A1(n_3279),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_3505)
);

OAI221xp5_ASAP7_75t_L g3506 ( 
.A1(n_3292),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.C(n_418),
.Y(n_3506)
);

OR2x2_ASAP7_75t_L g3507 ( 
.A(n_3257),
.B(n_419),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3254),
.B(n_420),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3276),
.B(n_421),
.Y(n_3509)
);

NAND3xp33_ASAP7_75t_SL g3510 ( 
.A(n_3276),
.B(n_421),
.C(n_422),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3276),
.B(n_423),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3299),
.A2(n_424),
.B(n_425),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3276),
.B(n_424),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_L g3514 ( 
.A(n_3360),
.B(n_425),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3317),
.Y(n_3515)
);

NAND3x1_ASAP7_75t_L g3516 ( 
.A(n_3286),
.B(n_426),
.C(n_427),
.Y(n_3516)
);

AOI211xp5_ASAP7_75t_L g3517 ( 
.A1(n_3360),
.A2(n_429),
.B(n_427),
.C(n_428),
.Y(n_3517)
);

OAI22xp33_ASAP7_75t_L g3518 ( 
.A1(n_3279),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_3518)
);

INVx1_ASAP7_75t_SL g3519 ( 
.A(n_3276),
.Y(n_3519)
);

OAI22xp5_ASAP7_75t_L g3520 ( 
.A1(n_3360),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3317),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3317),
.Y(n_3522)
);

AOI322xp5_ASAP7_75t_L g3523 ( 
.A1(n_3274),
.A2(n_431),
.A3(n_432),
.B1(n_433),
.B2(n_434),
.C1(n_436),
.C2(n_437),
.Y(n_3523)
);

AOI31xp33_ASAP7_75t_L g3524 ( 
.A1(n_3360),
.A2(n_438),
.A3(n_433),
.B(n_434),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3317),
.Y(n_3525)
);

AOI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3292),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_3526)
);

OAI22xp5_ASAP7_75t_L g3527 ( 
.A1(n_3360),
.A2(n_442),
.B1(n_439),
.B2(n_441),
.Y(n_3527)
);

AOI22xp33_ASAP7_75t_L g3528 ( 
.A1(n_3366),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3317),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_L g3530 ( 
.A(n_3519),
.B(n_443),
.Y(n_3530)
);

AOI221xp5_ASAP7_75t_L g3531 ( 
.A1(n_3428),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.C(n_447),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3419),
.B(n_445),
.Y(n_3532)
);

NOR2xp33_ASAP7_75t_L g3533 ( 
.A(n_3419),
.B(n_447),
.Y(n_3533)
);

OA22x2_ASAP7_75t_L g3534 ( 
.A1(n_3403),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_3534)
);

OAI221xp5_ASAP7_75t_SL g3535 ( 
.A1(n_3410),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.C(n_451),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3386),
.Y(n_3536)
);

NAND3xp33_ASAP7_75t_SL g3537 ( 
.A(n_3504),
.B(n_451),
.C(n_453),
.Y(n_3537)
);

INVx2_ASAP7_75t_SL g3538 ( 
.A(n_3425),
.Y(n_3538)
);

NOR4xp75_ASAP7_75t_L g3539 ( 
.A(n_3384),
.B(n_457),
.C(n_454),
.D(n_455),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3470),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3526),
.B(n_454),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3431),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3526),
.B(n_458),
.Y(n_3543)
);

AOI21xp33_ASAP7_75t_L g3544 ( 
.A1(n_3452),
.A2(n_458),
.B(n_459),
.Y(n_3544)
);

NOR2xp33_ASAP7_75t_L g3545 ( 
.A(n_3524),
.B(n_3510),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3512),
.B(n_459),
.Y(n_3546)
);

OAI322xp33_ASAP7_75t_L g3547 ( 
.A1(n_3469),
.A2(n_460),
.A3(n_461),
.B1(n_462),
.B2(n_463),
.C1(n_464),
.C2(n_465),
.Y(n_3547)
);

AOI211xp5_ASAP7_75t_L g3548 ( 
.A1(n_3377),
.A2(n_467),
.B(n_465),
.C(n_466),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3454),
.B(n_468),
.Y(n_3549)
);

NAND3xp33_ASAP7_75t_L g3550 ( 
.A(n_3441),
.B(n_468),
.C(n_469),
.Y(n_3550)
);

OAI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3382),
.A2(n_470),
.B(n_471),
.Y(n_3551)
);

NAND3xp33_ASAP7_75t_L g3552 ( 
.A(n_3388),
.B(n_470),
.C(n_472),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3427),
.B(n_473),
.Y(n_3553)
);

OAI21xp33_ASAP7_75t_SL g3554 ( 
.A1(n_3378),
.A2(n_473),
.B(n_474),
.Y(n_3554)
);

NOR3xp33_ASAP7_75t_SL g3555 ( 
.A(n_3414),
.B(n_474),
.C(n_475),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3416),
.A2(n_475),
.B(n_476),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_SL g3557 ( 
.A(n_3420),
.B(n_476),
.Y(n_3557)
);

OAI221xp5_ASAP7_75t_SL g3558 ( 
.A1(n_3380),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.C(n_481),
.Y(n_3558)
);

OR2x2_ASAP7_75t_L g3559 ( 
.A(n_3399),
.B(n_478),
.Y(n_3559)
);

HB1xp67_ASAP7_75t_L g3560 ( 
.A(n_3408),
.Y(n_3560)
);

AOI211xp5_ASAP7_75t_L g3561 ( 
.A1(n_3433),
.A2(n_485),
.B(n_481),
.C(n_484),
.Y(n_3561)
);

OAI21xp33_ASAP7_75t_L g3562 ( 
.A1(n_3444),
.A2(n_484),
.B(n_487),
.Y(n_3562)
);

NAND3xp33_ASAP7_75t_SL g3563 ( 
.A(n_3502),
.B(n_487),
.C(n_488),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3516),
.Y(n_3564)
);

INVx1_ASAP7_75t_SL g3565 ( 
.A(n_3508),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3387),
.B(n_488),
.Y(n_3566)
);

AOI221xp5_ASAP7_75t_L g3567 ( 
.A1(n_3383),
.A2(n_491),
.B1(n_489),
.B2(n_490),
.C(n_492),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3409),
.B(n_494),
.Y(n_3568)
);

OAI221xp5_ASAP7_75t_SL g3569 ( 
.A1(n_3503),
.A2(n_497),
.B1(n_494),
.B2(n_496),
.C(n_498),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_SL g3570 ( 
.A(n_3505),
.B(n_497),
.Y(n_3570)
);

AOI211xp5_ASAP7_75t_L g3571 ( 
.A1(n_3496),
.A2(n_501),
.B(n_499),
.C(n_500),
.Y(n_3571)
);

XOR2x2_ASAP7_75t_L g3572 ( 
.A(n_3379),
.B(n_499),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3389),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3507),
.Y(n_3574)
);

AOI211xp5_ASAP7_75t_L g3575 ( 
.A1(n_3498),
.A2(n_503),
.B(n_500),
.C(n_502),
.Y(n_3575)
);

NOR2xp33_ASAP7_75t_SL g3576 ( 
.A(n_3417),
.B(n_503),
.Y(n_3576)
);

AOI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_3453),
.A2(n_504),
.B(n_505),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3406),
.Y(n_3578)
);

NOR3xp33_ASAP7_75t_L g3579 ( 
.A(n_3395),
.B(n_507),
.C(n_508),
.Y(n_3579)
);

OA22x2_ASAP7_75t_L g3580 ( 
.A1(n_3423),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.Y(n_3580)
);

HB1xp67_ASAP7_75t_L g3581 ( 
.A(n_3429),
.Y(n_3581)
);

NOR2x1_ASAP7_75t_L g3582 ( 
.A(n_3392),
.B(n_509),
.Y(n_3582)
);

AND2x2_ASAP7_75t_L g3583 ( 
.A(n_3390),
.B(n_3397),
.Y(n_3583)
);

OR2x2_ASAP7_75t_L g3584 ( 
.A(n_3463),
.B(n_512),
.Y(n_3584)
);

OR2x2_ASAP7_75t_L g3585 ( 
.A(n_3442),
.B(n_512),
.Y(n_3585)
);

NOR3xp33_ASAP7_75t_L g3586 ( 
.A(n_3402),
.B(n_513),
.C(n_515),
.Y(n_3586)
);

NOR2x1_ASAP7_75t_L g3587 ( 
.A(n_3520),
.B(n_513),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3501),
.B(n_515),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3514),
.B(n_516),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3451),
.B(n_517),
.Y(n_3590)
);

OR2x2_ASAP7_75t_L g3591 ( 
.A(n_3430),
.B(n_517),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3412),
.A2(n_518),
.B(n_519),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3418),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3400),
.B(n_518),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3506),
.B(n_520),
.Y(n_3595)
);

INVx2_ASAP7_75t_SL g3596 ( 
.A(n_3439),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3405),
.B(n_522),
.Y(n_3597)
);

OA22x2_ASAP7_75t_L g3598 ( 
.A1(n_3459),
.A2(n_527),
.B1(n_524),
.B2(n_525),
.Y(n_3598)
);

AOI211xp5_ASAP7_75t_L g3599 ( 
.A1(n_3472),
.A2(n_528),
.B(n_525),
.C(n_527),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3474),
.B(n_529),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_3438),
.A2(n_529),
.B(n_530),
.Y(n_3601)
);

NAND3xp33_ASAP7_75t_L g3602 ( 
.A(n_3443),
.B(n_531),
.C(n_533),
.Y(n_3602)
);

NAND3xp33_ASAP7_75t_L g3603 ( 
.A(n_3415),
.B(n_531),
.C(n_533),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3484),
.B(n_535),
.Y(n_3604)
);

NOR2xp33_ASAP7_75t_L g3605 ( 
.A(n_3432),
.B(n_535),
.Y(n_3605)
);

INVxp67_ASAP7_75t_SL g3606 ( 
.A(n_3404),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3411),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3422),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3468),
.B(n_536),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3462),
.B(n_536),
.Y(n_3610)
);

OR2x2_ASAP7_75t_L g3611 ( 
.A(n_3381),
.B(n_538),
.Y(n_3611)
);

AOI21xp33_ASAP7_75t_L g3612 ( 
.A1(n_3458),
.A2(n_538),
.B(n_539),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3424),
.B(n_539),
.Y(n_3613)
);

NOR3x1_ASAP7_75t_L g3614 ( 
.A(n_3437),
.B(n_540),
.C(n_541),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3434),
.B(n_542),
.Y(n_3615)
);

XNOR2xp5_ASAP7_75t_L g3616 ( 
.A(n_3517),
.B(n_542),
.Y(n_3616)
);

OAI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_3455),
.A2(n_543),
.B(n_544),
.Y(n_3617)
);

XNOR2x1_ASAP7_75t_L g3618 ( 
.A(n_3385),
.B(n_543),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3445),
.Y(n_3619)
);

AOI211xp5_ASAP7_75t_L g3620 ( 
.A1(n_3515),
.A2(n_548),
.B(n_544),
.C(n_546),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3560),
.Y(n_3621)
);

NOR2xp67_ASAP7_75t_L g3622 ( 
.A(n_3538),
.B(n_3446),
.Y(n_3622)
);

AOI322xp5_ASAP7_75t_L g3623 ( 
.A1(n_3554),
.A2(n_3426),
.A3(n_3447),
.B1(n_3440),
.B2(n_3449),
.C1(n_3466),
.C2(n_3457),
.Y(n_3623)
);

OR2x2_ASAP7_75t_L g3624 ( 
.A(n_3540),
.B(n_3521),
.Y(n_3624)
);

OAI22xp5_ASAP7_75t_L g3625 ( 
.A1(n_3596),
.A2(n_3528),
.B1(n_3525),
.B2(n_3522),
.Y(n_3625)
);

NAND3xp33_ASAP7_75t_SL g3626 ( 
.A(n_3565),
.B(n_3539),
.C(n_3551),
.Y(n_3626)
);

OAI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3554),
.A2(n_3482),
.B(n_3461),
.Y(n_3627)
);

NAND3xp33_ASAP7_75t_L g3628 ( 
.A(n_3548),
.B(n_3393),
.C(n_3460),
.Y(n_3628)
);

AOI22xp33_ASAP7_75t_L g3629 ( 
.A1(n_3607),
.A2(n_3464),
.B1(n_3485),
.B2(n_3413),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3532),
.B(n_3523),
.Y(n_3630)
);

NOR3x1_ASAP7_75t_L g3631 ( 
.A(n_3617),
.B(n_3529),
.C(n_3435),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3581),
.Y(n_3632)
);

OAI221xp5_ASAP7_75t_L g3633 ( 
.A1(n_3545),
.A2(n_3497),
.B1(n_3511),
.B2(n_3509),
.C(n_3499),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_3573),
.A2(n_3471),
.B1(n_3490),
.B2(n_3493),
.Y(n_3634)
);

AOI211x1_ASAP7_75t_L g3635 ( 
.A1(n_3557),
.A2(n_3473),
.B(n_3487),
.C(n_3480),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3582),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3533),
.B(n_3486),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_3546),
.A2(n_3513),
.B(n_3527),
.Y(n_3638)
);

AOI22xp5_ASAP7_75t_L g3639 ( 
.A1(n_3530),
.A2(n_3483),
.B1(n_3436),
.B2(n_3479),
.Y(n_3639)
);

NOR3xp33_ASAP7_75t_L g3640 ( 
.A(n_3612),
.B(n_3478),
.C(n_3407),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3572),
.Y(n_3641)
);

AOI211xp5_ASAP7_75t_L g3642 ( 
.A1(n_3536),
.A2(n_3489),
.B(n_3467),
.C(n_3518),
.Y(n_3642)
);

AO22x1_ASAP7_75t_L g3643 ( 
.A1(n_3542),
.A2(n_3450),
.B1(n_3456),
.B2(n_3475),
.Y(n_3643)
);

AOI211xp5_ASAP7_75t_L g3644 ( 
.A1(n_3583),
.A2(n_3477),
.B(n_3491),
.C(n_3396),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3618),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3598),
.Y(n_3646)
);

AOI221xp5_ASAP7_75t_SL g3647 ( 
.A1(n_3592),
.A2(n_3476),
.B1(n_3494),
.B2(n_3492),
.C(n_3448),
.Y(n_3647)
);

A2O1A1Ixp33_ASAP7_75t_L g3648 ( 
.A1(n_3577),
.A2(n_3401),
.B(n_3394),
.C(n_3398),
.Y(n_3648)
);

OAI21xp5_ASAP7_75t_L g3649 ( 
.A1(n_3550),
.A2(n_3500),
.B(n_3391),
.Y(n_3649)
);

AOI221x1_ASAP7_75t_L g3650 ( 
.A1(n_3615),
.A2(n_3495),
.B1(n_3488),
.B2(n_3481),
.C(n_3465),
.Y(n_3650)
);

NOR2x1_ASAP7_75t_L g3651 ( 
.A(n_3559),
.B(n_3421),
.Y(n_3651)
);

O2A1O1Ixp33_ASAP7_75t_L g3652 ( 
.A1(n_3558),
.A2(n_551),
.B(n_549),
.C(n_550),
.Y(n_3652)
);

OAI211xp5_ASAP7_75t_SL g3653 ( 
.A1(n_3564),
.A2(n_552),
.B(n_549),
.C(n_550),
.Y(n_3653)
);

OAI221xp5_ASAP7_75t_L g3654 ( 
.A1(n_3549),
.A2(n_553),
.B1(n_555),
.B2(n_556),
.C(n_557),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3534),
.Y(n_3655)
);

AOI21xp33_ASAP7_75t_L g3656 ( 
.A1(n_3606),
.A2(n_556),
.B(n_557),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3555),
.B(n_558),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3590),
.Y(n_3658)
);

OAI31xp33_ASAP7_75t_L g3659 ( 
.A1(n_3552),
.A2(n_562),
.A3(n_559),
.B(n_560),
.Y(n_3659)
);

NAND4xp25_ASAP7_75t_L g3660 ( 
.A(n_3599),
.B(n_562),
.C(n_559),
.D(n_560),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_3537),
.B(n_563),
.Y(n_3661)
);

AOI222xp33_ASAP7_75t_L g3662 ( 
.A1(n_3608),
.A2(n_3619),
.B1(n_3593),
.B2(n_3574),
.C1(n_3578),
.C2(n_3563),
.Y(n_3662)
);

OAI21xp5_ASAP7_75t_SL g3663 ( 
.A1(n_3553),
.A2(n_563),
.B(n_564),
.Y(n_3663)
);

OAI21xp5_ASAP7_75t_L g3664 ( 
.A1(n_3556),
.A2(n_565),
.B(n_566),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3609),
.B(n_568),
.Y(n_3665)
);

NOR2xp33_ASAP7_75t_L g3666 ( 
.A(n_3604),
.B(n_568),
.Y(n_3666)
);

AOI22xp5_ASAP7_75t_L g3667 ( 
.A1(n_3576),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_3667)
);

AOI22xp5_ASAP7_75t_L g3668 ( 
.A1(n_3600),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_3668)
);

AOI322xp5_ASAP7_75t_L g3669 ( 
.A1(n_3587),
.A2(n_573),
.A3(n_575),
.B1(n_576),
.B2(n_577),
.C1(n_578),
.C2(n_579),
.Y(n_3669)
);

OAI21xp5_ASAP7_75t_SL g3670 ( 
.A1(n_3616),
.A2(n_3611),
.B(n_3605),
.Y(n_3670)
);

OAI21xp33_ASAP7_75t_L g3671 ( 
.A1(n_3570),
.A2(n_577),
.B(n_578),
.Y(n_3671)
);

OAI222xp33_ASAP7_75t_L g3672 ( 
.A1(n_3580),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.C1(n_583),
.C2(n_584),
.Y(n_3672)
);

AOI311xp33_ASAP7_75t_L g3673 ( 
.A1(n_3620),
.A2(n_581),
.A3(n_583),
.B(n_584),
.C(n_585),
.Y(n_3673)
);

NAND3xp33_ASAP7_75t_L g3674 ( 
.A(n_3579),
.B(n_585),
.C(n_586),
.Y(n_3674)
);

O2A1O1Ixp33_ASAP7_75t_L g3675 ( 
.A1(n_3613),
.A2(n_588),
.B(n_589),
.C(n_590),
.Y(n_3675)
);

NAND2x1_ASAP7_75t_L g3676 ( 
.A(n_3588),
.B(n_588),
.Y(n_3676)
);

NAND3xp33_ASAP7_75t_L g3677 ( 
.A(n_3586),
.B(n_590),
.C(n_591),
.Y(n_3677)
);

OAI21xp5_ASAP7_75t_L g3678 ( 
.A1(n_3601),
.A2(n_592),
.B(n_593),
.Y(n_3678)
);

NAND3xp33_ASAP7_75t_L g3679 ( 
.A(n_3561),
.B(n_592),
.C(n_593),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3539),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3621),
.Y(n_3681)
);

OAI22x1_ASAP7_75t_L g3682 ( 
.A1(n_3680),
.A2(n_3602),
.B1(n_3603),
.B2(n_3595),
.Y(n_3682)
);

AOI22xp5_ASAP7_75t_L g3683 ( 
.A1(n_3666),
.A2(n_3562),
.B1(n_3568),
.B2(n_3589),
.Y(n_3683)
);

AO22x1_ASAP7_75t_L g3684 ( 
.A1(n_3632),
.A2(n_3614),
.B1(n_3610),
.B2(n_3597),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3636),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3635),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3676),
.Y(n_3687)
);

A2O1A1Ixp33_ASAP7_75t_L g3688 ( 
.A1(n_3661),
.A2(n_3638),
.B(n_3675),
.C(n_3637),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3665),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3657),
.Y(n_3690)
);

CKINVDCx5p33_ASAP7_75t_R g3691 ( 
.A(n_3641),
.Y(n_3691)
);

INVxp67_ASAP7_75t_SL g3692 ( 
.A(n_3622),
.Y(n_3692)
);

AOI22xp5_ASAP7_75t_L g3693 ( 
.A1(n_3630),
.A2(n_3594),
.B1(n_3566),
.B2(n_3541),
.Y(n_3693)
);

AOI221xp5_ASAP7_75t_L g3694 ( 
.A1(n_3633),
.A2(n_3544),
.B1(n_3543),
.B2(n_3531),
.C(n_3591),
.Y(n_3694)
);

INVx2_ASAP7_75t_SL g3695 ( 
.A(n_3624),
.Y(n_3695)
);

OA22x2_ASAP7_75t_L g3696 ( 
.A1(n_3667),
.A2(n_3535),
.B1(n_3575),
.B2(n_3571),
.Y(n_3696)
);

AO22x1_ASAP7_75t_L g3697 ( 
.A1(n_3631),
.A2(n_3569),
.B1(n_3547),
.B2(n_3567),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3646),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3655),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3651),
.Y(n_3700)
);

INVxp67_ASAP7_75t_SL g3701 ( 
.A(n_3652),
.Y(n_3701)
);

AOI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3626),
.A2(n_3585),
.B1(n_3584),
.B2(n_597),
.Y(n_3702)
);

AOI221xp5_ASAP7_75t_L g3703 ( 
.A1(n_3625),
.A2(n_594),
.B1(n_596),
.B2(n_597),
.C(n_598),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3645),
.Y(n_3704)
);

AOI221x1_ASAP7_75t_SL g3705 ( 
.A1(n_3642),
.A2(n_594),
.B1(n_596),
.B2(n_598),
.C(n_599),
.Y(n_3705)
);

OAI31xp33_ASAP7_75t_SL g3706 ( 
.A1(n_3628),
.A2(n_600),
.A3(n_601),
.B(n_602),
.Y(n_3706)
);

O2A1O1Ixp33_ASAP7_75t_SL g3707 ( 
.A1(n_3648),
.A2(n_600),
.B(n_601),
.C(n_603),
.Y(n_3707)
);

OAI22xp5_ASAP7_75t_L g3708 ( 
.A1(n_3639),
.A2(n_604),
.B1(n_605),
.B2(n_606),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3653),
.Y(n_3709)
);

OAI22xp5_ASAP7_75t_L g3710 ( 
.A1(n_3679),
.A2(n_607),
.B1(n_608),
.B2(n_609),
.Y(n_3710)
);

NOR4xp25_ASAP7_75t_L g3711 ( 
.A(n_3670),
.B(n_3629),
.C(n_3627),
.D(n_3634),
.Y(n_3711)
);

AOI22xp5_ASAP7_75t_L g3712 ( 
.A1(n_3668),
.A2(n_607),
.B1(n_608),
.B2(n_609),
.Y(n_3712)
);

OAI22x1_ASAP7_75t_L g3713 ( 
.A1(n_3674),
.A2(n_610),
.B1(n_611),
.B2(n_612),
.Y(n_3713)
);

NAND5xp2_ASAP7_75t_SL g3714 ( 
.A(n_3662),
.B(n_614),
.C(n_615),
.D(n_616),
.E(n_618),
.Y(n_3714)
);

BUFx2_ASAP7_75t_L g3715 ( 
.A(n_3678),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3658),
.Y(n_3716)
);

AOI221x1_ASAP7_75t_L g3717 ( 
.A1(n_3686),
.A2(n_3640),
.B1(n_3671),
.B2(n_3656),
.C(n_3664),
.Y(n_3717)
);

OAI221xp5_ASAP7_75t_L g3718 ( 
.A1(n_3695),
.A2(n_3659),
.B1(n_3644),
.B2(n_3649),
.C(n_3663),
.Y(n_3718)
);

NOR2xp33_ASAP7_75t_R g3719 ( 
.A(n_3681),
.B(n_3623),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3700),
.Y(n_3720)
);

AOI221xp5_ASAP7_75t_L g3721 ( 
.A1(n_3711),
.A2(n_3690),
.B1(n_3684),
.B2(n_3699),
.C(n_3698),
.Y(n_3721)
);

NOR2xp33_ASAP7_75t_L g3722 ( 
.A(n_3687),
.B(n_3672),
.Y(n_3722)
);

AOI211xp5_ASAP7_75t_L g3723 ( 
.A1(n_3685),
.A2(n_3697),
.B(n_3643),
.C(n_3691),
.Y(n_3723)
);

AOI221xp5_ASAP7_75t_L g3724 ( 
.A1(n_3704),
.A2(n_3647),
.B1(n_3677),
.B2(n_3660),
.C(n_3654),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3709),
.Y(n_3725)
);

OAI211xp5_ASAP7_75t_L g3726 ( 
.A1(n_3703),
.A2(n_3669),
.B(n_3673),
.C(n_3650),
.Y(n_3726)
);

AOI221xp5_ASAP7_75t_L g3727 ( 
.A1(n_3701),
.A2(n_3660),
.B1(n_616),
.B2(n_618),
.C(n_619),
.Y(n_3727)
);

AOI22xp33_ASAP7_75t_L g3728 ( 
.A1(n_3689),
.A2(n_614),
.B1(n_619),
.B2(n_620),
.Y(n_3728)
);

AOI22xp5_ASAP7_75t_L g3729 ( 
.A1(n_3683),
.A2(n_3702),
.B1(n_3692),
.B2(n_3693),
.Y(n_3729)
);

NAND5xp2_ASAP7_75t_L g3730 ( 
.A(n_3694),
.B(n_622),
.C(n_623),
.D(n_624),
.E(n_625),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3706),
.B(n_623),
.Y(n_3731)
);

NOR2xp33_ASAP7_75t_R g3732 ( 
.A(n_3714),
.B(n_624),
.Y(n_3732)
);

AOI222xp33_ASAP7_75t_L g3733 ( 
.A1(n_3682),
.A2(n_626),
.B1(n_627),
.B2(n_628),
.C1(n_629),
.C2(n_630),
.Y(n_3733)
);

NAND5xp2_ASAP7_75t_L g3734 ( 
.A(n_3688),
.B(n_628),
.C(n_629),
.D(n_630),
.E(n_631),
.Y(n_3734)
);

INVx2_ASAP7_75t_SL g3735 ( 
.A(n_3715),
.Y(n_3735)
);

NAND3xp33_ASAP7_75t_SL g3736 ( 
.A(n_3723),
.B(n_3721),
.C(n_3719),
.Y(n_3736)
);

AOI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_3722),
.A2(n_3716),
.B1(n_3696),
.B2(n_3710),
.Y(n_3737)
);

AOI221xp5_ASAP7_75t_L g3738 ( 
.A1(n_3720),
.A2(n_3705),
.B1(n_3707),
.B2(n_3713),
.C(n_3708),
.Y(n_3738)
);

AOI211xp5_ASAP7_75t_L g3739 ( 
.A1(n_3726),
.A2(n_3712),
.B(n_632),
.C(n_633),
.Y(n_3739)
);

AOI211xp5_ASAP7_75t_SL g3740 ( 
.A1(n_3718),
.A2(n_3712),
.B(n_632),
.C(n_633),
.Y(n_3740)
);

AOI211xp5_ASAP7_75t_L g3741 ( 
.A1(n_3724),
.A2(n_631),
.B(n_634),
.C(n_635),
.Y(n_3741)
);

OAI221xp5_ASAP7_75t_L g3742 ( 
.A1(n_3735),
.A2(n_636),
.B1(n_637),
.B2(n_639),
.C(n_640),
.Y(n_3742)
);

XNOR2x1_ASAP7_75t_L g3743 ( 
.A(n_3729),
.B(n_640),
.Y(n_3743)
);

NOR2xp33_ASAP7_75t_L g3744 ( 
.A(n_3734),
.B(n_641),
.Y(n_3744)
);

NAND5xp2_ASAP7_75t_L g3745 ( 
.A(n_3727),
.B(n_641),
.C(n_643),
.D(n_644),
.E(n_645),
.Y(n_3745)
);

A2O1A1Ixp33_ASAP7_75t_L g3746 ( 
.A1(n_3731),
.A2(n_644),
.B(n_645),
.C(n_646),
.Y(n_3746)
);

OAI221xp5_ASAP7_75t_SL g3747 ( 
.A1(n_3725),
.A2(n_647),
.B1(n_648),
.B2(n_649),
.C(n_650),
.Y(n_3747)
);

AOI221x1_ASAP7_75t_L g3748 ( 
.A1(n_3730),
.A2(n_651),
.B1(n_652),
.B2(n_653),
.C(n_654),
.Y(n_3748)
);

OAI21xp33_ASAP7_75t_L g3749 ( 
.A1(n_3736),
.A2(n_3732),
.B(n_3733),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3744),
.Y(n_3750)
);

NAND3xp33_ASAP7_75t_L g3751 ( 
.A(n_3739),
.B(n_3717),
.C(n_3728),
.Y(n_3751)
);

AND3x1_ASAP7_75t_L g3752 ( 
.A(n_3741),
.B(n_651),
.C(n_652),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3748),
.B(n_653),
.Y(n_3753)
);

AOI21xp33_ASAP7_75t_L g3754 ( 
.A1(n_3743),
.A2(n_654),
.B(n_655),
.Y(n_3754)
);

OAI22xp5_ASAP7_75t_L g3755 ( 
.A1(n_3737),
.A2(n_656),
.B1(n_657),
.B2(n_658),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3740),
.B(n_656),
.Y(n_3756)
);

NAND3xp33_ASAP7_75t_SL g3757 ( 
.A(n_3738),
.B(n_658),
.C(n_659),
.Y(n_3757)
);

NAND3xp33_ASAP7_75t_L g3758 ( 
.A(n_3746),
.B(n_660),
.C(n_661),
.Y(n_3758)
);

INVxp67_ASAP7_75t_SL g3759 ( 
.A(n_3753),
.Y(n_3759)
);

OAI221xp5_ASAP7_75t_SL g3760 ( 
.A1(n_3749),
.A2(n_3742),
.B1(n_3745),
.B2(n_3747),
.C(n_663),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3752),
.Y(n_3761)
);

OR2x2_ASAP7_75t_L g3762 ( 
.A(n_3756),
.B(n_660),
.Y(n_3762)
);

AOI211xp5_ASAP7_75t_SL g3763 ( 
.A1(n_3760),
.A2(n_3755),
.B(n_3750),
.C(n_3754),
.Y(n_3763)
);

NAND4xp75_ASAP7_75t_L g3764 ( 
.A(n_3761),
.B(n_3757),
.C(n_3751),
.D(n_3758),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3759),
.B(n_661),
.Y(n_3765)
);

XNOR2xp5_ASAP7_75t_L g3766 ( 
.A(n_3764),
.B(n_3762),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3766),
.Y(n_3767)
);

OAI31xp33_ASAP7_75t_L g3768 ( 
.A1(n_3767),
.A2(n_3763),
.A3(n_3765),
.B(n_664),
.Y(n_3768)
);

AOI22xp5_ASAP7_75t_L g3769 ( 
.A1(n_3768),
.A2(n_662),
.B1(n_663),
.B2(n_664),
.Y(n_3769)
);

AOI31xp33_ASAP7_75t_L g3770 ( 
.A1(n_3769),
.A2(n_665),
.A3(n_666),
.B(n_667),
.Y(n_3770)
);

AOI22xp5_ASAP7_75t_L g3771 ( 
.A1(n_3770),
.A2(n_665),
.B1(n_666),
.B2(n_667),
.Y(n_3771)
);

OAI21xp33_ASAP7_75t_SL g3772 ( 
.A1(n_3771),
.A2(n_668),
.B(n_670),
.Y(n_3772)
);

OAI222xp33_ASAP7_75t_L g3773 ( 
.A1(n_3772),
.A2(n_670),
.B1(n_671),
.B2(n_672),
.C1(n_673),
.C2(n_674),
.Y(n_3773)
);

OAI21xp5_ASAP7_75t_L g3774 ( 
.A1(n_3772),
.A2(n_671),
.B(n_672),
.Y(n_3774)
);

INVx2_ASAP7_75t_SL g3775 ( 
.A(n_3774),
.Y(n_3775)
);

HB1xp67_ASAP7_75t_L g3776 ( 
.A(n_3773),
.Y(n_3776)
);

NAND2x2_ASAP7_75t_L g3777 ( 
.A(n_3775),
.B(n_674),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3777),
.A2(n_3776),
.B(n_676),
.Y(n_3778)
);

AOI211xp5_ASAP7_75t_L g3779 ( 
.A1(n_3778),
.A2(n_675),
.B(n_677),
.C(n_679),
.Y(n_3779)
);


endmodule