module fake_netlist_5_2163_n_1524 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1524);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1524;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_1517;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_968;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_783;
wire n_555;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_232),
.B(n_171),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_261),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_109),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_243),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_177),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_203),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_357),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_302),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_221),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_280),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_40),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_312),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_23),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_85),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_142),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_266),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_137),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_170),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_214),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_92),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_150),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_288),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_188),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_218),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_354),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_163),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_262),
.Y(n_415)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_110),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_19),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_148),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_75),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_191),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_146),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_257),
.Y(n_423)
);

BUFx8_ASAP7_75t_SL g424 ( 
.A(n_17),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_366),
.Y(n_425)
);

BUFx5_ASAP7_75t_L g426 ( 
.A(n_161),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_26),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_281),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_166),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_328),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_8),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_98),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_77),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_87),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_387),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_199),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_258),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_363),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_16),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_121),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_240),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_348),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_289),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_47),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_67),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_37),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_117),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_274),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_369),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_160),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_6),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_336),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_186),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_133),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_386),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_310),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_200),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_40),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_337),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_107),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_164),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_119),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_223),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_5),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_335),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_157),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_383),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_96),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_189),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_388),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_81),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_11),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_144),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_0),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_377),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_250),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_307),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_87),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_3),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_64),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_128),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_206),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_265),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_64),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_138),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_318),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_153),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_32),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_2),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_219),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_233),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_174),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_169),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_33),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_356),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_81),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_194),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_381),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_26),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_129),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_239),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_317),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_220),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_254),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_43),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_179),
.B(n_48),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_234),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_105),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_314),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_190),
.B(n_244),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_116),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_216),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_367),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_241),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_210),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_119),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_275),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_320),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_63),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_361),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_117),
.Y(n_523)
);

BUFx5_ASAP7_75t_L g524 ( 
.A(n_222),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_253),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_208),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_152),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_323),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_105),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_141),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_184),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_143),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_134),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_248),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_83),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_202),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_197),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_324),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_79),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_44),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_116),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_151),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_230),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_55),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_83),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_293),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_100),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_334),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_149),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_311),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_126),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_140),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_108),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_209),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_175),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_115),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_38),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_204),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_48),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_47),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_362),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_115),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_24),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_205),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_88),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_2),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_168),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_91),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_380),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_401),
.B(n_0),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_424),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_397),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_397),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_401),
.B(n_1),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_416),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_397),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_397),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_535),
.Y(n_578)
);

OAI21x1_ASAP7_75t_L g579 ( 
.A1(n_393),
.A2(n_131),
.B(n_130),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_392),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_529),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_391),
.Y(n_582)
);

BUFx8_ASAP7_75t_SL g583 ( 
.A(n_446),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_409),
.B(n_4),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_450),
.B(n_5),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_416),
.B(n_6),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_416),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_513),
.B(n_7),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_416),
.Y(n_589)
);

INVx6_ASAP7_75t_L g590 ( 
.A(n_396),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_416),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_493),
.B(n_8),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_427),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_449),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_416),
.B(n_9),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_427),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_399),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_393),
.B(n_10),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_432),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_449),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_463),
.B(n_461),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_463),
.B(n_10),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_464),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_449),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_467),
.Y(n_605)
);

OA21x2_ASAP7_75t_L g606 ( 
.A1(n_395),
.A2(n_11),
.B(n_12),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_536),
.B(n_12),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_426),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_408),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_440),
.Y(n_610)
);

AND2x2_ASAP7_75t_SL g611 ( 
.A(n_452),
.B(n_13),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_467),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_460),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_410),
.B(n_14),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_402),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_392),
.B(n_15),
.Y(n_616)
);

BUFx12f_ASAP7_75t_L g617 ( 
.A(n_529),
.Y(n_617)
);

BUFx12f_ASAP7_75t_L g618 ( 
.A(n_396),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_467),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_478),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_444),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_466),
.Y(n_622)
);

BUFx12f_ASAP7_75t_L g623 ( 
.A(n_420),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_435),
.B(n_16),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_431),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_426),
.Y(n_626)
);

NOR2x1_ASAP7_75t_L g627 ( 
.A(n_389),
.B(n_132),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_478),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_473),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_478),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_545),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_426),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_426),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_434),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_561),
.B(n_18),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_451),
.B(n_20),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_400),
.B(n_20),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_404),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_481),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_426),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_426),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_435),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_548),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_524),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_486),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_562),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_491),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_414),
.B(n_21),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_601),
.B(n_418),
.Y(n_650)
);

NOR2x1p5_ASAP7_75t_L g651 ( 
.A(n_601),
.B(n_433),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_572),
.Y(n_652)
);

AOI21x1_ASAP7_75t_L g653 ( 
.A1(n_587),
.A2(n_406),
.B(n_405),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_572),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_572),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_573),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_573),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_616),
.B(n_423),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_647),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_647),
.Y(n_660)
);

AND2x2_ASAP7_75t_SL g661 ( 
.A(n_611),
.B(n_531),
.Y(n_661)
);

INVxp33_ASAP7_75t_L g662 ( 
.A(n_578),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_596),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_573),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_590),
.B(n_525),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_576),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_590),
.B(n_525),
.Y(n_667)
);

AND3x1_ASAP7_75t_L g668 ( 
.A(n_588),
.B(n_470),
.C(n_462),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_639),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_577),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_577),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_624),
.B(n_468),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_597),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_570),
.B(n_508),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_574),
.B(n_508),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_594),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_594),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_603),
.B(n_417),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_594),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_604),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_588),
.B(n_407),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_590),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_609),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_604),
.Y(n_684)
);

CKINVDCx14_ASAP7_75t_R g685 ( 
.A(n_571),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_604),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_611),
.B(n_429),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_593),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_589),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_625),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_605),
.Y(n_691)
);

BUFx6f_ASAP7_75t_SL g692 ( 
.A(n_614),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_605),
.Y(n_693)
);

BUFx6f_ASAP7_75t_SL g694 ( 
.A(n_614),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_603),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_605),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_591),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_612),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_612),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_689),
.B(n_697),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_658),
.B(n_575),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_655),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_678),
.B(n_635),
.Y(n_703)
);

INVxp33_ASAP7_75t_L g704 ( 
.A(n_662),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_676),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_683),
.B(n_597),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_672),
.B(n_575),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g708 ( 
.A(n_674),
.B(n_598),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_678),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_676),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_650),
.B(n_626),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_665),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_683),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_690),
.B(n_581),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_690),
.B(n_602),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_675),
.B(n_598),
.Y(n_716)
);

AND2x6_ASAP7_75t_L g717 ( 
.A(n_667),
.B(n_584),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_661),
.B(n_602),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_695),
.B(n_637),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_669),
.B(n_639),
.Y(n_720)
);

BUFx6f_ASAP7_75t_SL g721 ( 
.A(n_661),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_652),
.B(n_608),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_699),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_699),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_652),
.B(n_608),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_673),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_654),
.B(n_633),
.Y(n_727)
);

NAND2x1p5_ASAP7_75t_L g728 ( 
.A(n_668),
.B(n_606),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_654),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_691),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_681),
.B(n_636),
.Y(n_731)
);

INVx8_ASAP7_75t_L g732 ( 
.A(n_692),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_669),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_662),
.B(n_637),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_682),
.B(n_636),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_664),
.B(n_633),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_664),
.B(n_634),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_666),
.B(n_634),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_666),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_687),
.B(n_643),
.C(n_580),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_673),
.B(n_585),
.C(n_584),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_655),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_692),
.B(n_618),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_670),
.B(n_671),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_671),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_682),
.B(n_585),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_677),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_679),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_680),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_692),
.B(n_623),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_651),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_680),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_684),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_688),
.B(n_592),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_686),
.B(n_641),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_694),
.B(n_617),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_686),
.B(n_641),
.Y(n_758)
);

OAI22xp33_ASAP7_75t_L g759 ( 
.A1(n_663),
.A2(n_568),
.B1(n_490),
.B2(n_445),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_694),
.A2(n_649),
.B1(n_638),
.B2(n_592),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_685),
.B(n_632),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_693),
.B(n_642),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_693),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_696),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_653),
.B(n_607),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_765),
.A2(n_579),
.B(n_653),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_712),
.B(n_704),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_741),
.A2(n_694),
.B1(n_403),
.B2(n_428),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_729),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_719),
.A2(n_760),
.B1(n_718),
.B2(n_731),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_709),
.B(n_582),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_739),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_740),
.B(n_595),
.C(n_586),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_733),
.B(n_610),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_708),
.B(n_613),
.C(n_599),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_748),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_707),
.B(n_698),
.Y(n_777)
);

INVx11_ASAP7_75t_L g778 ( 
.A(n_717),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_749),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_711),
.B(n_698),
.Y(n_780)
);

NAND2x1p5_ASAP7_75t_L g781 ( 
.A(n_713),
.B(n_512),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_703),
.B(n_582),
.Y(n_782)
);

AO21x1_ASAP7_75t_L g783 ( 
.A1(n_728),
.A2(n_649),
.B(n_638),
.Y(n_783)
);

NOR2xp67_ASAP7_75t_L g784 ( 
.A(n_726),
.B(n_734),
.Y(n_784)
);

NOR2x1_ASAP7_75t_L g785 ( 
.A(n_706),
.B(n_398),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_716),
.A2(n_700),
.B(n_746),
.Y(n_786)
);

AOI21xp33_ASAP7_75t_L g787 ( 
.A1(n_715),
.A2(n_613),
.B(n_552),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_720),
.B(n_621),
.Y(n_788)
);

AO21x1_ASAP7_75t_L g789 ( 
.A1(n_700),
.A2(n_413),
.B(n_411),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_717),
.A2(n_606),
.B(n_627),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_714),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_717),
.A2(n_552),
.B(n_537),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_752),
.A2(n_567),
.B1(n_487),
.B2(n_537),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_721),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_735),
.B(n_599),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_744),
.A2(n_644),
.B(n_600),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_754),
.Y(n_797)
);

OAI21xp33_ASAP7_75t_L g798 ( 
.A1(n_755),
.A2(n_501),
.B(n_498),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_732),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_717),
.A2(n_522),
.B1(n_550),
.B2(n_484),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_722),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_721),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_717),
.B(n_415),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_725),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_751),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_743),
.B(n_622),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_757),
.B(n_469),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_727),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_736),
.A2(n_448),
.B(n_441),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_763),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_730),
.B(n_745),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_759),
.B(n_472),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_737),
.A2(n_756),
.B(n_738),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_747),
.B(n_750),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_753),
.A2(n_503),
.B1(n_511),
.B2(n_497),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_738),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_764),
.B(n_629),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_756),
.A2(n_657),
.B(n_656),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_705),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_702),
.A2(n_645),
.B(n_642),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_SL g821 ( 
.A1(n_758),
.A2(n_762),
.B(n_454),
.C(n_455),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_732),
.B(n_390),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_732),
.B(n_394),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_761),
.B(n_640),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_710),
.B(n_583),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_723),
.B(n_648),
.C(n_646),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_742),
.B(n_457),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_724),
.B(n_447),
.C(n_439),
.Y(n_828)
);

AOI33xp33_ASAP7_75t_L g829 ( 
.A1(n_761),
.A2(n_566),
.A3(n_560),
.B1(n_563),
.B2(n_559),
.B3(n_480),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_761),
.A2(n_620),
.B(n_619),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_732),
.B(n_553),
.Y(n_831)
);

AO21x1_ASAP7_75t_L g832 ( 
.A1(n_728),
.A2(n_471),
.B(n_465),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_740),
.B(n_476),
.C(n_474),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_741),
.A2(n_485),
.B1(n_488),
.B2(n_479),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_765),
.A2(n_630),
.B(n_628),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_708),
.A2(n_492),
.B1(n_495),
.B2(n_494),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_709),
.B(n_615),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_712),
.B(n_583),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_709),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_708),
.A2(n_557),
.B(n_500),
.C(n_502),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_708),
.A2(n_505),
.B(n_506),
.C(n_499),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_708),
.A2(n_514),
.B(n_516),
.C(n_509),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_733),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_709),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_740),
.A2(n_530),
.B1(n_533),
.B2(n_527),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_708),
.A2(n_538),
.B(n_542),
.C(n_534),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_701),
.B(n_543),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_709),
.B(n_615),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_712),
.B(n_659),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_701),
.B(n_546),
.Y(n_850)
);

BUFx8_ASAP7_75t_L g851 ( 
.A(n_721),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_722),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_709),
.B(n_412),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_701),
.B(n_564),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_721),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_712),
.B(n_659),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_733),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_701),
.B(n_569),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_765),
.A2(n_631),
.B(n_532),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_801),
.B(n_419),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_804),
.B(n_421),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_769),
.Y(n_862)
);

OAI22x1_ASAP7_75t_L g863 ( 
.A1(n_775),
.A2(n_660),
.B1(n_496),
.B2(n_507),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_813),
.A2(n_524),
.B(n_135),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_772),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_776),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_766),
.A2(n_425),
.B(n_422),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_773),
.A2(n_436),
.B(n_430),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_786),
.A2(n_438),
.B(n_442),
.C(n_437),
.Y(n_869)
);

OAI21x1_ASAP7_75t_L g870 ( 
.A1(n_790),
.A2(n_524),
.B(n_136),
.Y(n_870)
);

OAI21x1_ASAP7_75t_SL g871 ( 
.A1(n_783),
.A2(n_524),
.B(n_139),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_770),
.A2(n_800),
.B1(n_792),
.B2(n_778),
.Y(n_872)
);

NOR2x1_ASAP7_75t_R g873 ( 
.A(n_799),
.B(n_482),
.Y(n_873)
);

AO31x2_ASAP7_75t_L g874 ( 
.A1(n_832),
.A2(n_28),
.A3(n_25),
.B(n_27),
.Y(n_874)
);

AOI211x1_ASAP7_75t_L g875 ( 
.A1(n_789),
.A2(n_847),
.B(n_854),
.C(n_850),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_818),
.A2(n_147),
.B(n_145),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_808),
.B(n_443),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_843),
.Y(n_878)
);

INVx6_ASAP7_75t_L g879 ( 
.A(n_819),
.Y(n_879)
);

AND2x2_ASAP7_75t_SL g880 ( 
.A(n_849),
.B(n_660),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_814),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_816),
.A2(n_456),
.B(n_453),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_794),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_852),
.B(n_458),
.Y(n_884)
);

AND2x2_ASAP7_75t_SL g885 ( 
.A(n_856),
.B(n_27),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_777),
.A2(n_475),
.B(n_459),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_859),
.A2(n_780),
.B(n_811),
.Y(n_887)
);

CKINVDCx11_ASAP7_75t_R g888 ( 
.A(n_805),
.Y(n_888)
);

OAI22x1_ASAP7_75t_L g889 ( 
.A1(n_767),
.A2(n_518),
.B1(n_521),
.B2(n_510),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_858),
.A2(n_483),
.B(n_477),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_784),
.B(n_489),
.Y(n_891)
);

AOI221x1_ASAP7_75t_L g892 ( 
.A1(n_842),
.A2(n_517),
.B1(n_519),
.B2(n_515),
.C(n_504),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_779),
.Y(n_893)
);

INVx8_ASAP7_75t_L g894 ( 
.A(n_831),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_791),
.B(n_520),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_843),
.B(n_526),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_839),
.Y(n_897)
);

OAI21x1_ASAP7_75t_L g898 ( 
.A1(n_835),
.A2(n_155),
.B(n_154),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_836),
.B(n_549),
.C(n_528),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_809),
.A2(n_555),
.B(n_554),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_797),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_837),
.B(n_558),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_844),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_848),
.B(n_523),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_843),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_845),
.A2(n_540),
.B1(n_541),
.B2(n_539),
.Y(n_906)
);

OAI21x1_ASAP7_75t_L g907 ( 
.A1(n_779),
.A2(n_810),
.B(n_827),
.Y(n_907)
);

O2A1O1Ixp5_ASAP7_75t_L g908 ( 
.A1(n_846),
.A2(n_547),
.B(n_551),
.C(n_544),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_857),
.B(n_156),
.Y(n_909)
);

AOI21xp33_ASAP7_75t_L g910 ( 
.A1(n_785),
.A2(n_565),
.B(n_556),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_781),
.A2(n_159),
.B1(n_162),
.B2(n_158),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_787),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_788),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_788),
.Y(n_914)
);

AOI221xp5_ASAP7_75t_L g915 ( 
.A1(n_793),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.C(n_33),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_821),
.A2(n_167),
.B(n_165),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_795),
.B(n_31),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_841),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_840),
.A2(n_173),
.B(n_172),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_782),
.B(n_34),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_774),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_853),
.A2(n_178),
.B(n_176),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_857),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_857),
.B(n_180),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_796),
.A2(n_182),
.B(n_181),
.Y(n_925)
);

OAI21x1_ASAP7_75t_SL g926 ( 
.A1(n_830),
.A2(n_185),
.B(n_183),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_774),
.B(n_187),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_833),
.A2(n_193),
.B(n_192),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_822),
.A2(n_196),
.B(n_195),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_806),
.B(n_35),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_823),
.A2(n_201),
.B(n_198),
.Y(n_931)
);

AOI221x1_ASAP7_75t_L g932 ( 
.A1(n_834),
.A2(n_251),
.B1(n_385),
.B2(n_384),
.C(n_382),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_829),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_771),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_824),
.B(n_36),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_819),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_831),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_798),
.B(n_812),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_768),
.A2(n_211),
.B(n_207),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_798),
.A2(n_213),
.B(n_212),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_807),
.A2(n_217),
.B(n_215),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_828),
.A2(n_826),
.B(n_831),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_802),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_815),
.A2(n_225),
.B(n_224),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_SL g945 ( 
.A(n_838),
.B(n_37),
.C(n_38),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_SL g946 ( 
.A(n_855),
.B(n_39),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_825),
.A2(n_227),
.B1(n_228),
.B2(n_226),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_851),
.B(n_39),
.Y(n_948)
);

OAI21x1_ASAP7_75t_L g949 ( 
.A1(n_851),
.A2(n_231),
.B(n_229),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_790),
.A2(n_236),
.B(n_235),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_770),
.B(n_237),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_790),
.A2(n_242),
.B(n_238),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_773),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_953)
);

AOI221xp5_ASAP7_75t_L g954 ( 
.A1(n_787),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.C(n_45),
.Y(n_954)
);

OAI21x1_ASAP7_75t_SL g955 ( 
.A1(n_783),
.A2(n_246),
.B(n_245),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_779),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_839),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_801),
.B(n_45),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_801),
.B(n_46),
.Y(n_959)
);

NOR2x1_ASAP7_75t_SL g960 ( 
.A(n_803),
.B(n_247),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_817),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_801),
.B(n_46),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_801),
.B(n_49),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_773),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_790),
.A2(n_252),
.B(n_249),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_769),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_767),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_767),
.B(n_50),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_790),
.A2(n_256),
.B(n_255),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_801),
.B(n_51),
.Y(n_970)
);

O2A1O1Ixp5_ASAP7_75t_L g971 ( 
.A1(n_832),
.A2(n_285),
.B(n_376),
.C(n_375),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_820),
.A2(n_378),
.B(n_260),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_801),
.B(n_52),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_767),
.B(n_52),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_801),
.B(n_53),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_843),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_813),
.A2(n_263),
.B(n_259),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_801),
.B(n_53),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_817),
.Y(n_979)
);

CKINVDCx8_ASAP7_75t_R g980 ( 
.A(n_794),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_769),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_790),
.A2(n_267),
.B(n_264),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_839),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_820),
.A2(n_374),
.B(n_269),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_820),
.A2(n_373),
.B(n_270),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_817),
.Y(n_986)
);

AO21x1_ASAP7_75t_L g987 ( 
.A1(n_792),
.A2(n_54),
.B(n_55),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_773),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_988)
);

AOI221xp5_ASAP7_75t_L g989 ( 
.A1(n_787),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.C(n_59),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_801),
.B(n_58),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_813),
.A2(n_271),
.B(n_268),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_801),
.B(n_59),
.Y(n_992)
);

OAI22x1_ASAP7_75t_L g993 ( 
.A1(n_775),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_790),
.A2(n_273),
.B(n_272),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_813),
.A2(n_277),
.B(n_276),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_801),
.B(n_60),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_771),
.B(n_61),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_SL g998 ( 
.A(n_792),
.B(n_63),
.Y(n_998)
);

NOR2xp67_ASAP7_75t_L g999 ( 
.A(n_786),
.B(n_278),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_773),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_801),
.B(n_65),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_801),
.B(n_66),
.Y(n_1002)
);

INVxp67_ASAP7_75t_SL g1003 ( 
.A(n_843),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_769),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_769),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_907),
.A2(n_282),
.B(n_279),
.Y(n_1006)
);

OA21x2_ASAP7_75t_L g1007 ( 
.A1(n_870),
.A2(n_284),
.B(n_283),
.Y(n_1007)
);

NOR2xp67_ASAP7_75t_L g1008 ( 
.A(n_881),
.B(n_372),
.Y(n_1008)
);

NAND2x1_ASAP7_75t_L g1009 ( 
.A(n_878),
.B(n_905),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_967),
.B(n_68),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_862),
.Y(n_1011)
);

AO21x2_ASAP7_75t_L g1012 ( 
.A1(n_867),
.A2(n_287),
.B(n_286),
.Y(n_1012)
);

AO21x2_ASAP7_75t_L g1013 ( 
.A1(n_867),
.A2(n_291),
.B(n_290),
.Y(n_1013)
);

AO21x2_ASAP7_75t_L g1014 ( 
.A1(n_951),
.A2(n_999),
.B(n_991),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_894),
.B(n_292),
.Y(n_1015)
);

AO21x2_ASAP7_75t_L g1016 ( 
.A1(n_999),
.A2(n_295),
.B(n_294),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_865),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_897),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_864),
.A2(n_305),
.B(n_370),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_888),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_866),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_901),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_872),
.A2(n_371),
.B(n_304),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_903),
.Y(n_1024)
);

INVx6_ASAP7_75t_L g1025 ( 
.A(n_879),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_998),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_883),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_875),
.B(n_296),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_957),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_966),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_981),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_943),
.Y(n_1032)
);

AO21x2_ASAP7_75t_L g1033 ( 
.A1(n_977),
.A2(n_306),
.B(n_364),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_950),
.A2(n_365),
.B(n_303),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1004),
.Y(n_1035)
);

AO21x2_ASAP7_75t_L g1036 ( 
.A1(n_995),
.A2(n_919),
.B(n_871),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_998),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_1037)
);

AO21x1_ASAP7_75t_L g1038 ( 
.A1(n_952),
.A2(n_71),
.B(n_72),
.Y(n_1038)
);

BUFx12f_ASAP7_75t_L g1039 ( 
.A(n_879),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_983),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_913),
.B(n_297),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_887),
.A2(n_308),
.B(n_359),
.Y(n_1042)
);

OR2x6_ASAP7_75t_L g1043 ( 
.A(n_894),
.B(n_298),
.Y(n_1043)
);

INVx5_ASAP7_75t_L g1044 ( 
.A(n_878),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_980),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_878),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_965),
.A2(n_301),
.B(n_358),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1005),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_938),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_934),
.B(n_73),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_936),
.Y(n_1051)
);

AO222x2_ASAP7_75t_L g1052 ( 
.A1(n_997),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.C1(n_77),
.C2(n_78),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_972),
.A2(n_313),
.B(n_355),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_921),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_984),
.A2(n_309),
.B(n_353),
.Y(n_1055)
);

NOR2x1_ASAP7_75t_R g1056 ( 
.A(n_937),
.B(n_76),
.Y(n_1056)
);

AO21x2_ASAP7_75t_L g1057 ( 
.A1(n_869),
.A2(n_315),
.B(n_352),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_914),
.B(n_299),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_905),
.Y(n_1059)
);

NOR2xp67_ASAP7_75t_L g1060 ( 
.A(n_860),
.B(n_360),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_893),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_880),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_905),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_969),
.A2(n_300),
.B(n_350),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_976),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_1003),
.B(n_316),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_893),
.Y(n_1067)
);

CKINVDCx11_ASAP7_75t_R g1068 ( 
.A(n_894),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_976),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_976),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_982),
.A2(n_351),
.B(n_349),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_861),
.B(n_347),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_985),
.A2(n_346),
.B(n_345),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_917),
.B(n_78),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_SL g1075 ( 
.A1(n_955),
.A2(n_344),
.B(n_343),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_956),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_882),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_1077)
);

AO21x2_ASAP7_75t_L g1078 ( 
.A1(n_882),
.A2(n_994),
.B(n_928),
.Y(n_1078)
);

OAI321xp33_ASAP7_75t_L g1079 ( 
.A1(n_954),
.A2(n_80),
.A3(n_82),
.B1(n_84),
.B2(n_85),
.C(n_86),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_877),
.B(n_84),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_956),
.Y(n_1081)
);

OAI22xp33_ASAP7_75t_SL g1082 ( 
.A1(n_968),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_935),
.Y(n_1083)
);

AO21x2_ASAP7_75t_L g1084 ( 
.A1(n_928),
.A2(n_342),
.B(n_341),
.Y(n_1084)
);

INVx6_ASAP7_75t_L g1085 ( 
.A(n_937),
.Y(n_1085)
);

OA21x2_ASAP7_75t_L g1086 ( 
.A1(n_876),
.A2(n_340),
.B(n_339),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_895),
.B(n_89),
.Y(n_1087)
);

AO21x2_ASAP7_75t_L g1088 ( 
.A1(n_890),
.A2(n_338),
.B(n_333),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_923),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_885),
.B(n_90),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_961),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_974),
.Y(n_1092)
);

BUFx2_ASAP7_75t_SL g1093 ( 
.A(n_923),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_L g1094 ( 
.A(n_890),
.B(n_90),
.C(n_91),
.Y(n_1094)
);

AO21x2_ASAP7_75t_L g1095 ( 
.A1(n_900),
.A2(n_332),
.B(n_331),
.Y(n_1095)
);

INVxp67_ASAP7_75t_L g1096 ( 
.A(n_920),
.Y(n_1096)
);

OA21x2_ASAP7_75t_L g1097 ( 
.A1(n_940),
.A2(n_330),
.B(n_329),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_979),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_941),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_927),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_884),
.B(n_92),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_986),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_932),
.A2(n_327),
.B(n_325),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_927),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_958),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_863),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_898),
.A2(n_322),
.B(n_321),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_959),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_900),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_1109)
);

NAND2x1p5_ASAP7_75t_L g1110 ( 
.A(n_896),
.B(n_319),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_962),
.Y(n_1111)
);

BUFx5_ASAP7_75t_L g1112 ( 
.A(n_933),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_930),
.B(n_963),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_970),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_868),
.A2(n_127),
.B(n_94),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_973),
.Y(n_1116)
);

NAND3xp33_ASAP7_75t_L g1117 ( 
.A(n_989),
.B(n_93),
.C(n_95),
.Y(n_1117)
);

AO21x2_ASAP7_75t_L g1118 ( 
.A1(n_868),
.A2(n_916),
.B(n_944),
.Y(n_1118)
);

OA21x2_ASAP7_75t_L g1119 ( 
.A1(n_892),
.A2(n_96),
.B(n_97),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_975),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_971),
.A2(n_99),
.B(n_101),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_889),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1002),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_948),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_949),
.Y(n_1125)
);

BUFx4f_ASAP7_75t_SL g1126 ( 
.A(n_891),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_978),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_875),
.B(n_102),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_910),
.A2(n_103),
.B(n_104),
.C(n_106),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_SL g1130 ( 
.A1(n_926),
.A2(n_106),
.B(n_107),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_909),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_902),
.A2(n_108),
.B(n_109),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_908),
.A2(n_110),
.B(n_111),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_990),
.Y(n_1134)
);

AO21x2_ASAP7_75t_L g1135 ( 
.A1(n_992),
.A2(n_127),
.B(n_112),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_996),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_904),
.B(n_111),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_R g1138 ( 
.A(n_947),
.B(n_113),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_924),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1001),
.A2(n_113),
.B(n_114),
.Y(n_1140)
);

BUFx12f_ASAP7_75t_L g1141 ( 
.A(n_873),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_873),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_942),
.B(n_114),
.Y(n_1143)
);

CKINVDCx6p67_ASAP7_75t_R g1144 ( 
.A(n_993),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_939),
.A2(n_118),
.B(n_120),
.C(n_121),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_SL g1146 ( 
.A1(n_987),
.A2(n_960),
.B(n_931),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_906),
.B(n_118),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_953),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_906),
.B(n_122),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_918),
.A2(n_123),
.B(n_124),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_988),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_922),
.A2(n_929),
.B(n_925),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_946),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1000),
.A2(n_915),
.B1(n_947),
.B2(n_945),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_911),
.B(n_964),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_912),
.A2(n_899),
.B(n_886),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_874),
.B(n_946),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1113),
.B(n_874),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1054),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1017),
.Y(n_1160)
);

CKINVDCx6p67_ASAP7_75t_R g1161 ( 
.A(n_1039),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1011),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1021),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1022),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1031),
.Y(n_1165)
);

AOI221xp5_ASAP7_75t_L g1166 ( 
.A1(n_1147),
.A2(n_1149),
.B1(n_1079),
.B2(n_1117),
.C(n_1151),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1024),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1111),
.B(n_1114),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1030),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1035),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1083),
.B(n_1090),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1083),
.B(n_1092),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1100),
.B(n_1104),
.Y(n_1173)
);

OAI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_1154),
.A2(n_1140),
.B1(n_1109),
.B2(n_1077),
.C(n_1026),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1032),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1048),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1154),
.A2(n_1074),
.B1(n_1151),
.B2(n_1094),
.Y(n_1177)
);

CKINVDCx11_ASAP7_75t_R g1178 ( 
.A(n_1045),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_1018),
.Y(n_1179)
);

AO21x1_ASAP7_75t_L g1180 ( 
.A1(n_1023),
.A2(n_1047),
.B(n_1034),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1091),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1040),
.Y(n_1182)
);

OAI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1117),
.A2(n_1010),
.B(n_1137),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1098),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1094),
.A2(n_1140),
.B1(n_1150),
.B2(n_1148),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1102),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1076),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1067),
.Y(n_1188)
);

AO21x1_ASAP7_75t_L g1189 ( 
.A1(n_1023),
.A2(n_1047),
.B(n_1034),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1150),
.A2(n_1143),
.B1(n_1115),
.B2(n_1082),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1064),
.A2(n_1071),
.B(n_1133),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1050),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1028),
.A2(n_1071),
.B(n_1064),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1116),
.B(n_1127),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1105),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1108),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1143),
.A2(n_1115),
.B1(n_1082),
.B2(n_1087),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1123),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1134),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1061),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1136),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1052),
.A2(n_1153),
.B1(n_1062),
.B2(n_1079),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1061),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1152),
.A2(n_1042),
.B(n_1006),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1143),
.A2(n_1155),
.B1(n_1078),
.B2(n_1038),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1081),
.Y(n_1206)
);

INVxp67_ASAP7_75t_SL g1207 ( 
.A(n_1112),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1081),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1112),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1112),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1029),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1041),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1120),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1018),
.Y(n_1214)
);

AO21x2_ASAP7_75t_L g1215 ( 
.A1(n_1078),
.A2(n_1118),
.B(n_1036),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1027),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1044),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1058),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1120),
.Y(n_1219)
);

BUFx4f_ASAP7_75t_L g1220 ( 
.A(n_1025),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1044),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1104),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1096),
.B(n_1124),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1153),
.B(n_1144),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1058),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_1044),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1104),
.Y(n_1227)
);

AO21x2_ASAP7_75t_L g1228 ( 
.A1(n_1118),
.A2(n_1036),
.B(n_1014),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1093),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1157),
.A2(n_1103),
.B1(n_1084),
.B2(n_1138),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1100),
.B(n_1106),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1066),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1155),
.A2(n_1156),
.B(n_1060),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1103),
.A2(n_1155),
.B1(n_1157),
.B2(n_1037),
.Y(n_1234)
);

INVx4_ASAP7_75t_SL g1235 ( 
.A(n_1015),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1089),
.B(n_1131),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1025),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1066),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1128),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1084),
.A2(n_1132),
.B1(n_1119),
.B2(n_1128),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1063),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1065),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1046),
.Y(n_1243)
);

BUFx12f_ASAP7_75t_L g1244 ( 
.A(n_1068),
.Y(n_1244)
);

OAI221xp5_ASAP7_75t_L g1245 ( 
.A1(n_1129),
.A2(n_1049),
.B1(n_1145),
.B2(n_1101),
.C(n_1080),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1069),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1135),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1135),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1059),
.B(n_1122),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1065),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1009),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1051),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1070),
.B(n_1139),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1028),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1046),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1008),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1065),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1085),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1099),
.A2(n_1055),
.B(n_1053),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1085),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1008),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1015),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1126),
.A2(n_1043),
.B1(n_1015),
.B2(n_1060),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1043),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1014),
.A2(n_1156),
.B(n_1033),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1072),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1072),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1119),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1043),
.A2(n_1095),
.B1(n_1033),
.B2(n_1013),
.Y(n_1269)
);

AOI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1007),
.A2(n_1019),
.B(n_1073),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1110),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1095),
.A2(n_1012),
.B1(n_1013),
.B2(n_1088),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1130),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1007),
.A2(n_1019),
.B(n_1073),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1121),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1121),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1107),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1125),
.B(n_1142),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1141),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1012),
.B(n_1088),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1020),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1097),
.A2(n_1086),
.B1(n_1056),
.B2(n_1075),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1016),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1016),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1057),
.B(n_1086),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1056),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1078),
.A2(n_1146),
.B(n_1118),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1171),
.B(n_1172),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1180),
.A2(n_1189),
.A3(n_1280),
.B(n_1275),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1213),
.B(n_1219),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1224),
.B(n_1214),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1214),
.B(n_1192),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1179),
.B(n_1168),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1202),
.A2(n_1166),
.B1(n_1183),
.B2(n_1174),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1276),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1159),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1179),
.B(n_1194),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1182),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1202),
.A2(n_1185),
.B1(n_1177),
.B2(n_1166),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1167),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1223),
.B(n_1249),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1220),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1199),
.B(n_1201),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1183),
.A2(n_1174),
.B1(n_1177),
.B2(n_1185),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1195),
.B(n_1196),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1175),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1190),
.A2(n_1197),
.B1(n_1245),
.B2(n_1193),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1190),
.A2(n_1197),
.B1(n_1245),
.B2(n_1193),
.Y(n_1308)
);

AND2x4_ASAP7_75t_SL g1309 ( 
.A(n_1161),
.B(n_1236),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1181),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1184),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1232),
.B(n_1238),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1160),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1205),
.A2(n_1225),
.B1(n_1218),
.B2(n_1263),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1198),
.B(n_1162),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1235),
.B(n_1212),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1164),
.B(n_1165),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1241),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1163),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1209),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1176),
.B(n_1186),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1231),
.B(n_1246),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1211),
.B(n_1262),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1169),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1216),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1211),
.B(n_1170),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1226),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1264),
.B(n_1235),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1226),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1188),
.B(n_1222),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1234),
.A2(n_1286),
.B1(n_1207),
.B2(n_1191),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1263),
.A2(n_1278),
.B1(n_1271),
.B2(n_1267),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1236),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1253),
.B(n_1227),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1278),
.B(n_1173),
.Y(n_1335)
);

AO31x2_ASAP7_75t_L g1336 ( 
.A1(n_1280),
.A2(n_1284),
.A3(n_1283),
.B(n_1234),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1239),
.B(n_1254),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1220),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1173),
.B(n_1252),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1187),
.B(n_1229),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1200),
.B(n_1286),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1200),
.B(n_1286),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1203),
.B(n_1208),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1158),
.B(n_1206),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1260),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1251),
.B(n_1266),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1210),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1217),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1268),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1247),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1258),
.B(n_1158),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1258),
.B(n_1243),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1255),
.B(n_1221),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1205),
.B(n_1256),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1260),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1237),
.B(n_1281),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1217),
.B(n_1250),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1221),
.B(n_1242),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1242),
.B(n_1250),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1257),
.B(n_1178),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1248),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1260),
.B(n_1273),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1261),
.B(n_1240),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1244),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1240),
.B(n_1230),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1230),
.A2(n_1191),
.B1(n_1265),
.B2(n_1269),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1233),
.B(n_1269),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1279),
.B(n_1265),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1287),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1287),
.B(n_1215),
.Y(n_1370)
);

BUFx8_ASAP7_75t_L g1371 ( 
.A(n_1277),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1228),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1282),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1259),
.B(n_1285),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1349),
.B(n_1215),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1293),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1297),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1349),
.B(n_1228),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1368),
.B(n_1272),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1350),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1299),
.A2(n_1204),
.B1(n_1270),
.B2(n_1274),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1361),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1292),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1288),
.B(n_1294),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1307),
.B(n_1308),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1351),
.B(n_1290),
.Y(n_1386)
);

AOI211xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1314),
.A2(n_1354),
.B(n_1332),
.C(n_1365),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1307),
.B(n_1308),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1295),
.B(n_1344),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1294),
.A2(n_1304),
.B1(n_1367),
.B2(n_1371),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1291),
.B(n_1301),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1304),
.B(n_1315),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1326),
.B(n_1311),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1296),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1289),
.B(n_1373),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1340),
.B(n_1300),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1298),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1310),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1334),
.B(n_1324),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1305),
.B(n_1321),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1303),
.B(n_1317),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1313),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1338),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1347),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1323),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1312),
.B(n_1337),
.Y(n_1406)
);

NOR2xp67_ASAP7_75t_L g1407 ( 
.A(n_1345),
.B(n_1355),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1289),
.B(n_1363),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1289),
.B(n_1336),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1319),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1312),
.B(n_1330),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1289),
.B(n_1331),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1331),
.B(n_1347),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1371),
.A2(n_1328),
.B1(n_1316),
.B2(n_1362),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1322),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1370),
.B(n_1343),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1312),
.B(n_1318),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1357),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1333),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1352),
.B(n_1353),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1318),
.A2(n_1302),
.B1(n_1348),
.B2(n_1306),
.Y(n_1421)
);

NOR3xp33_ASAP7_75t_L g1422 ( 
.A(n_1345),
.B(n_1355),
.C(n_1360),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1348),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1376),
.B(n_1358),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1380),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1389),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1377),
.B(n_1359),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1382),
.Y(n_1428)
);

NAND4xp25_ASAP7_75t_L g1429 ( 
.A(n_1387),
.B(n_1341),
.C(n_1342),
.D(n_1366),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1383),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1403),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1416),
.B(n_1336),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1413),
.B(n_1374),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1413),
.B(n_1374),
.Y(n_1434)
);

INVxp67_ASAP7_75t_SL g1435 ( 
.A(n_1423),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1404),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1394),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1416),
.B(n_1336),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1386),
.B(n_1320),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1379),
.B(n_1408),
.Y(n_1440)
);

NOR2xp67_ASAP7_75t_L g1441 ( 
.A(n_1407),
.B(n_1339),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1379),
.B(n_1336),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1408),
.B(n_1372),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1412),
.B(n_1372),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1418),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1412),
.B(n_1375),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1395),
.B(n_1369),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1445),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1431),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1431),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1435),
.B(n_1420),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1436),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1430),
.B(n_1420),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1424),
.B(n_1405),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1427),
.B(n_1406),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1425),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1425),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1439),
.B(n_1396),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1443),
.B(n_1446),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1443),
.B(n_1409),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1428),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1440),
.B(n_1432),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1440),
.B(n_1378),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1438),
.B(n_1366),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1438),
.B(n_1395),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1426),
.B(n_1399),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1426),
.B(n_1393),
.Y(n_1467)
);

BUFx2_ASAP7_75t_SL g1468 ( 
.A(n_1441),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1456),
.Y(n_1469)
);

OAI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1448),
.A2(n_1390),
.B1(n_1429),
.B2(n_1422),
.C(n_1384),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1457),
.Y(n_1471)
);

OAI32xp33_ASAP7_75t_L g1472 ( 
.A1(n_1460),
.A2(n_1415),
.A3(n_1447),
.B1(n_1385),
.B2(n_1388),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1461),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1453),
.Y(n_1474)
);

OAI321xp33_ASAP7_75t_L g1475 ( 
.A1(n_1451),
.A2(n_1385),
.A3(n_1388),
.B1(n_1381),
.B2(n_1421),
.C(n_1392),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1452),
.Y(n_1476)
);

NAND2x1_ASAP7_75t_SL g1477 ( 
.A(n_1464),
.B(n_1442),
.Y(n_1477)
);

OAI21xp33_ASAP7_75t_L g1478 ( 
.A1(n_1464),
.A2(n_1442),
.B(n_1381),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1466),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1449),
.B(n_1433),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1465),
.B(n_1444),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1459),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1463),
.B(n_1434),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1449),
.B(n_1431),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1475),
.A2(n_1433),
.B1(n_1462),
.B2(n_1459),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1474),
.B(n_1467),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1469),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1471),
.Y(n_1488)
);

OAI321xp33_ASAP7_75t_L g1489 ( 
.A1(n_1478),
.A2(n_1470),
.A3(n_1433),
.B1(n_1484),
.B2(n_1479),
.C(n_1473),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1470),
.A2(n_1468),
.B1(n_1434),
.B2(n_1433),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1475),
.A2(n_1454),
.B1(n_1458),
.B2(n_1397),
.C(n_1455),
.Y(n_1491)
);

XOR2x2_ASAP7_75t_L g1492 ( 
.A(n_1477),
.B(n_1356),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1487),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1490),
.A2(n_1481),
.B1(n_1482),
.B2(n_1462),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1488),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1489),
.A2(n_1472),
.B(n_1484),
.C(n_1403),
.Y(n_1496)
);

OAI22x1_ASAP7_75t_L g1497 ( 
.A1(n_1486),
.A2(n_1480),
.B1(n_1450),
.B2(n_1483),
.Y(n_1497)
);

NAND5xp2_ASAP7_75t_L g1498 ( 
.A(n_1496),
.B(n_1491),
.C(n_1414),
.D(n_1485),
.E(n_1335),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1493),
.B(n_1492),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1495),
.Y(n_1500)
);

NOR4xp25_ASAP7_75t_L g1501 ( 
.A(n_1494),
.B(n_1391),
.C(n_1410),
.D(n_1402),
.Y(n_1501)
);

NAND4xp25_ASAP7_75t_L g1502 ( 
.A(n_1497),
.B(n_1419),
.C(n_1417),
.D(n_1400),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1496),
.A2(n_1364),
.B(n_1309),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1501),
.B(n_1481),
.Y(n_1504)
);

NAND5xp2_ASAP7_75t_L g1505 ( 
.A(n_1503),
.B(n_1401),
.C(n_1398),
.D(n_1411),
.E(n_1444),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1500),
.B(n_1371),
.C(n_1437),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1504),
.B(n_1499),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1506),
.Y(n_1508)
);

NAND4xp75_ASAP7_75t_L g1509 ( 
.A(n_1508),
.B(n_1498),
.C(n_1325),
.D(n_1450),
.Y(n_1509)
);

NAND4xp75_ASAP7_75t_L g1510 ( 
.A(n_1509),
.B(n_1507),
.C(n_1325),
.D(n_1364),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1510),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1510),
.B(n_1364),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1511),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1512),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1513),
.A2(n_1512),
.B(n_1502),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1514),
.A2(n_1302),
.B(n_1505),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1515),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1516),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1517),
.A2(n_1364),
.B(n_1309),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1518),
.A2(n_1346),
.B(n_1327),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1519),
.A2(n_1346),
.B(n_1480),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1520),
.B(n_1346),
.Y(n_1522)
);

AO21x2_ASAP7_75t_L g1523 ( 
.A1(n_1521),
.A2(n_1316),
.B(n_1476),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1523),
.A2(n_1522),
.B1(n_1329),
.B2(n_1327),
.Y(n_1524)
);


endmodule