module fake_jpeg_18206_n_120 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_1),
.Y(n_65)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_72),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_47),
.B1(n_54),
.B2(n_33),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_70),
.B1(n_55),
.B2(n_38),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_51),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_49),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_57),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_73),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_87),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_46),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_82),
.B1(n_80),
.B2(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_52),
.B1(n_50),
.B2(n_45),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_97),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_3),
.C(n_4),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_4),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_43),
.B1(n_35),
.B2(n_7),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_3),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_15),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_105),
.Y(n_109)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_97),
.B1(n_88),
.B2(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_110),
.Y(n_111)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_104),
.B(n_96),
.CON(n_110),
.SN(n_110)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_104),
.B(n_109),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_110),
.B1(n_101),
.B2(n_100),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_107),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_114),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_103),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_91),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_9),
.B(n_10),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_11),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_12),
.Y(n_120)
);


endmodule