module fake_ibex_1682_n_904 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_904);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_904;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_506;
wire n_564;
wire n_562;
wire n_444;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_298;
wire n_202;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_109),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_60),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_47),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_104),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_50),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_49),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_58),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_5),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_92),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_160),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_70),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_9),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_51),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_22),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_31),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_94),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_45),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_64),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_28),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_76),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_63),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_19),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_73),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_125),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_158),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_L g219 ( 
.A(n_102),
.B(n_142),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_96),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_78),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_122),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_108),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_57),
.B(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_117),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_132),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_72),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_59),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_105),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_56),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_68),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_170),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_166),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_55),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_148),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_28),
.B(n_129),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_19),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_114),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_69),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_L g244 ( 
.A(n_27),
.B(n_79),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_27),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_146),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_173),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_52),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_3),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_29),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_34),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_9),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_112),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_87),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_131),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_2),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_167),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_89),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_20),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_81),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_44),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_39),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_141),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_86),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_20),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_46),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_165),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_175),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_140),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_130),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g273 ( 
.A(n_121),
.B(n_25),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_95),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_82),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_161),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_37),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_143),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_22),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_11),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_11),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_75),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_48),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_31),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_145),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_29),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_162),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_119),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_38),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_99),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_90),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_150),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_197),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_252),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_0),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_197),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_199),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_179),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_197),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_179),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_228),
.B(n_1),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_182),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_245),
.B(n_4),
.Y(n_306)
);

OA21x2_ASAP7_75t_L g307 ( 
.A1(n_182),
.A2(n_98),
.B(n_174),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

OA21x2_ASAP7_75t_L g310 ( 
.A1(n_203),
.A2(n_97),
.B(n_171),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_203),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_229),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_4),
.Y(n_314)
);

CKINVDCx6p67_ASAP7_75t_R g315 ( 
.A(n_272),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_229),
.B(n_6),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_211),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_237),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_211),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_287),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_242),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_242),
.B(n_40),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_255),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_177),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_193),
.B(n_6),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_188),
.B(n_7),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_198),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_214),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_255),
.B(n_7),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_180),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_181),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_183),
.B(n_8),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_186),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_187),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_189),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_191),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_194),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_195),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_277),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_200),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_201),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_205),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_206),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_207),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_209),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_240),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_251),
.Y(n_350)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_193),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_277),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_266),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_210),
.B(n_8),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_193),
.B(n_10),
.Y(n_355)
);

OAI22x1_ASAP7_75t_SL g356 ( 
.A1(n_196),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_212),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_284),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_358)
);

BUFx8_ASAP7_75t_L g359 ( 
.A(n_225),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_215),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_216),
.Y(n_361)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_178),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_220),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_286),
.B(n_15),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_222),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_223),
.B(n_16),
.Y(n_366)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_224),
.B(n_41),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_226),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_306),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_306),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_300),
.B(n_282),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_314),
.B(n_227),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_323),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_317),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_351),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_184),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_317),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_294),
.A2(n_249),
.B1(n_208),
.B2(n_260),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_364),
.A2(n_257),
.B1(n_291),
.B2(n_290),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_352),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_322),
.B(n_230),
.Y(n_385)
);

BUFx4f_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_185),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_232),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_342),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_296),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_293),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_235),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_298),
.B(n_259),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_292),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_331),
.B(n_279),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_314),
.B(n_244),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_327),
.B(n_236),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_327),
.B(n_340),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_367),
.Y(n_402)
);

OAI22xp33_ASAP7_75t_L g403 ( 
.A1(n_358),
.A2(n_196),
.B1(n_281),
.B2(n_280),
.Y(n_403)
);

OAI21xp33_ASAP7_75t_SL g404 ( 
.A1(n_340),
.A2(n_346),
.B(n_341),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_360),
.B(n_185),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_359),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_349),
.B(n_263),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_305),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_359),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_330),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_328),
.B(n_259),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_346),
.B(n_241),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_347),
.B(n_243),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_293),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_293),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

OR2x6_ASAP7_75t_L g419 ( 
.A(n_355),
.B(n_239),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g423 ( 
.A(n_348),
.B(n_248),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_348),
.A2(n_363),
.B1(n_367),
.B2(n_333),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_350),
.B(n_259),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_303),
.A2(n_254),
.B1(n_238),
.B2(n_234),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_299),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_297),
.Y(n_429)
);

AND3x2_ASAP7_75t_L g430 ( 
.A(n_356),
.B(n_267),
.C(n_265),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_363),
.B(n_269),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_318),
.B(n_234),
.Y(n_432)
);

NAND2xp33_ASAP7_75t_R g433 ( 
.A(n_307),
.B(n_289),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_338),
.B(n_270),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_297),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_333),
.B(n_271),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_338),
.B(n_275),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_299),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_302),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_334),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_302),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_325),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_353),
.A2(n_254),
.B1(n_238),
.B2(n_281),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_318),
.B(n_190),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_304),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_312),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_297),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_335),
.A2(n_354),
.B1(n_329),
.B2(n_366),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_L g450 ( 
.A(n_367),
.B(n_325),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_334),
.B(n_190),
.C(n_285),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_312),
.Y(n_452)
);

BUFx8_ASAP7_75t_SL g453 ( 
.A(n_321),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_337),
.B(n_274),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_412),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_410),
.B(n_368),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_389),
.B(n_339),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_378),
.A2(n_368),
.B1(n_361),
.B2(n_357),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_425),
.B(n_344),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_379),
.B(n_344),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g461 ( 
.A(n_386),
.B(n_307),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_387),
.B(n_449),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_413),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_436),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_276),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

NOR3xp33_ASAP7_75t_L g467 ( 
.A(n_382),
.B(n_332),
.C(n_311),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_422),
.B(n_278),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_405),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_400),
.B(n_372),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_436),
.B(n_283),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_384),
.B(n_311),
.Y(n_472)
);

BUFx6f_ASAP7_75t_SL g473 ( 
.A(n_384),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_372),
.B(n_383),
.Y(n_474)
);

INVx8_ASAP7_75t_L g475 ( 
.A(n_419),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_408),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_383),
.B(n_285),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_428),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_418),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_424),
.B(n_192),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_395),
.B(n_202),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_295),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_395),
.B(n_204),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_396),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_407),
.B(n_308),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_393),
.B(n_308),
.Y(n_487)
);

OR2x6_ASAP7_75t_L g488 ( 
.A(n_406),
.B(n_273),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_399),
.B(n_213),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_376),
.Y(n_491)
);

OAI221xp5_ASAP7_75t_L g492 ( 
.A1(n_404),
.A2(n_326),
.B1(n_324),
.B2(n_320),
.C(n_313),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_401),
.B(n_217),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_390),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_397),
.B(n_218),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_381),
.A2(n_324),
.B1(n_326),
.B2(n_320),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_385),
.B(n_221),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_385),
.B(n_231),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_440),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_445),
.B(n_343),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_442),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_369),
.B(n_233),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_370),
.A2(n_345),
.B1(n_307),
.B2(n_310),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_446),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_447),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_452),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g508 ( 
.A(n_451),
.B(n_16),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_375),
.B(n_246),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_430),
.B(n_253),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_373),
.B(n_392),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_423),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_423),
.A2(n_261),
.B1(n_258),
.B2(n_288),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_423),
.A2(n_310),
.B1(n_301),
.B2(n_319),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_431),
.B(n_262),
.Y(n_515)
);

AND2x2_ASAP7_75t_SL g516 ( 
.A(n_427),
.B(n_310),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_431),
.B(n_264),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_398),
.A2(n_310),
.B(n_219),
.Y(n_518)
);

O2A1O1Ixp33_ASAP7_75t_L g519 ( 
.A1(n_398),
.A2(n_17),
.B(n_18),
.C(n_21),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_414),
.B(n_309),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_414),
.B(n_18),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_415),
.B(n_377),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_415),
.B(n_309),
.Y(n_523)
);

O2A1O1Ixp5_ASAP7_75t_L g524 ( 
.A1(n_518),
.A2(n_388),
.B(n_434),
.C(n_438),
.Y(n_524)
);

A2O1A1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_462),
.A2(n_388),
.B(n_438),
.C(n_434),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_L g526 ( 
.A1(n_511),
.A2(n_443),
.B(n_426),
.C(n_421),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_469),
.B(n_437),
.Y(n_527)
);

AO21x1_ASAP7_75t_L g528 ( 
.A1(n_519),
.A2(n_433),
.B(n_371),
.Y(n_528)
);

O2A1O1Ixp33_ASAP7_75t_L g529 ( 
.A1(n_474),
.A2(n_403),
.B(n_426),
.C(n_420),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_469),
.B(n_437),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_432),
.Y(n_531)
);

AOI21xp33_ASAP7_75t_L g532 ( 
.A1(n_477),
.A2(n_433),
.B(n_403),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_486),
.B(n_432),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_512),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_463),
.B(n_453),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_463),
.B(n_23),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_475),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_461),
.A2(n_470),
.B(n_504),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_459),
.B(n_430),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_473),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_494),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_472),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_459),
.B(n_24),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_491),
.B(n_24),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_491),
.A2(n_516),
.B1(n_458),
.B2(n_492),
.Y(n_545)
);

CKINVDCx10_ASAP7_75t_R g546 ( 
.A(n_473),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_461),
.A2(n_380),
.B(n_374),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_475),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_475),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_464),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_504),
.A2(n_416),
.B(n_391),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_487),
.B(n_26),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_500),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_522),
.A2(n_460),
.B(n_514),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_466),
.B(n_26),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_499),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_456),
.B(n_30),
.Y(n_558)
);

NAND2x1p5_ASAP7_75t_L g559 ( 
.A(n_521),
.B(n_309),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_465),
.Y(n_560)
);

AOI21x1_ASAP7_75t_L g561 ( 
.A1(n_481),
.A2(n_417),
.B(n_435),
.Y(n_561)
);

OA22x2_ASAP7_75t_L g562 ( 
.A1(n_488),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_562)
);

AO22x1_ASAP7_75t_L g563 ( 
.A1(n_521),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_563)
);

A2O1A1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_457),
.A2(n_319),
.B(n_316),
.C(n_429),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_478),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_468),
.A2(n_493),
.B(n_489),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_458),
.A2(n_496),
.B1(n_490),
.B2(n_506),
.Y(n_567)
);

OAI21xp33_ASAP7_75t_L g568 ( 
.A1(n_497),
.A2(n_319),
.B(n_316),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_496),
.A2(n_319),
.B1(n_316),
.B2(n_448),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_495),
.B(n_42),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_479),
.A2(n_448),
.B(n_316),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_510),
.B(n_43),
.Y(n_572)
);

BUFx8_ASAP7_75t_L g573 ( 
.A(n_501),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_488),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_503),
.A2(n_53),
.B(n_54),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_515),
.B(n_176),
.Y(n_576)
);

OAI221xp5_ASAP7_75t_L g577 ( 
.A1(n_467),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.C(n_66),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_480),
.A2(n_67),
.B(n_71),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_483),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_509),
.A2(n_74),
.B(n_77),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_471),
.A2(n_80),
.B(n_83),
.Y(n_581)
);

A2O1A1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_505),
.A2(n_84),
.B(n_88),
.C(n_91),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_502),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_517),
.A2(n_100),
.B(n_101),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_498),
.B(n_103),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_513),
.B(n_107),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_488),
.B(n_110),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_476),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_507),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_520),
.A2(n_118),
.B(n_123),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_538),
.A2(n_484),
.B(n_482),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_555),
.A2(n_523),
.B(n_520),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_540),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_542),
.B(n_508),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_547),
.B(n_523),
.Y(n_595)
);

OAI22x1_ASAP7_75t_L g596 ( 
.A1(n_535),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_565),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_560),
.B(n_128),
.Y(n_598)
);

AO21x2_ASAP7_75t_L g599 ( 
.A1(n_528),
.A2(n_133),
.B(n_134),
.Y(n_599)
);

OAI22x1_ASAP7_75t_L g600 ( 
.A1(n_574),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_566),
.A2(n_147),
.B(n_149),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_524),
.A2(n_151),
.B(n_156),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_550),
.B(n_537),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_540),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_545),
.A2(n_559),
.B1(n_544),
.B2(n_553),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_565),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_525),
.A2(n_567),
.B(n_529),
.Y(n_607)
);

AOI211x1_ASAP7_75t_L g608 ( 
.A1(n_532),
.A2(n_545),
.B(n_563),
.C(n_577),
.Y(n_608)
);

AO21x2_ASAP7_75t_L g609 ( 
.A1(n_578),
.A2(n_564),
.B(n_590),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_SL g610 ( 
.A(n_533),
.B(n_531),
.C(n_572),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_549),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_557),
.B(n_554),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_573),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_573),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_589),
.B(n_558),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_536),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_587),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_527),
.A2(n_530),
.B(n_576),
.Y(n_618)
);

AO21x2_ASAP7_75t_L g619 ( 
.A1(n_590),
.A2(n_571),
.B(n_568),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_588),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_551),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_541),
.B(n_543),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_539),
.B(n_556),
.Y(n_623)
);

AO21x1_ASAP7_75t_L g624 ( 
.A1(n_586),
.A2(n_584),
.B(n_575),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_546),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_562),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_551),
.B(n_570),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_534),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_562),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_534),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_580),
.A2(n_569),
.B(n_581),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_545),
.A2(n_559),
.B1(n_516),
.B2(n_544),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_583),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_589),
.Y(n_634)
);

A2O1A1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_529),
.A2(n_462),
.B(n_566),
.C(n_511),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_583),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_548),
.A2(n_552),
.B(n_561),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_579),
.B(n_462),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_538),
.A2(n_462),
.B(n_555),
.Y(n_639)
);

NOR3xp33_ASAP7_75t_L g640 ( 
.A(n_533),
.B(n_531),
.C(n_535),
.Y(n_640)
);

AO31x2_ASAP7_75t_L g641 ( 
.A1(n_528),
.A2(n_538),
.A3(n_545),
.B(n_564),
.Y(n_641)
);

AO22x2_ASAP7_75t_L g642 ( 
.A1(n_545),
.A2(n_444),
.B1(n_536),
.B2(n_485),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_589),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_583),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_572),
.B(n_402),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_540),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_579),
.B(n_462),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_538),
.A2(n_450),
.B(n_394),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_579),
.B(n_550),
.Y(n_649)
);

AO31x2_ASAP7_75t_L g650 ( 
.A1(n_528),
.A2(n_538),
.A3(n_545),
.B(n_564),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_572),
.B(n_402),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_538),
.A2(n_450),
.B(n_394),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_542),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_538),
.A2(n_450),
.B(n_394),
.Y(n_654)
);

OAI22x1_ASAP7_75t_L g655 ( 
.A1(n_535),
.A2(n_318),
.B1(n_321),
.B2(n_427),
.Y(n_655)
);

BUFx2_ASAP7_75t_R g656 ( 
.A(n_549),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_589),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_579),
.B(n_462),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_583),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_573),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_SL g661 ( 
.A1(n_576),
.A2(n_585),
.B(n_526),
.C(n_582),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_579),
.B(n_462),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_565),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_613),
.Y(n_664)
);

AOI21xp33_ASAP7_75t_SL g665 ( 
.A1(n_625),
.A2(n_614),
.B(n_655),
.Y(n_665)
);

NOR2xp67_ASAP7_75t_L g666 ( 
.A(n_593),
.B(n_646),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_638),
.B(n_647),
.Y(n_667)
);

AO31x2_ASAP7_75t_L g668 ( 
.A1(n_605),
.A2(n_632),
.A3(n_635),
.B(n_624),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_662),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_660),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_653),
.B(n_623),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_616),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_634),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_636),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_644),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_626),
.B(n_629),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_642),
.B(n_615),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_659),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_620),
.Y(n_679)
);

OA21x2_ASAP7_75t_L g680 ( 
.A1(n_607),
.A2(n_639),
.B(n_602),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_643),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_657),
.Y(n_682)
);

NAND2x1p5_ASAP7_75t_L g683 ( 
.A(n_597),
.B(n_606),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_642),
.B(n_640),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_603),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g686 ( 
.A1(n_648),
.A2(n_654),
.B(n_652),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_592),
.A2(n_591),
.B(n_595),
.Y(n_687)
);

CKINVDCx6p67_ASAP7_75t_R g688 ( 
.A(n_604),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_603),
.B(n_612),
.Y(n_689)
);

OA21x2_ASAP7_75t_L g690 ( 
.A1(n_592),
.A2(n_631),
.B(n_618),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_622),
.B(n_595),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_663),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_645),
.A2(n_651),
.B(n_610),
.C(n_601),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_611),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_617),
.B(n_612),
.Y(n_695)
);

OR3x4_ASAP7_75t_SL g696 ( 
.A(n_656),
.B(n_611),
.C(n_617),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_608),
.B(n_650),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_594),
.A2(n_598),
.B(n_650),
.Y(n_698)
);

OA21x2_ASAP7_75t_L g699 ( 
.A1(n_641),
.A2(n_650),
.B(n_599),
.Y(n_699)
);

AO31x2_ASAP7_75t_L g700 ( 
.A1(n_600),
.A2(n_596),
.A3(n_641),
.B(n_609),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_645),
.A2(n_651),
.B(n_661),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_628),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_630),
.B(n_641),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_627),
.Y(n_704)
);

AO21x2_ASAP7_75t_L g705 ( 
.A1(n_609),
.A2(n_599),
.B(n_619),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_627),
.A2(n_608),
.B(n_619),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_635),
.A2(n_538),
.B(n_639),
.Y(n_707)
);

AO31x2_ASAP7_75t_L g708 ( 
.A1(n_605),
.A2(n_632),
.A3(n_528),
.B(n_635),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_621),
.Y(n_709)
);

BUFx4_ASAP7_75t_SL g710 ( 
.A(n_613),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_634),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_613),
.Y(n_712)
);

OA21x2_ASAP7_75t_L g713 ( 
.A1(n_607),
.A2(n_639),
.B(n_637),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_649),
.B(n_579),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_649),
.B(n_579),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_642),
.A2(n_640),
.B1(n_626),
.B2(n_629),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_633),
.Y(n_717)
);

AO21x2_ASAP7_75t_L g718 ( 
.A1(n_607),
.A2(n_639),
.B(n_605),
.Y(n_718)
);

OA21x2_ASAP7_75t_L g719 ( 
.A1(n_607),
.A2(n_639),
.B(n_637),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_649),
.B(n_579),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_613),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_638),
.B(n_647),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_633),
.Y(n_723)
);

AO21x2_ASAP7_75t_L g724 ( 
.A1(n_607),
.A2(n_639),
.B(n_605),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_633),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_638),
.B(n_647),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_633),
.Y(n_727)
);

BUFx4f_ASAP7_75t_SL g728 ( 
.A(n_625),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_653),
.B(n_485),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_633),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_638),
.B(n_647),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_633),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_676),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_704),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_674),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_675),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_684),
.B(n_677),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_671),
.B(n_673),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_671),
.B(n_681),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_678),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_679),
.Y(n_741)
);

BUFx2_ASAP7_75t_SL g742 ( 
.A(n_666),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_717),
.Y(n_743)
);

AO21x2_ASAP7_75t_L g744 ( 
.A1(n_686),
.A2(n_707),
.B(n_706),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_682),
.B(n_711),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_723),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_665),
.B(n_695),
.C(n_722),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_725),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_727),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_709),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_709),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_688),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_730),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_710),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_732),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_716),
.B(n_691),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_710),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_667),
.A2(n_731),
.B1(n_726),
.B2(n_669),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_691),
.B(n_676),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_731),
.B(n_667),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_672),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_709),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_714),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_729),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_669),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_703),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_728),
.Y(n_768)
);

BUFx2_ASAP7_75t_SL g769 ( 
.A(n_714),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_715),
.Y(n_770)
);

OA21x2_ASAP7_75t_L g771 ( 
.A1(n_706),
.A2(n_707),
.B(n_698),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_701),
.B(n_687),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_704),
.B(n_683),
.Y(n_773)
);

NOR2x1_ASAP7_75t_R g774 ( 
.A(n_664),
.B(n_670),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_720),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_704),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_689),
.B(n_712),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_718),
.B(n_724),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_695),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_702),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_697),
.B(n_718),
.Y(n_781)
);

AO21x2_ASAP7_75t_L g782 ( 
.A1(n_705),
.A2(n_693),
.B(n_724),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_685),
.Y(n_783)
);

INVx4_ASAP7_75t_R g784 ( 
.A(n_755),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_778),
.B(n_708),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_781),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_761),
.B(n_708),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_733),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_761),
.B(n_708),
.Y(n_789)
);

INVx3_ASAP7_75t_SL g790 ( 
.A(n_773),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_766),
.B(n_664),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_757),
.A2(n_721),
.B1(n_670),
.B2(n_680),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_747),
.B(n_694),
.C(n_692),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_778),
.B(n_719),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_767),
.B(n_737),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_738),
.B(n_713),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_774),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_739),
.B(n_744),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_739),
.B(n_668),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_765),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_SL g801 ( 
.A(n_758),
.B(n_728),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_748),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_760),
.B(n_700),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_760),
.B(n_699),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_759),
.B(n_699),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_769),
.B(n_690),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_741),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_745),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_745),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_801),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_798),
.B(n_804),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_808),
.B(n_809),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_787),
.A2(n_779),
.B1(n_762),
.B2(n_755),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_798),
.B(n_771),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_788),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_804),
.B(n_771),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_788),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_803),
.B(n_771),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_802),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_803),
.B(n_782),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_807),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_800),
.B(n_754),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_799),
.B(n_782),
.Y(n_823)
);

AND2x2_ASAP7_75t_SL g824 ( 
.A(n_807),
.B(n_734),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_787),
.B(n_756),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_789),
.B(n_746),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_790),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_811),
.B(n_794),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_824),
.A2(n_806),
.B(n_772),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_811),
.B(n_818),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_818),
.B(n_794),
.Y(n_831)
);

INVxp67_ASAP7_75t_SL g832 ( 
.A(n_821),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_819),
.B(n_789),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_815),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_815),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_814),
.B(n_785),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_814),
.B(n_785),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_817),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_825),
.B(n_795),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_816),
.B(n_785),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_820),
.B(n_796),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_826),
.B(n_786),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_830),
.B(n_831),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_834),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_834),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_830),
.B(n_812),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_832),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_841),
.B(n_823),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_835),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_835),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_828),
.B(n_820),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_838),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_829),
.A2(n_824),
.B(n_797),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_841),
.B(n_828),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_847),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_853),
.A2(n_810),
.B1(n_824),
.B2(n_833),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_846),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_843),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_851),
.A2(n_836),
.B1(n_837),
.B2(n_840),
.Y(n_859)
);

OAI21xp33_ASAP7_75t_L g860 ( 
.A1(n_843),
.A2(n_836),
.B(n_837),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_844),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_SL g862 ( 
.A1(n_845),
.A2(n_793),
.B(n_780),
.C(n_777),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_851),
.B(n_831),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_849),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_L g865 ( 
.A(n_850),
.B(n_822),
.C(n_813),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_846),
.Y(n_866)
);

AOI211xp5_ASAP7_75t_SL g867 ( 
.A1(n_856),
.A2(n_784),
.B(n_696),
.C(n_805),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_860),
.B(n_827),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_861),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_859),
.A2(n_854),
.B1(n_848),
.B2(n_827),
.Y(n_870)
);

AOI211xp5_ASAP7_75t_L g871 ( 
.A1(n_862),
.A2(n_790),
.B(n_753),
.C(n_768),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_857),
.A2(n_827),
.B1(n_790),
.B2(n_839),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_858),
.B(n_866),
.Y(n_873)
);

OAI221xp5_ASAP7_75t_L g874 ( 
.A1(n_867),
.A2(n_855),
.B1(n_862),
.B2(n_865),
.C(n_864),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_869),
.B(n_855),
.Y(n_875)
);

AOI211xp5_ASAP7_75t_L g876 ( 
.A1(n_872),
.A2(n_871),
.B(n_868),
.C(n_870),
.Y(n_876)
);

OAI211xp5_ASAP7_75t_SL g877 ( 
.A1(n_876),
.A2(n_792),
.B(n_873),
.C(n_791),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_875),
.Y(n_878)
);

NAND4xp75_ASAP7_75t_L g879 ( 
.A(n_877),
.B(n_696),
.C(n_874),
.D(n_753),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_SL g880 ( 
.A(n_878),
.B(n_768),
.C(n_784),
.Y(n_880)
);

AND3x4_ASAP7_75t_L g881 ( 
.A(n_880),
.B(n_764),
.C(n_775),
.Y(n_881)
);

NAND4xp75_ASAP7_75t_L g882 ( 
.A(n_879),
.B(n_742),
.C(n_776),
.D(n_863),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_882),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_881),
.Y(n_884)
);

XNOR2x1_ASAP7_75t_L g885 ( 
.A(n_883),
.B(n_742),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_884),
.B(n_842),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_883),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_887),
.B(n_852),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_885),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_886),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_887),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_SL g892 ( 
.A1(n_887),
.A2(n_734),
.B1(n_776),
.B2(n_773),
.Y(n_892)
);

XNOR2xp5_ASAP7_75t_L g893 ( 
.A(n_889),
.B(n_770),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_892),
.A2(n_734),
.B1(n_769),
.B2(n_783),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_891),
.A2(n_752),
.B(n_763),
.Y(n_895)
);

AOI22x1_ASAP7_75t_L g896 ( 
.A1(n_890),
.A2(n_752),
.B1(n_751),
.B2(n_763),
.Y(n_896)
);

AOI21xp33_ASAP7_75t_L g897 ( 
.A1(n_888),
.A2(n_749),
.B(n_743),
.Y(n_897)
);

OR2x6_ASAP7_75t_L g898 ( 
.A(n_891),
.B(n_773),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_896),
.Y(n_899)
);

AOI21xp33_ASAP7_75t_L g900 ( 
.A1(n_893),
.A2(n_735),
.B(n_740),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_895),
.A2(n_750),
.B(n_736),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_899),
.B(n_898),
.Y(n_902)
);

OA21x2_ASAP7_75t_L g903 ( 
.A1(n_902),
.A2(n_900),
.B(n_897),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_903),
.A2(n_901),
.B(n_894),
.Y(n_904)
);


endmodule