module fake_jpeg_32161_n_455 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_455);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_455;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_51),
.B(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_45),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_17),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_89),
.Y(n_111)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_70),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_86),
.Y(n_133)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_30),
.Y(n_131)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_37),
.B(n_16),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_45),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_131),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_53),
.B(n_0),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_20),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_67),
.A2(n_46),
.B1(n_44),
.B2(n_19),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_46),
.B1(n_31),
.B2(n_38),
.Y(n_141)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

AO21x2_ASAP7_75t_SL g192 ( 
.A1(n_141),
.A2(n_143),
.B(n_114),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_60),
.B1(n_66),
.B2(n_62),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_147),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_65),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_172),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_102),
.A2(n_54),
.B1(n_80),
.B2(n_85),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_149),
.A2(n_164),
.B1(n_169),
.B2(n_114),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_151),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_98),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_153),
.B(n_155),
.Y(n_207)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_30),
.B(n_31),
.C(n_20),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_75),
.B1(n_74),
.B2(n_63),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_171),
.B1(n_175),
.B2(n_36),
.Y(n_182)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_157),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_160),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_46),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_50),
.B1(n_31),
.B2(n_44),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_140),
.B1(n_137),
.B2(n_121),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_113),
.A2(n_19),
.B1(n_44),
.B2(n_23),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_168),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_117),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_105),
.A2(n_26),
.B1(n_38),
.B2(n_36),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_24),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_124),
.B(n_42),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_174),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_115),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_116),
.A2(n_23),
.B1(n_38),
.B2(n_36),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_138),
.B(n_42),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_32),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_51),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_177),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_192),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_119),
.B1(n_116),
.B2(n_130),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_96),
.B(n_136),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_176),
.B(n_160),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_195),
.B(n_145),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_138),
.C(n_98),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_143),
.C(n_151),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_143),
.A2(n_119),
.B1(n_130),
.B2(n_137),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_204),
.B1(n_147),
.B2(n_162),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_200),
.A2(n_170),
.B1(n_144),
.B2(n_178),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_140),
.B1(n_103),
.B2(n_134),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_20),
.B(n_19),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_155),
.B(n_148),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_100),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_147),
.Y(n_221)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_210),
.A2(n_212),
.B(n_214),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_230),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_174),
.B1(n_143),
.B2(n_152),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_213),
.A2(n_225),
.B(n_189),
.Y(n_252)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_142),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_223),
.Y(n_253)
);

BUFx4f_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_219),
.A2(n_189),
.B1(n_179),
.B2(n_199),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_187),
.B1(n_162),
.B2(n_166),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_221),
.B(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_183),
.B(n_145),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_173),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_228),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_157),
.B(n_178),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_152),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_193),
.B(n_158),
.Y(n_228)
);

NAND2x1p5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_127),
.Y(n_229)
);

AO21x2_ASAP7_75t_SL g242 ( 
.A1(n_229),
.A2(n_221),
.B(n_230),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_167),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_168),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_193),
.C(n_203),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_154),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_226),
.A2(n_192),
.B1(n_200),
.B2(n_198),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_256),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_186),
.B(n_192),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_211),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_210),
.A2(n_205),
.B(n_190),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_237),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_240),
.C(n_246),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_203),
.C(n_197),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_242),
.A2(n_247),
.B(n_252),
.Y(n_285)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_194),
.C(n_185),
.Y(n_246)
);

AO21x2_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_182),
.B(n_204),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_195),
.C(n_184),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_255),
.C(n_227),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_187),
.C(n_161),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_202),
.B(n_189),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_226),
.B1(n_239),
.B2(n_215),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_SL g258 ( 
.A(n_237),
.B(n_229),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_258),
.A2(n_259),
.B(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_262),
.A2(n_267),
.B1(n_247),
.B2(n_240),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_248),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_263),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_222),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_264),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_254),
.B(n_228),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_265),
.B(n_269),
.Y(n_289)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_212),
.B1(n_232),
.B2(n_220),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_248),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_270),
.B(n_255),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_235),
.A2(n_229),
.B1(n_208),
.B2(n_217),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_247),
.B1(n_257),
.B2(n_242),
.Y(n_293)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

OAI22x1_ASAP7_75t_L g274 ( 
.A1(n_236),
.A2(n_217),
.B1(n_202),
.B2(n_209),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_217),
.Y(n_275)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_246),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_280),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_245),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_284),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_201),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_283),
.B(n_250),
.Y(n_305)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_245),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_219),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_268),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_278),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_233),
.C(n_238),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_308),
.C(n_314),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_293),
.A2(n_300),
.B1(n_307),
.B2(n_312),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_233),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_310),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_271),
.A2(n_247),
.B1(n_242),
.B2(n_250),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_302),
.B(n_263),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_291),
.B1(n_303),
.B2(n_316),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_285),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_247),
.B1(n_242),
.B2(n_253),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_253),
.C(n_243),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_188),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_179),
.B1(n_181),
.B2(n_199),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_313),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_267),
.B(n_188),
.C(n_152),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_139),
.C(n_218),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_316),
.C(n_284),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_136),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_317),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_318),
.A2(n_327),
.B1(n_335),
.B2(n_320),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_264),
.Y(n_319)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_319),
.Y(n_358)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_294),
.A2(n_265),
.B(n_275),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g364 ( 
.A(n_321),
.B(n_16),
.C(n_15),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_281),
.Y(n_322)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_307),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_336),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_269),
.C(n_279),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_331),
.C(n_332),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_285),
.B1(n_262),
.B2(n_277),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_329),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_308),
.B(n_260),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_285),
.C(n_273),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_272),
.C(n_266),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_334),
.A2(n_191),
.B(n_96),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_291),
.A2(n_277),
.B1(n_278),
.B2(n_179),
.Y(n_335)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_24),
.C(n_22),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_302),
.B(n_290),
.C(n_314),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_299),
.C(n_139),
.Y(n_353)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_340),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_341),
.A2(n_301),
.B1(n_332),
.B2(n_335),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_334),
.A2(n_313),
.B(n_315),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_342),
.B(n_353),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_326),
.B(n_295),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_362),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_359),
.C(n_337),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_330),
.A2(n_300),
.B1(n_293),
.B2(n_306),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_347),
.A2(n_350),
.B1(n_355),
.B2(n_356),
.Y(n_378)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_348),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_349),
.A2(n_99),
.B1(n_22),
.B2(n_95),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_299),
.B1(n_297),
.B2(n_312),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_334),
.A2(n_199),
.B1(n_191),
.B2(n_166),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_327),
.A2(n_191),
.B1(n_169),
.B2(n_165),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_337),
.C(n_331),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_324),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_16),
.B(n_15),
.Y(n_362)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_97),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_365),
.B(n_159),
.Y(n_369)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_366),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_369),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_358),
.A2(n_338),
.B1(n_336),
.B2(n_325),
.Y(n_368)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_368),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_349),
.A2(n_165),
.B1(n_146),
.B2(n_169),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_370),
.A2(n_373),
.B1(n_375),
.B2(n_382),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_360),
.Y(n_371)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_357),
.A2(n_146),
.B1(n_112),
.B2(n_104),
.Y(n_373)
);

A2O1A1Ixp33_ASAP7_75t_SL g375 ( 
.A1(n_347),
.A2(n_112),
.B(n_104),
.C(n_159),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_99),
.C(n_93),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_385),
.C(n_359),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_363),
.B(n_24),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_381),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_350),
.A2(n_93),
.B1(n_22),
.B2(n_23),
.Y(n_381)
);

XOR2x1_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_0),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_383),
.A2(n_384),
.B(n_355),
.Y(n_398)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_123),
.C(n_94),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_362),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_373),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_387),
.B(n_389),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_345),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_374),
.A2(n_342),
.B(n_352),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_391),
.A2(n_396),
.B(n_399),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_365),
.C(n_353),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_393),
.C(n_401),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_346),
.Y(n_393)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_394),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_378),
.A2(n_352),
.B(n_361),
.Y(n_396)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_398),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_356),
.B(n_351),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_354),
.C(n_26),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_402),
.A2(n_400),
.B1(n_390),
.B2(n_395),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_388),
.A2(n_372),
.B(n_385),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_406),
.A2(n_2),
.B(n_4),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_391),
.A2(n_396),
.B(n_399),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_1),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g410 ( 
.A(n_403),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_410),
.B(n_2),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_402),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_370),
.C(n_382),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_412),
.B(n_1),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_394),
.A2(n_371),
.B1(n_375),
.B2(n_383),
.Y(n_413)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_413),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_387),
.B(n_386),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_409),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_400),
.A2(n_375),
.B1(n_2),
.B2(n_3),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_416),
.A2(n_408),
.B1(n_375),
.B2(n_397),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_420),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_419),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_414),
.B(n_392),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_409),
.A2(n_401),
.B(n_393),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_416),
.B(n_6),
.Y(n_435)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_422),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_424),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_1),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_426),
.Y(n_436)
);

AOI31xp33_ASAP7_75t_L g427 ( 
.A1(n_410),
.A2(n_404),
.A3(n_407),
.B(n_405),
.Y(n_427)
);

AOI322xp5_ASAP7_75t_L g431 ( 
.A1(n_427),
.A2(n_417),
.A3(n_405),
.B1(n_419),
.B2(n_422),
.C1(n_418),
.C2(n_411),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_428),
.B(n_5),
.Y(n_438)
);

OAI21x1_ASAP7_75t_SL g441 ( 
.A1(n_431),
.A2(n_5),
.B(n_7),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_412),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_432),
.B(n_437),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_435),
.A2(n_5),
.B(n_7),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_5),
.C(n_6),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_438),
.B(n_429),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g448 ( 
.A1(n_439),
.A2(n_441),
.B(n_443),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_430),
.Y(n_440)
);

AOI322xp5_ASAP7_75t_L g446 ( 
.A1(n_440),
.A2(n_433),
.A3(n_436),
.B1(n_10),
.B2(n_11),
.C1(n_8),
.C2(n_14),
.Y(n_446)
);

AOI21x1_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_7),
.B(n_8),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_442),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_437),
.B(n_8),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_444),
.A2(n_433),
.B1(n_10),
.B2(n_11),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_449),
.C(n_445),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_450),
.Y(n_452)
);

AOI321xp33_ASAP7_75t_L g451 ( 
.A1(n_447),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_448),
.C(n_427),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_451),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_453),
.B(n_9),
.Y(n_454)
);

BUFx24_ASAP7_75t_SL g455 ( 
.A(n_454),
.Y(n_455)
);


endmodule