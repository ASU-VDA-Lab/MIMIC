module real_jpeg_1916_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_11;
wire n_14;
wire n_7;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

AND2x2_ASAP7_75t_SL g14 ( 
.A(n_1),
.B(n_15),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_10),
.Y(n_9)
);

NAND2x1_ASAP7_75t_SL g11 ( 
.A(n_5),
.B(n_10),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_12),
.B1(n_13),
.B2(n_21),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_9),
.B(n_11),
.Y(n_7)
);

CKINVDCx14_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_17),
.B(n_18),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_16),
.B(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);


endmodule