module fake_aes_2703_n_668 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_668);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_668;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx14_ASAP7_75t_R g77 ( .A(n_12), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_59), .Y(n_78) );
NOR2xp67_ASAP7_75t_L g79 ( .A(n_4), .B(n_41), .Y(n_79) );
BUFx6f_ASAP7_75t_L g80 ( .A(n_68), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_1), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_17), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_50), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_53), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_3), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_40), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_63), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_75), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_27), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_20), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_65), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_76), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_36), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_38), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_3), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_43), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_67), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_74), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_52), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_62), .Y(n_100) );
INVxp33_ASAP7_75t_L g101 ( .A(n_46), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_71), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_19), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_6), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_73), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_48), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_45), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_16), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_15), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_25), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_5), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_1), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_47), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_60), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_44), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_15), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_14), .Y(n_118) );
XNOR2xp5_ASAP7_75t_L g119 ( .A(n_37), .B(n_35), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_72), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_54), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_56), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_26), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_82), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_78), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_77), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_104), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_83), .Y(n_132) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_107), .A2(n_28), .B(n_69), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_81), .B(n_0), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_87), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_87), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_105), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_80), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_105), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_99), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_81), .B(n_2), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_94), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_84), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_107), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_84), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_85), .B(n_2), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_95), .B(n_4), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_94), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_88), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_95), .B(n_5), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_119), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_119), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_117), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_99), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_90), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_90), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_91), .B(n_6), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_101), .B(n_7), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
BUFx4_ASAP7_75t_L g166 ( .A(n_134), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_150), .B(n_117), .Y(n_167) );
NAND2x1p5_ASAP7_75t_L g168 ( .A(n_125), .B(n_123), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
INVx3_ASAP7_75t_R g170 ( .A(n_149), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_136), .B(n_111), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_130), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_150), .B(n_109), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_125), .B(n_112), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_126), .B(n_118), .Y(n_176) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_164), .B(n_113), .C(n_122), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_146), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_137), .B(n_103), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_126), .B(n_122), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
OAI221xp5_ASAP7_75t_L g186 ( .A1(n_134), .A2(n_110), .B1(n_89), .B2(n_120), .C(n_121), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_132), .B(n_123), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_160), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_131), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_164), .A2(n_120), .B1(n_91), .B2(n_92), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_132), .B(n_121), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_164), .B(n_116), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_135), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_154), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_157), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_135), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_135), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_138), .B(n_92), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_140), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_138), .B(n_115), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_146), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_145), .B(n_98), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_144), .B(n_114), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_145), .B(n_97), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_153), .B(n_108), .Y(n_211) );
NAND3x1_ASAP7_75t_L g212 ( .A(n_143), .B(n_93), .C(n_102), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_129), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_129), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_147), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_140), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_127), .B(n_106), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_147), .B(n_100), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_152), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_152), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_161), .B(n_93), .Y(n_222) );
OR2x6_ASAP7_75t_L g223 ( .A(n_166), .B(n_143), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_168), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_179), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_177), .B(n_151), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_179), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_168), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_167), .B(n_151), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_187), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_181), .Y(n_232) );
AND2x6_ASAP7_75t_L g233 ( .A(n_193), .B(n_162), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_181), .Y(n_234) );
BUFx4f_ASAP7_75t_SL g235 ( .A(n_190), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_187), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_173), .B(n_128), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g238 ( .A(n_186), .B(n_162), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_173), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_188), .Y(n_240) );
NOR2xp33_ASAP7_75t_R g241 ( .A(n_190), .B(n_156), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_188), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_194), .B(n_161), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_179), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_183), .B(n_124), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_182), .Y(n_246) );
BUFx4f_ASAP7_75t_SL g247 ( .A(n_167), .Y(n_247) );
INVxp67_ASAP7_75t_SL g248 ( .A(n_166), .Y(n_248) );
NAND2xp33_ASAP7_75t_L g249 ( .A(n_212), .B(n_96), .Y(n_249) );
NOR3xp33_ASAP7_75t_SL g250 ( .A(n_171), .B(n_158), .C(n_163), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_193), .B(n_142), .Y(n_251) );
NOR3xp33_ASAP7_75t_SL g252 ( .A(n_209), .B(n_148), .C(n_155), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_193), .B(n_155), .Y(n_253) );
BUFx2_ASAP7_75t_L g254 ( .A(n_212), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_222), .B(n_176), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_167), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_222), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_211), .B(n_148), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_182), .Y(n_259) );
NOR3xp33_ASAP7_75t_SL g260 ( .A(n_218), .B(n_79), .C(n_8), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_195), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_182), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_195), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_185), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_176), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_196), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_174), .B(n_133), .Y(n_267) );
XNOR2xp5_ASAP7_75t_L g268 ( .A(n_192), .B(n_7), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_174), .B(n_133), .Y(n_269) );
INVxp67_ASAP7_75t_L g270 ( .A(n_204), .Y(n_270) );
BUFx12f_ASAP7_75t_L g271 ( .A(n_222), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_176), .B(n_159), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_176), .B(n_159), .Y(n_273) );
NOR3xp33_ASAP7_75t_SL g274 ( .A(n_219), .B(n_9), .C(n_10), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_174), .B(n_159), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_184), .B(n_159), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_196), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_198), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_184), .B(n_141), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_204), .B(n_139), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_184), .A2(n_141), .B1(n_139), .B2(n_133), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_184), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_189), .B(n_141), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_230), .B(n_189), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_224), .B(n_189), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_226), .B(n_189), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_229), .B(n_221), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_271), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_233), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_265), .B(n_221), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_265), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_230), .A2(n_220), .B1(n_216), .B2(n_200), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_282), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_239), .A2(n_206), .B1(n_208), .B2(n_210), .C(n_220), .Y(n_294) );
AND3x1_ASAP7_75t_SL g295 ( .A(n_268), .B(n_216), .C(n_207), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_237), .Y(n_296) );
AOI21xp5_ASAP7_75t_SL g297 ( .A1(n_267), .A2(n_185), .B(n_198), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_257), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_233), .Y(n_299) );
NAND2x2_ASAP7_75t_L g300 ( .A(n_241), .B(n_9), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_270), .B(n_207), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_230), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_271), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_227), .B(n_201), .Y(n_304) );
INVx5_ASAP7_75t_L g305 ( .A(n_233), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_282), .A2(n_199), .B1(n_139), .B2(n_141), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_223), .B(n_139), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_267), .A2(n_269), .B(n_253), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_233), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_248), .B(n_10), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_223), .B(n_11), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_233), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_256), .B(n_11), .Y(n_313) );
NOR2x1_ASAP7_75t_SL g314 ( .A(n_223), .B(n_170), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_232), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_243), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_236), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_247), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_252), .B(n_12), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_267), .B(n_217), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_236), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_256), .B(n_13), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_227), .B(n_13), .Y(n_323) );
OR2x6_ASAP7_75t_L g324 ( .A(n_255), .B(n_170), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_241), .B(n_14), .Y(n_325) );
NAND2x1_ASAP7_75t_L g326 ( .A(n_263), .B(n_217), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_269), .B(n_191), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_247), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_227), .B(n_280), .Y(n_329) );
AND2x2_ASAP7_75t_SL g330 ( .A(n_254), .B(n_16), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_235), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_317), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_316), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_297), .A2(n_281), .B(n_251), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_329), .A2(n_249), .B1(n_238), .B2(n_258), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_298), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_301), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_317), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_329), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_296), .B(n_272), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_293), .B(n_329), .Y(n_341) );
OR2x6_ASAP7_75t_L g342 ( .A(n_289), .B(n_269), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_330), .A2(n_249), .B1(n_258), .B2(n_245), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_293), .Y(n_344) );
NAND3xp33_ASAP7_75t_L g345 ( .A(n_294), .B(n_260), .C(n_250), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_292), .B(n_275), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_288), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_321), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_330), .A2(n_313), .B1(n_322), .B2(n_319), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_308), .A2(n_279), .B(n_276), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_292), .B(n_263), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_288), .B(n_273), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_320), .A2(n_231), .B(n_277), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_303), .B(n_278), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_289), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_289), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_311), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_300), .A2(n_235), .B1(n_278), .B2(n_266), .Y(n_358) );
OR2x6_ASAP7_75t_L g359 ( .A(n_289), .B(n_275), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_309), .B(n_283), .Y(n_360) );
AND2x6_ASAP7_75t_L g361 ( .A(n_309), .B(n_283), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_285), .A2(n_245), .B1(n_225), .B2(n_262), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_351), .B(n_287), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_345), .A2(n_319), .B1(n_307), .B2(n_325), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_337), .B(n_302), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_349), .A2(n_319), .B1(n_307), .B2(n_300), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_351), .B(n_287), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_342), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_346), .A2(n_307), .B1(n_323), .B2(n_310), .Y(n_369) );
INVxp33_ASAP7_75t_SL g370 ( .A(n_344), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_334), .A2(n_327), .B(n_320), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_332), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_334), .A2(n_327), .B(n_304), .Y(n_374) );
AO21x2_ASAP7_75t_L g375 ( .A1(n_350), .A2(n_321), .B(n_306), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_332), .A2(n_287), .B(n_284), .Y(n_376) );
NOR2xp67_ASAP7_75t_SL g377 ( .A(n_355), .B(n_305), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_343), .A2(n_286), .B1(n_285), .B2(n_302), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_338), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_333), .A2(n_285), .B1(n_286), .B2(n_318), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_357), .A2(n_286), .B1(n_291), .B2(n_261), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_358), .B(n_305), .Y(n_382) );
OAI21xp5_ASAP7_75t_SL g383 ( .A1(n_335), .A2(n_295), .B(n_331), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_339), .A2(n_328), .B1(n_312), .B2(n_225), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_341), .A2(n_312), .B1(n_259), .B2(n_262), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_338), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_341), .A2(n_295), .B1(n_314), .B2(n_305), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_342), .Y(n_388) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_359), .A2(n_324), .B(n_315), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_363), .B(n_354), .Y(n_390) );
BUFx2_ASAP7_75t_L g391 ( .A(n_372), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_387), .B(n_305), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_363), .B(n_342), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_365), .B(n_336), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_373), .Y(n_395) );
OAI21xp33_ASAP7_75t_L g396 ( .A1(n_364), .A2(n_274), .B(n_348), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_367), .B(n_348), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_365), .B(n_340), .Y(n_399) );
OAI221xp5_ASAP7_75t_SL g400 ( .A1(n_383), .A2(n_340), .B1(n_354), .B2(n_352), .C(n_362), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_366), .A2(n_347), .B1(n_352), .B2(n_353), .C(n_240), .Y(n_401) );
NOR3xp33_ASAP7_75t_L g402 ( .A(n_383), .B(n_350), .C(n_246), .Y(n_402) );
AND4x1_ASAP7_75t_L g403 ( .A(n_380), .B(n_242), .C(n_361), .D(n_324), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_379), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_369), .A2(n_360), .B1(n_359), .B2(n_290), .C(n_324), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_376), .A2(n_175), .B(n_165), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_378), .A2(n_360), .B1(n_359), .B2(n_290), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_376), .A2(n_299), .B(n_356), .C(n_246), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_379), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_373), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_368), .A2(n_360), .B1(n_359), .B2(n_299), .Y(n_412) );
AO21x2_ASAP7_75t_L g413 ( .A1(n_375), .A2(n_169), .B(n_165), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_369), .B(n_244), .C(n_259), .D(n_228), .Y(n_414) );
OA21x2_ASAP7_75t_L g415 ( .A1(n_371), .A2(n_169), .B(n_172), .Y(n_415) );
AND2x6_ASAP7_75t_L g416 ( .A(n_367), .B(n_355), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_386), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_386), .Y(n_418) );
OR2x6_ASAP7_75t_L g419 ( .A(n_368), .B(n_360), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_386), .B(n_356), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_387), .B(n_355), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_375), .Y(n_422) );
NAND3xp33_ASAP7_75t_SL g423 ( .A(n_381), .B(n_384), .C(n_382), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_411), .B(n_375), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_381), .B1(n_385), .B2(n_372), .C(n_388), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_395), .Y(n_427) );
BUFx12f_ASAP7_75t_L g428 ( .A(n_390), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_404), .Y(n_429) );
INVx4_ASAP7_75t_L g430 ( .A(n_416), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_411), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_410), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_395), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_418), .B(n_375), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_418), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_399), .B(n_390), .Y(n_436) );
INVx5_ASAP7_75t_L g437 ( .A(n_416), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_400), .B(n_389), .C(n_388), .D(n_244), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_410), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_423), .A2(n_361), .B1(n_388), .B2(n_374), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_394), .B(n_388), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_398), .B(n_406), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_416), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_398), .B(n_374), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_391), .Y(n_445) );
INVxp67_ASAP7_75t_L g446 ( .A(n_391), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_406), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_417), .B(n_374), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_421), .B(n_419), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_417), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g451 ( .A1(n_396), .A2(n_389), .B1(n_228), .B2(n_326), .C(n_234), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_403), .B(n_228), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_401), .A2(n_129), .B1(n_374), .B2(n_213), .C(n_205), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
INVxp67_ASAP7_75t_L g455 ( .A(n_420), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_422), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_421), .B(n_371), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_422), .B(n_371), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_419), .B(n_355), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_419), .B(n_315), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_402), .B(n_129), .C(n_377), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_419), .B(n_413), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_413), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_393), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_413), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_393), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_393), .B(n_129), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_403), .B(n_361), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_408), .B(n_361), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_407), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_407), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_436), .B(n_416), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_442), .B(n_416), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_429), .B(n_416), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_439), .Y(n_475) );
NAND2xp33_ASAP7_75t_SL g476 ( .A(n_430), .B(n_392), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_442), .B(n_407), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
NAND3xp33_ASAP7_75t_SL g479 ( .A(n_461), .B(n_405), .C(n_409), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_449), .B(n_18), .Y(n_481) );
NAND2xp33_ASAP7_75t_SL g482 ( .A(n_430), .B(n_377), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_432), .Y(n_483) );
NAND2x1_ASAP7_75t_L g484 ( .A(n_430), .B(n_415), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_445), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_427), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_428), .Y(n_487) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_435), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_428), .B(n_414), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_454), .B(n_412), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_462), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_455), .B(n_415), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_441), .B(n_415), .Y(n_493) );
NAND2xp33_ASAP7_75t_R g494 ( .A(n_443), .B(n_415), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_456), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_449), .B(n_21), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_464), .B(n_315), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_446), .B(n_315), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_456), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_447), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_466), .B(n_22), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_427), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_450), .B(n_23), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_433), .Y(n_504) );
INVx5_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_433), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_444), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_449), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_467), .B(n_24), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_444), .B(n_29), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_426), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_467), .B(n_30), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_448), .Y(n_513) );
NAND4xp25_ASAP7_75t_SL g514 ( .A(n_440), .B(n_361), .C(n_32), .D(n_33), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_448), .Y(n_515) );
INVx3_ASAP7_75t_L g516 ( .A(n_437), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_457), .B(n_31), .Y(n_517) );
OAI21xp5_ASAP7_75t_SL g518 ( .A1(n_438), .A2(n_468), .B(n_443), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_471), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_458), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_458), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_457), .B(n_34), .Y(n_522) );
INVx4_ASAP7_75t_L g523 ( .A(n_437), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_462), .B(n_39), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_459), .B(n_42), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_424), .B(n_361), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_424), .B(n_49), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_470), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_489), .A2(n_452), .B1(n_425), .B2(n_469), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_489), .A2(n_443), .B1(n_437), .B2(n_434), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_483), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_473), .B(n_434), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_475), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_480), .Y(n_534) );
INVx3_ASAP7_75t_L g535 ( .A(n_523), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_485), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g537 ( .A1(n_524), .A2(n_470), .B(n_465), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_495), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_506), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_499), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_507), .B(n_465), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_478), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_506), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_478), .Y(n_544) );
NOR2xp67_ASAP7_75t_L g545 ( .A(n_505), .B(n_437), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_520), .B(n_463), .Y(n_546) );
NAND2xp33_ASAP7_75t_L g547 ( .A(n_487), .B(n_459), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_511), .Y(n_548) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_523), .B(n_463), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_488), .B(n_460), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_500), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_505), .B(n_453), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_508), .B(n_460), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_518), .A2(n_451), .B1(n_264), .B2(n_232), .Y(n_554) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_476), .A2(n_180), .B1(n_191), .B2(n_197), .C(n_175), .Y(n_555) );
OAI31xp33_ASAP7_75t_L g556 ( .A1(n_476), .A2(n_234), .A3(n_180), .B(n_213), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_488), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_521), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_513), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_515), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_477), .B(n_51), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_528), .B(n_203), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_474), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_486), .Y(n_564) );
INVxp33_ASAP7_75t_L g565 ( .A(n_509), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_486), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_502), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_491), .B(n_203), .Y(n_568) );
AOI32xp33_ASAP7_75t_L g569 ( .A1(n_482), .A2(n_55), .A3(n_57), .B1(n_58), .B2(n_61), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_505), .A2(n_264), .B1(n_232), .B2(n_70), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_472), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_491), .B(n_202), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_505), .B(n_264), .Y(n_573) );
NAND2xp33_ASAP7_75t_L g574 ( .A(n_482), .B(n_264), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_517), .B(n_64), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_502), .Y(n_576) );
AOI311xp33_ASAP7_75t_L g577 ( .A1(n_490), .A2(n_66), .A3(n_215), .B(n_178), .C(n_214), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_504), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_172), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_531), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_542), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_544), .Y(n_582) );
INVx3_ASAP7_75t_L g583 ( .A(n_535), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_558), .B(n_519), .Y(n_584) );
XOR2x2_ASAP7_75t_L g585 ( .A(n_545), .B(n_481), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_550), .B(n_516), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_551), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_532), .B(n_519), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_548), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_571), .B(n_493), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_535), .B(n_516), .Y(n_591) );
NAND2xp33_ASAP7_75t_SL g592 ( .A(n_565), .B(n_494), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_536), .B(n_479), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_559), .B(n_504), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_557), .B(n_526), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_553), .B(n_527), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_547), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_533), .Y(n_598) );
A2O1A1O1Ixp25_ASAP7_75t_L g599 ( .A1(n_537), .A2(n_514), .B(n_479), .C(n_494), .D(n_496), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_534), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_538), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_540), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_563), .B(n_484), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_546), .B(n_522), .Y(n_604) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_574), .B(n_496), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_560), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_550), .Y(n_607) );
OAI211xp5_ASAP7_75t_L g608 ( .A1(n_569), .A2(n_510), .B(n_512), .C(n_525), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_552), .A2(n_481), .B(n_503), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_546), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_529), .A2(n_501), .B(n_498), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_541), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_541), .B(n_497), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_539), .B(n_197), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_543), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_610), .B(n_566), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g617 ( .A1(n_608), .A2(n_537), .B(n_570), .C(n_556), .Y(n_617) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_608), .A2(n_530), .B(n_554), .C(n_577), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_615), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_584), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_590), .B(n_607), .Y(n_621) );
AOI322xp5_ASAP7_75t_L g622 ( .A1(n_593), .A2(n_549), .A3(n_575), .B1(n_576), .B2(n_564), .C1(n_568), .C2(n_572), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_612), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_593), .A2(n_572), .B1(n_568), .B2(n_570), .C(n_578), .Y(n_624) );
XOR2x2_ASAP7_75t_L g625 ( .A(n_585), .B(n_597), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_580), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_588), .B(n_567), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_585), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_587), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_581), .B(n_579), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_598), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_611), .A2(n_561), .B1(n_562), .B2(n_573), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_599), .A2(n_562), .B(n_555), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_591), .A2(n_232), .B(n_202), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_592), .A2(n_178), .B1(n_214), .B2(n_215), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_600), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_582), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_631), .Y(n_638) );
CKINVDCx6p67_ASAP7_75t_R g639 ( .A(n_628), .Y(n_639) );
OAI22xp5_ASAP7_75t_SL g640 ( .A1(n_625), .A2(n_605), .B1(n_583), .B2(n_609), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_627), .B(n_621), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_620), .B(n_586), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_625), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_616), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_618), .A2(n_591), .B(n_592), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_617), .A2(n_596), .B1(n_603), .B2(n_586), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_637), .B(n_603), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_633), .A2(n_586), .B1(n_613), .B2(n_589), .Y(n_648) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_630), .B(n_595), .Y(n_649) );
NAND3xp33_ASAP7_75t_SL g650 ( .A(n_622), .B(n_604), .C(n_594), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_632), .A2(n_624), .B1(n_637), .B2(n_635), .C(n_623), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_626), .A2(n_602), .B(n_601), .C(n_606), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_629), .B(n_583), .C(n_614), .Y(n_653) );
OAI22x1_ASAP7_75t_L g654 ( .A1(n_636), .A2(n_205), .B1(n_178), .B2(n_214), .Y(n_654) );
NAND5xp2_ASAP7_75t_L g655 ( .A(n_634), .B(n_178), .C(n_214), .D(n_215), .E(n_619), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_619), .A2(n_215), .B1(n_628), .B2(n_625), .Y(n_656) );
NOR3xp33_ASAP7_75t_SL g657 ( .A(n_640), .B(n_645), .C(n_651), .Y(n_657) );
NAND2x1_ASAP7_75t_SL g658 ( .A(n_656), .B(n_646), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_643), .B(n_639), .Y(n_659) );
INVx5_ASAP7_75t_L g660 ( .A(n_641), .Y(n_660) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_659), .B(n_645), .C(n_648), .D(n_639), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_660), .Y(n_662) );
OA22x2_ASAP7_75t_L g663 ( .A1(n_657), .A2(n_647), .B1(n_644), .B2(n_649), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_662), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_661), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_664), .B(n_665), .Y(n_666) );
AOI322xp5_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_663), .A3(n_650), .B1(n_647), .B2(n_658), .C1(n_653), .C2(n_642), .Y(n_667) );
AOI221xp5_ASAP7_75t_SL g668 ( .A1(n_667), .A2(n_652), .B1(n_655), .B2(n_654), .C(n_638), .Y(n_668) );
endmodule