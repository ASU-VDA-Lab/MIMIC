module fake_ibex_630_n_963 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_963);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_963;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_510;
wire n_418;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_317;
wire n_375;
wire n_340;
wire n_280;
wire n_708;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_899;
wire n_843;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_874;
wire n_890;
wire n_921;
wire n_912;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_298;
wire n_202;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g197 ( 
.A(n_92),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_65),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_111),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_L g205 ( 
.A(n_68),
.B(n_23),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_159),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_90),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_18),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_18),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_1),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_15),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_79),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_84),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_55),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_114),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_88),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_50),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_59),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_75),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_83),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_154),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_91),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_138),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_93),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_177),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_3),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_171),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_53),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_66),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_33),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_30),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_28),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_179),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_74),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_46),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_112),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_70),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_97),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_141),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_4),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_94),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_99),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_6),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_166),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_6),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_109),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_85),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_186),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_170),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_62),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_125),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_121),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_72),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_40),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_86),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_139),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_51),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_156),
.B(n_22),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_17),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_95),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_67),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_47),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_49),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_103),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_80),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_8),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_165),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_168),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_96),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_21),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_189),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_122),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_157),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_115),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_117),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_158),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_19),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_35),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_11),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_100),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_116),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_110),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_135),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_173),
.B(n_63),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g294 ( 
.A(n_118),
.B(n_131),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_183),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_196),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_160),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_17),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_43),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_36),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_82),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_123),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_19),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_107),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_137),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_29),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_133),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_126),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_71),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_188),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_56),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_32),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_180),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_30),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_41),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_12),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_52),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_181),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_28),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_113),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_81),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_193),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_98),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_237),
.B(n_0),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_1),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_240),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_208),
.B(n_2),
.Y(n_327)
);

OA21x2_ASAP7_75t_L g328 ( 
.A1(n_215),
.A2(n_104),
.B(n_191),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_232),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_238),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_212),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_212),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_223),
.A2(n_102),
.B(n_190),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_212),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_215),
.A2(n_246),
.B(n_245),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_208),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_224),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_238),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_229),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_223),
.B(n_5),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_7),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_235),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_307),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_307),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_245),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_209),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_209),
.B(n_9),
.Y(n_348)
);

OAI21x1_ASAP7_75t_L g349 ( 
.A1(n_246),
.A2(n_105),
.B(n_187),
.Y(n_349)
);

BUFx8_ASAP7_75t_SL g350 ( 
.A(n_232),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_206),
.B(n_9),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_240),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_249),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_262),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_213),
.Y(n_355)
);

OA21x2_ASAP7_75t_L g356 ( 
.A1(n_249),
.A2(n_108),
.B(n_185),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_213),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_282),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_210),
.Y(n_359)
);

OAI22x1_ASAP7_75t_R g360 ( 
.A1(n_312),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_235),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_258),
.B(n_13),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_251),
.B(n_14),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_251),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_253),
.B(n_15),
.Y(n_365)
);

INVx6_ASAP7_75t_L g366 ( 
.A(n_262),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_282),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_308),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_247),
.Y(n_369)
);

AND2x2_ASAP7_75t_SL g370 ( 
.A(n_276),
.B(n_284),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_323),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_197),
.B(n_16),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_262),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_312),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_211),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_241),
.B(n_24),
.Y(n_376)
);

OAI22x1_ASAP7_75t_R g377 ( 
.A1(n_201),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_377)
);

AND2x6_ASAP7_75t_L g378 ( 
.A(n_239),
.B(n_44),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_241),
.B(n_25),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_235),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_263),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_308),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_263),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_279),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_225),
.B(n_26),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_268),
.B(n_300),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_235),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_281),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_268),
.Y(n_390)
);

BUFx8_ASAP7_75t_L g391 ( 
.A(n_317),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_300),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_248),
.B(n_27),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_314),
.B(n_27),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_198),
.A2(n_119),
.B(n_184),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_275),
.B(n_29),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_366),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_370),
.A2(n_302),
.B1(n_204),
.B2(n_219),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

NAND3xp33_ASAP7_75t_L g407 ( 
.A(n_338),
.B(n_298),
.C(n_287),
.Y(n_407)
);

OAI22x1_ASAP7_75t_L g408 ( 
.A1(n_326),
.A2(n_315),
.B1(n_319),
.B2(n_303),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_341),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_341),
.B(n_199),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_336),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_354),
.B(n_271),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_341),
.B(n_200),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_R g416 ( 
.A(n_371),
.B(n_271),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_342),
.B(n_203),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_359),
.B(n_201),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_359),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_354),
.B(n_214),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_376),
.B(n_204),
.Y(n_422)
);

BUFx10_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_378),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_366),
.B(n_214),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_376),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_335),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_340),
.B(n_316),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_331),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_379),
.Y(n_432)
);

OR2x6_ASAP7_75t_L g433 ( 
.A(n_329),
.B(n_288),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_335),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_370),
.B(n_255),
.Y(n_435)
);

NOR3xp33_ASAP7_75t_L g436 ( 
.A(n_374),
.B(n_306),
.C(n_264),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_335),
.Y(n_437)
);

OA22x2_ASAP7_75t_L g438 ( 
.A1(n_386),
.A2(n_255),
.B1(n_299),
.B2(n_304),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_348),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_348),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_384),
.B(n_304),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_373),
.B(n_216),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_380),
.Y(n_443)
);

BUFx6f_ASAP7_75t_SL g444 ( 
.A(n_363),
.Y(n_444)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_391),
.B(n_218),
.C(n_217),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_365),
.Y(n_447)
);

OAI22x1_ASAP7_75t_L g448 ( 
.A1(n_360),
.A2(n_274),
.B1(n_321),
.B2(n_318),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_365),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_333),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_333),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_373),
.B(n_220),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_344),
.B(n_222),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_350),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_330),
.B(n_202),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_339),
.B(n_231),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_339),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_337),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_391),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_386),
.B(n_205),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_378),
.A2(n_322),
.B1(n_233),
.B2(n_234),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_324),
.A2(n_243),
.B1(n_242),
.B2(n_313),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_391),
.B(n_221),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_344),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_351),
.B(n_320),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_328),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_345),
.B(n_236),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_362),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_324),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_372),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_345),
.B(n_226),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_325),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_364),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_328),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_346),
.B(n_227),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_347),
.B(n_244),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_328),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_353),
.B(n_250),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_353),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_355),
.B(n_252),
.Y(n_483)
);

AO21x2_ASAP7_75t_L g484 ( 
.A1(n_349),
.A2(n_207),
.B(n_254),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_364),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_463),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_427),
.B(n_325),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_402),
.B(n_398),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_403),
.B(n_385),
.Y(n_489)
);

BUFx8_ASAP7_75t_L g490 ( 
.A(n_455),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_476),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_393),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_438),
.A2(n_358),
.B1(n_367),
.B2(n_368),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_463),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_404),
.B(n_410),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_485),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_357),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_432),
.B(n_459),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_425),
.B(n_228),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_425),
.B(n_256),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_444),
.A2(n_242),
.B1(n_243),
.B2(n_352),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_432),
.B(n_381),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_404),
.B(n_410),
.Y(n_503)
);

NOR3xp33_ASAP7_75t_L g504 ( 
.A(n_422),
.B(n_375),
.C(n_392),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_420),
.B(n_383),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_444),
.A2(n_367),
.B1(n_358),
.B2(n_368),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_390),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_406),
.B(n_382),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_419),
.B(n_392),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_460),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_438),
.A2(n_382),
.B1(n_388),
.B2(n_395),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_467),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_414),
.B(n_392),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_441),
.B(n_473),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_423),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_472),
.Y(n_516)
);

O2A1O1Ixp5_ASAP7_75t_L g517 ( 
.A1(n_469),
.A2(n_283),
.B(n_257),
.C(n_259),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_482),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_409),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_424),
.B(n_388),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_473),
.B(n_397),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_450),
.B(n_334),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_426),
.B(n_230),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_400),
.B(n_356),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_439),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_465),
.B(n_31),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_458),
.B(n_265),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_L g529 ( 
.A1(n_440),
.A2(n_396),
.B(n_260),
.C(n_261),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_450),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_L g531 ( 
.A1(n_447),
.A2(n_291),
.B(n_266),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_449),
.A2(n_296),
.B1(n_301),
.B2(n_269),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_442),
.B(n_270),
.Y(n_533)
);

AOI221xp5_ASAP7_75t_L g534 ( 
.A1(n_408),
.A2(n_310),
.B1(n_309),
.B2(n_292),
.C(n_277),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_422),
.Y(n_535)
);

NOR3xp33_ASAP7_75t_L g536 ( 
.A(n_436),
.B(n_377),
.C(n_267),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_456),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_412),
.B(n_278),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g539 ( 
.A1(n_405),
.A2(n_239),
.B1(n_272),
.B2(n_273),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_435),
.A2(n_311),
.B1(n_295),
.B2(n_280),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_415),
.B(n_289),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_445),
.B(n_290),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_475),
.B(n_31),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_411),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_417),
.B(n_305),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_466),
.B(n_293),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_416),
.B(n_272),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_431),
.B(n_273),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_413),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_453),
.A2(n_285),
.B1(n_294),
.B2(n_281),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_448),
.B(n_32),
.Y(n_551)
);

NAND2x1_ASAP7_75t_L g552 ( 
.A(n_464),
.B(n_281),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_413),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_464),
.B(n_285),
.Y(n_554)
);

AOI221xp5_ASAP7_75t_L g555 ( 
.A1(n_430),
.A2(n_297),
.B1(n_387),
.B2(n_361),
.C(n_343),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_484),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_462),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_484),
.Y(n_558)
);

O2A1O1Ixp33_ASAP7_75t_L g559 ( 
.A1(n_430),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_407),
.B(n_297),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_462),
.B(n_297),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_483),
.B(n_343),
.Y(n_562)
);

INVxp33_ASAP7_75t_L g563 ( 
.A(n_479),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_478),
.A2(n_389),
.B1(n_387),
.B2(n_361),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_474),
.B(n_343),
.Y(n_565)
);

NOR3xp33_ASAP7_75t_L g566 ( 
.A(n_468),
.B(n_36),
.C(n_37),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_514),
.B(n_433),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_487),
.B(n_479),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_556),
.A2(n_469),
.B(n_480),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_497),
.B(n_477),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_558),
.A2(n_480),
.B(n_477),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_495),
.Y(n_572)
);

OAI22xp33_ASAP7_75t_L g573 ( 
.A1(n_501),
.A2(n_433),
.B1(n_470),
.B2(n_454),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_487),
.A2(n_433),
.B1(n_483),
.B2(n_481),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_530),
.B(n_481),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_497),
.B(n_454),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_496),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_516),
.B(n_470),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_492),
.B(n_37),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_544),
.A2(n_553),
.B(n_549),
.Y(n_580)
);

CKINVDCx10_ASAP7_75t_R g581 ( 
.A(n_490),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_488),
.B(n_38),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_488),
.B(n_489),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_515),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_524),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_503),
.B(n_38),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_535),
.A2(n_361),
.B1(n_387),
.B2(n_389),
.Y(n_587)
);

AOI21xp33_ASAP7_75t_L g588 ( 
.A1(n_563),
.A2(n_39),
.B(n_40),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_486),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_507),
.B(n_39),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_496),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_517),
.A2(n_529),
.B(n_525),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_509),
.B(n_41),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_498),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_521),
.B(n_42),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g596 ( 
.A1(n_527),
.A2(n_42),
.B(n_434),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_502),
.B(n_45),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_493),
.A2(n_434),
.B1(n_421),
.B2(n_446),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_510),
.Y(n_599)
);

AO22x1_ASAP7_75t_L g600 ( 
.A1(n_490),
.A2(n_48),
.B1(n_54),
.B2(n_57),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_498),
.B(n_58),
.Y(n_601)
);

CKINVDCx8_ASAP7_75t_R g602 ( 
.A(n_502),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_522),
.A2(n_451),
.B(n_437),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_540),
.B(n_60),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_543),
.B(n_61),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_519),
.A2(n_429),
.B1(n_446),
.B2(n_443),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_508),
.A2(n_520),
.B(n_565),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_508),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_505),
.A2(n_428),
.B(n_401),
.C(n_452),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_511),
.B(n_428),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_L g611 ( 
.A(n_536),
.B(n_64),
.C(n_69),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_520),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_526),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_537),
.Y(n_614)
);

NOR3xp33_ASAP7_75t_L g615 ( 
.A(n_539),
.B(n_73),
.C(n_76),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_504),
.A2(n_401),
.B1(n_452),
.B2(n_87),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_557),
.A2(n_452),
.B1(n_78),
.B2(n_89),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_524),
.B(n_77),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_532),
.B(n_106),
.Y(n_619)
);

NAND3xp33_ASAP7_75t_L g620 ( 
.A(n_566),
.B(n_534),
.C(n_561),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_528),
.B(n_192),
.Y(n_621)
);

O2A1O1Ixp33_ASAP7_75t_SL g622 ( 
.A1(n_552),
.A2(n_120),
.B(n_124),
.C(n_127),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_513),
.B(n_182),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_518),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_554),
.A2(n_132),
.B(n_134),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_506),
.B(n_136),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_547),
.B(n_140),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_494),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_538),
.B(n_142),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_512),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_SL g631 ( 
.A1(n_542),
.A2(n_143),
.B(n_144),
.C(n_147),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_541),
.B(n_148),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_541),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_533),
.B(n_523),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_551),
.B(n_162),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_559),
.B(n_163),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_545),
.B(n_175),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_562),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_491),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_583),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_634),
.A2(n_560),
.B(n_550),
.C(n_548),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_602),
.B(n_531),
.Y(n_642)
);

BUFx4f_ASAP7_75t_L g643 ( 
.A(n_601),
.Y(n_643)
);

BUFx5_ASAP7_75t_L g644 ( 
.A(n_618),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_599),
.Y(n_645)
);

AOI221x1_ASAP7_75t_L g646 ( 
.A1(n_592),
.A2(n_562),
.B1(n_546),
.B2(n_555),
.C(n_564),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_568),
.B(n_562),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_601),
.B(n_499),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_596),
.A2(n_500),
.B(n_167),
.C(n_169),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_630),
.Y(n_650)
);

CKINVDCx11_ASAP7_75t_R g651 ( 
.A(n_581),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_572),
.B(n_584),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_607),
.A2(n_603),
.B(n_620),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_594),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_585),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_586),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_574),
.B(n_613),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_614),
.B(n_573),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_584),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_620),
.A2(n_575),
.B(n_570),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_567),
.B(n_593),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_596),
.A2(n_629),
.B(n_632),
.C(n_582),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_576),
.B(n_628),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_578),
.B(n_579),
.Y(n_664)
);

NOR2xp67_ASAP7_75t_L g665 ( 
.A(n_604),
.B(n_597),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_636),
.B(n_605),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_589),
.Y(n_667)
);

BUFx5_ASAP7_75t_L g668 ( 
.A(n_618),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_577),
.Y(n_669)
);

OAI22x1_ASAP7_75t_L g670 ( 
.A1(n_595),
.A2(n_590),
.B1(n_600),
.B2(n_616),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_621),
.A2(n_615),
.B(n_637),
.C(n_619),
.Y(n_671)
);

AOI211x1_ASAP7_75t_L g672 ( 
.A1(n_588),
.A2(n_610),
.B(n_624),
.C(n_627),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_585),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_636),
.B(n_591),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_591),
.B(n_638),
.Y(n_675)
);

BUFx4f_ASAP7_75t_L g676 ( 
.A(n_636),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_639),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_611),
.B(n_633),
.C(n_625),
.Y(n_678)
);

BUFx4_ASAP7_75t_R g679 ( 
.A(n_635),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_626),
.B(n_623),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_598),
.Y(n_681)
);

AO21x2_ASAP7_75t_L g682 ( 
.A1(n_617),
.A2(n_622),
.B(n_631),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_585),
.B(n_606),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_587),
.B(n_583),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_583),
.B(n_608),
.Y(n_685)
);

AND2x2_ASAP7_75t_SL g686 ( 
.A(n_601),
.B(n_418),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_583),
.B(n_608),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_583),
.B(n_608),
.Y(n_688)
);

INVx5_ASAP7_75t_L g689 ( 
.A(n_584),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_583),
.B(n_608),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_584),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_583),
.B(n_608),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_599),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_596),
.A2(n_573),
.B1(n_567),
.B2(n_574),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_583),
.B(n_608),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_569),
.A2(n_571),
.B(n_580),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_599),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_583),
.B(n_601),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_569),
.A2(n_571),
.B(n_580),
.Y(n_699)
);

INVx5_ASAP7_75t_L g700 ( 
.A(n_584),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_583),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_583),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_583),
.B(n_495),
.Y(n_703)
);

AO31x2_ASAP7_75t_L g704 ( 
.A1(n_609),
.A2(n_529),
.A3(n_558),
.B(n_556),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_583),
.B(n_608),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_569),
.A2(n_571),
.B(n_580),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_583),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_583),
.A2(n_634),
.B(n_596),
.C(n_620),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_585),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_596),
.A2(n_573),
.B1(n_567),
.B2(n_574),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_583),
.B(n_608),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_583),
.A2(n_612),
.B1(n_608),
.B2(n_601),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_583),
.B(n_608),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_583),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_583),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_583),
.B(n_419),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_638),
.Y(n_717)
);

AO31x2_ASAP7_75t_L g718 ( 
.A1(n_609),
.A2(n_529),
.A3(n_558),
.B(n_556),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_640),
.B(n_714),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_SL g720 ( 
.A(n_676),
.B(n_643),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_685),
.B(n_687),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_707),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_712),
.A2(n_698),
.B1(n_694),
.B2(n_710),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_701),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_701),
.Y(n_725)
);

INVx8_ASAP7_75t_L g726 ( 
.A(n_689),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_702),
.B(n_715),
.Y(n_727)
);

AO31x2_ASAP7_75t_L g728 ( 
.A1(n_681),
.A2(n_670),
.A3(n_662),
.B(n_708),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_660),
.A2(n_657),
.B(n_678),
.Y(n_729)
);

AO31x2_ASAP7_75t_L g730 ( 
.A1(n_696),
.A2(n_706),
.A3(n_699),
.B(n_671),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_702),
.Y(n_731)
);

AO31x2_ASAP7_75t_L g732 ( 
.A1(n_646),
.A2(n_641),
.A3(n_680),
.B(n_683),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_715),
.B(n_686),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_688),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_690),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_716),
.B(n_703),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_689),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_692),
.Y(n_738)
);

BUFx2_ASAP7_75t_R g739 ( 
.A(n_651),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_689),
.Y(n_740)
);

AO21x2_ASAP7_75t_L g741 ( 
.A1(n_682),
.A2(n_678),
.B(n_694),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_691),
.Y(n_742)
);

NAND2x1p5_ASAP7_75t_L g743 ( 
.A(n_643),
.B(n_691),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_695),
.B(n_705),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_711),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_691),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_655),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_698),
.A2(n_713),
.B(n_664),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_700),
.Y(n_749)
);

OAI21x1_ASAP7_75t_SL g750 ( 
.A1(n_674),
.A2(n_710),
.B(n_649),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_645),
.Y(n_751)
);

OA21x2_ASAP7_75t_L g752 ( 
.A1(n_658),
.A2(n_647),
.B(n_684),
.Y(n_752)
);

AOI22x1_ASAP7_75t_L g753 ( 
.A1(n_656),
.A2(n_666),
.B1(n_648),
.B2(n_717),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_700),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_661),
.A2(n_665),
.B1(n_672),
.B2(n_650),
.Y(n_755)
);

CKINVDCx6p67_ASAP7_75t_R g756 ( 
.A(n_700),
.Y(n_756)
);

AO21x2_ASAP7_75t_L g757 ( 
.A1(n_682),
.A2(n_665),
.B(n_675),
.Y(n_757)
);

OAI21xp33_ASAP7_75t_SL g758 ( 
.A1(n_679),
.A2(n_697),
.B(n_693),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_667),
.Y(n_759)
);

BUFx10_ASAP7_75t_L g760 ( 
.A(n_659),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_648),
.B(n_669),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_654),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_655),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_673),
.A2(n_709),
.B(n_642),
.Y(n_764)
);

OA21x2_ASAP7_75t_L g765 ( 
.A1(n_704),
.A2(n_718),
.B(n_672),
.Y(n_765)
);

AO31x2_ASAP7_75t_L g766 ( 
.A1(n_718),
.A2(n_644),
.A3(n_668),
.B(n_673),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_677),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_644),
.A2(n_668),
.B(n_652),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_663),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_640),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_640),
.Y(n_771)
);

AO31x2_ASAP7_75t_L g772 ( 
.A1(n_681),
.A2(n_670),
.A3(n_529),
.B(n_662),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_689),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_640),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_655),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_708),
.A2(n_653),
.B(n_662),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_640),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_640),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_643),
.B(n_689),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_707),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_701),
.B(n_702),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_655),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_640),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_708),
.A2(n_653),
.B(n_662),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_640),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_640),
.B(n_714),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_727),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_747),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_745),
.B(n_738),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_727),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_721),
.B(n_744),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_730),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_745),
.B(n_734),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_726),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_721),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_724),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_721),
.B(n_744),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_733),
.B(n_719),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_744),
.B(n_781),
.Y(n_799)
);

AO21x1_ASAP7_75t_SL g800 ( 
.A1(n_723),
.A2(n_784),
.B(n_776),
.Y(n_800)
);

CKINVDCx11_ASAP7_75t_R g801 ( 
.A(n_749),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_735),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_725),
.Y(n_803)
);

INVxp33_ASAP7_75t_L g804 ( 
.A(n_777),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_726),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_731),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_781),
.B(n_736),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_780),
.B(n_722),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_723),
.B(n_786),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_752),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_748),
.B(n_759),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_770),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_752),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_771),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_748),
.B(n_751),
.Y(n_815)
);

INVxp33_ASAP7_75t_L g816 ( 
.A(n_743),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_774),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_768),
.B(n_766),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_784),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_726),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_728),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_772),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_729),
.B(n_765),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_729),
.B(n_765),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_758),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_772),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_766),
.B(n_757),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_755),
.B(n_769),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_778),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_772),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_747),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_720),
.B(n_758),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_783),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_732),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_815),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_800),
.B(n_741),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_815),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_800),
.B(n_811),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_805),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_810),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_809),
.A2(n_720),
.B1(n_797),
.B2(n_802),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_813),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_787),
.B(n_785),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_801),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_819),
.B(n_823),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_805),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_823),
.B(n_762),
.Y(n_847)
);

OAI221xp5_ASAP7_75t_L g848 ( 
.A1(n_798),
.A2(n_761),
.B1(n_753),
.B2(n_779),
.C(n_767),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_818),
.B(n_764),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_824),
.B(n_742),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_824),
.B(n_742),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_796),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_828),
.B(n_773),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_796),
.B(n_746),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_791),
.A2(n_756),
.B1(n_737),
.B2(n_740),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_804),
.B(n_739),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_805),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_787),
.B(n_761),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_818),
.B(n_764),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_790),
.B(n_767),
.Y(n_860)
);

OR2x6_ASAP7_75t_L g861 ( 
.A(n_825),
.B(n_832),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_789),
.B(n_803),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_803),
.B(n_806),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_797),
.A2(n_750),
.B1(n_737),
.B2(n_754),
.Y(n_864)
);

AND2x4_ASAP7_75t_SL g865 ( 
.A(n_799),
.B(n_795),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_808),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_SL g867 ( 
.A1(n_799),
.A2(n_760),
.B1(n_763),
.B2(n_775),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_840),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_849),
.B(n_827),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_839),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_835),
.B(n_837),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_845),
.B(n_821),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_839),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_845),
.B(n_834),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_838),
.B(n_792),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_838),
.B(n_792),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_850),
.B(n_826),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_842),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_862),
.B(n_830),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_850),
.B(n_822),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_851),
.B(n_822),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_856),
.B(n_739),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_868),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_868),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_874),
.B(n_862),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_874),
.B(n_836),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_874),
.B(n_836),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_877),
.B(n_851),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_872),
.B(n_866),
.Y(n_889)
);

AOI211xp5_ASAP7_75t_SL g890 ( 
.A1(n_882),
.A2(n_855),
.B(n_848),
.C(n_841),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_871),
.B(n_863),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_L g892 ( 
.A(n_878),
.B(n_857),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_880),
.B(n_847),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_872),
.B(n_847),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_871),
.B(n_844),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_881),
.B(n_853),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_879),
.B(n_863),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_869),
.B(n_859),
.Y(n_898)
);

NAND2x1_ASAP7_75t_L g899 ( 
.A(n_869),
.B(n_861),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_885),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_885),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_889),
.B(n_879),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_898),
.B(n_869),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_886),
.B(n_875),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_897),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_897),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_895),
.A2(n_841),
.B1(n_875),
.B2(n_876),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_891),
.Y(n_908)
);

INVx3_ASAP7_75t_SL g909 ( 
.A(n_891),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_883),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_884),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_888),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_886),
.B(n_875),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_908),
.A2(n_896),
.B1(n_888),
.B2(n_893),
.C(n_894),
.Y(n_914)
);

O2A1O1Ixp5_ASAP7_75t_L g915 ( 
.A1(n_903),
.A2(n_890),
.B(n_899),
.C(n_846),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_900),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_901),
.Y(n_917)
);

OAI21xp33_ASAP7_75t_L g918 ( 
.A1(n_907),
.A2(n_887),
.B(n_896),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_909),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_910),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_911),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_905),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_909),
.A2(n_898),
.B1(n_892),
.B2(n_887),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_906),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_916),
.B(n_902),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_919),
.Y(n_926)
);

OAI211xp5_ASAP7_75t_L g927 ( 
.A1(n_923),
.A2(n_846),
.B(n_899),
.C(n_864),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_914),
.B(n_893),
.Y(n_928)
);

AOI222xp33_ASAP7_75t_L g929 ( 
.A1(n_928),
.A2(n_918),
.B1(n_922),
.B2(n_924),
.C1(n_917),
.C2(n_921),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_927),
.A2(n_915),
.B(n_892),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_925),
.Y(n_931)
);

OAI21xp33_ASAP7_75t_L g932 ( 
.A1(n_929),
.A2(n_926),
.B(n_920),
.Y(n_932)
);

AOI211x1_ASAP7_75t_SL g933 ( 
.A1(n_930),
.A2(n_920),
.B(n_843),
.C(n_858),
.Y(n_933)
);

NOR4xp75_ASAP7_75t_L g934 ( 
.A(n_932),
.B(n_915),
.C(n_820),
.D(n_794),
.Y(n_934)
);

NOR2x1_ASAP7_75t_L g935 ( 
.A(n_933),
.B(n_846),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_934),
.B(n_931),
.C(n_793),
.Y(n_936)
);

OAI322xp33_ASAP7_75t_L g937 ( 
.A1(n_935),
.A2(n_912),
.A3(n_829),
.B1(n_833),
.B2(n_814),
.C1(n_812),
.C2(n_817),
.Y(n_937)
);

XNOR2xp5_ASAP7_75t_L g938 ( 
.A(n_936),
.B(n_816),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_937),
.B(n_904),
.Y(n_939)
);

AND2x2_ASAP7_75t_SL g940 ( 
.A(n_939),
.B(n_846),
.Y(n_940)
);

XOR2xp5_ASAP7_75t_L g941 ( 
.A(n_938),
.B(n_794),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_938),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_941),
.A2(n_820),
.B1(n_857),
.B2(n_867),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_942),
.A2(n_839),
.B1(n_903),
.B2(n_873),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_940),
.A2(n_860),
.B(n_807),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_942),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_940),
.B(n_852),
.Y(n_947)
);

AO21x2_ASAP7_75t_L g948 ( 
.A1(n_946),
.A2(n_806),
.B(n_808),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_944),
.B(n_904),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_943),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_947),
.A2(n_903),
.B1(n_873),
.B2(n_870),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_945),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_L g953 ( 
.A(n_946),
.B(n_775),
.C(n_782),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_946),
.B(n_870),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_954),
.A2(n_913),
.B1(n_873),
.B2(n_870),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_950),
.A2(n_913),
.B1(n_854),
.B2(n_898),
.Y(n_956)
);

INVxp33_ASAP7_75t_L g957 ( 
.A(n_953),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_948),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_957),
.A2(n_952),
.B(n_949),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_958),
.B(n_951),
.Y(n_960)
);

AOI22x1_ASAP7_75t_L g961 ( 
.A1(n_956),
.A2(n_854),
.B1(n_831),
.B2(n_788),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_959),
.B(n_955),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_962),
.A2(n_960),
.B1(n_961),
.B2(n_865),
.Y(n_963)
);


endmodule