module fake_jpeg_28293_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_9),
.B(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_17),
.B1(n_23),
.B2(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_56),
.B1(n_25),
.B2(n_23),
.Y(n_83)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_30),
.B1(n_26),
.B2(n_19),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_25),
.B1(n_27),
.B2(n_22),
.Y(n_85)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_59),
.Y(n_88)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_17),
.B1(n_23),
.B2(n_32),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_26),
.B1(n_19),
.B2(n_31),
.Y(n_57)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_73)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_40),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_24),
.B(n_17),
.C(n_28),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_72),
.B(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_30),
.B(n_43),
.C(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_94),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_40),
.C(n_43),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_60),
.C(n_48),
.Y(n_103)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

OAI22x1_ASAP7_75t_R g78 ( 
.A1(n_57),
.A2(n_52),
.B1(n_61),
.B2(n_65),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_78),
.A2(n_92),
.B1(n_34),
.B2(n_20),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_30),
.B(n_41),
.C(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_84),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_31),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_16),
.B1(n_28),
.B2(n_32),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_45),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_64),
.B1(n_58),
.B2(n_55),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_16),
.B1(n_31),
.B2(n_28),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_42),
.B1(n_34),
.B2(n_21),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_45),
.B1(n_66),
.B2(n_62),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_16),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_33),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_107),
.B1(n_111),
.B2(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_50),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_66),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_51),
.B1(n_53),
.B2(n_25),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_122),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_91),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

AO22x2_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_78),
.B1(n_72),
.B2(n_80),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_123),
.A2(n_125),
.B1(n_126),
.B2(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_133),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_78),
.B1(n_88),
.B2(n_72),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_80),
.B1(n_73),
.B2(n_74),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_68),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_22),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_91),
.C(n_69),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_113),
.C(n_101),
.Y(n_155)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_137),
.Y(n_153)
);

FAx1_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_91),
.CI(n_85),
.CON(n_136),
.SN(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_111),
.B(n_122),
.C(n_118),
.D(n_105),
.Y(n_158)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_96),
.B(n_120),
.C(n_116),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_121),
.B(n_108),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_93),
.B1(n_87),
.B2(n_79),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_144),
.B1(n_149),
.B2(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_142),
.Y(n_173)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_79),
.B1(n_77),
.B2(n_81),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_27),
.B1(n_18),
.B2(n_21),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_106),
.A2(n_84),
.B1(n_82),
.B2(n_76),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_152),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_76),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_105),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_92),
.B1(n_25),
.B2(n_33),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_102),
.A2(n_22),
.B1(n_18),
.B2(n_33),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_20),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_110),
.B1(n_99),
.B2(n_119),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_135),
.B(n_99),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_155),
.B(n_161),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_179),
.B(n_8),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_104),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_160),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_165),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_166),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_95),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_95),
.C(n_115),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_130),
.C(n_131),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_12),
.B(n_1),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_8),
.B(n_2),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_143),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_176),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_118),
.C(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_180),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_92),
.B1(n_121),
.B2(n_27),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_181),
.A2(n_185),
.B1(n_127),
.B2(n_34),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_184),
.B1(n_34),
.B2(n_0),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_21),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_132),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_34),
.C(n_21),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_152),
.B1(n_123),
.B2(n_136),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_191),
.B1(n_194),
.B2(n_201),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_123),
.A3(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_123),
.B1(n_150),
.B2(n_127),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_199),
.B1(n_175),
.B2(n_180),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_7),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_200),
.B(n_202),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_158),
.B1(n_179),
.B2(n_163),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_153),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_173),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_8),
.B(n_2),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_157),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_171),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_210),
.B1(n_154),
.B2(n_174),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_170),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_216),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_161),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_214),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_217),
.B(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_159),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_160),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_222),
.A2(n_223),
.B1(n_229),
.B2(n_234),
.Y(n_250)
);

INVxp33_ASAP7_75t_SL g224 ( 
.A(n_193),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_226),
.B(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_197),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_227),
.A2(n_230),
.B(n_233),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_166),
.C(n_165),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_240),
.C(n_4),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_186),
.A2(n_185),
.B1(n_172),
.B2(n_155),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_232),
.A2(n_237),
.B1(n_198),
.B2(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_156),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_236),
.A2(n_194),
.B1(n_212),
.B2(n_187),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_172),
.B1(n_183),
.B2(n_181),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_201),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_6),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_177),
.C(n_164),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_251),
.B1(n_257),
.B2(n_250),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_209),
.B(n_204),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_253),
.B(n_238),
.Y(n_267)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_221),
.B(n_192),
.CI(n_189),
.CON(n_244),
.SN(n_244)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_253),
.B(n_243),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_198),
.B1(n_187),
.B2(n_211),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_245),
.A2(n_252),
.B1(n_11),
.B2(n_12),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_216),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_258),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_234),
.C(n_238),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_232),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_249),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_219),
.A2(n_212),
.B1(n_192),
.B2(n_195),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_200),
.B1(n_202),
.B2(n_207),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_200),
.B(n_210),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_219),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_3),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_261),
.C(n_240),
.Y(n_264)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_256),
.Y(n_262)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_270),
.B1(n_273),
.B2(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_275),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_267),
.B(n_261),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_258),
.B1(n_246),
.B2(n_14),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_237),
.B1(n_220),
.B2(n_223),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_222),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_231),
.Y(n_272)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_7),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_274),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_244),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_265),
.B1(n_277),
.B2(n_276),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_259),
.C(n_242),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_264),
.C(n_269),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_245),
.B(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_242),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_287),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_244),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_11),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_294),
.B(n_303),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_282),
.C(n_293),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_271),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_305),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_281),
.A2(n_275),
.B1(n_278),
.B2(n_274),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_298),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_270),
.B1(n_263),
.B2(n_262),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_13),
.B(n_14),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_304),
.A2(n_290),
.B(n_289),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_13),
.CI(n_14),
.CON(n_305),
.SN(n_305)
);

AOI31xp33_ASAP7_75t_L g306 ( 
.A1(n_280),
.A2(n_13),
.A3(n_15),
.B(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_13),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_279),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_314),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_300),
.B(n_296),
.C(n_302),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_299),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_313),
.B(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_301),
.B(n_285),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_283),
.C(n_288),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_311),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_294),
.B(n_300),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_319),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_321),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_320),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_324),
.B(n_322),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_312),
.Y(n_328)
);

OAI321xp33_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_321),
.A3(n_304),
.B1(n_325),
.B2(n_283),
.C(n_305),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_305),
.B(n_15),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_330),
.Y(n_331)
);


endmodule