module real_jpeg_28386_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_1),
.A2(n_25),
.B1(n_28),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_73),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_25),
.B1(n_28),
.B2(n_73),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_76),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_4),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_85),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_85),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_4),
.A2(n_25),
.B1(n_28),
.B2(n_85),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_7),
.A2(n_25),
.B1(n_28),
.B2(n_39),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_8),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_8),
.A2(n_71),
.B1(n_76),
.B2(n_86),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_71),
.Y(n_177)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_9),
.B(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_9),
.B(n_65),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_9),
.A2(n_65),
.B(n_134),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_78),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_9),
.A2(n_25),
.B(n_29),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_9),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_9),
.A2(n_41),
.B1(n_50),
.B2(n_185),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_105)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_11),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_12),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_12),
.A2(n_25),
.B1(n_28),
.B2(n_56),
.Y(n_131)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_108),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_108),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_87),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_24),
.A2(n_36),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_24),
.A2(n_36),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_24),
.A2(n_36),
.B1(n_141),
.B2(n_160),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_24),
.B(n_78),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_27),
.A2(n_32),
.B(n_78),
.C(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_28),
.B(n_190),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g132 ( 
.A1(n_31),
.A2(n_66),
.A3(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_32),
.B(n_63),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_54),
.B(n_57),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_36),
.A2(n_142),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_47),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_41),
.A2(n_45),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_41),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_41),
.A2(n_177),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_42),
.B(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_42),
.A2(n_48),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_42),
.A2(n_107),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_50),
.A2(n_105),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_50),
.B(n_78),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.C(n_74),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_52),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_55),
.B(n_58),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_61),
.A2(n_69),
.B1(n_70),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_69),
.B1(n_116),
.B2(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_69),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_62)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_66),
.B1(n_80),
.B2(n_81),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_80),
.Y(n_103)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_75),
.B1(n_82),
.B2(n_103),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.CON(n_75),
.SN(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_80),
.B(n_82),
.C(n_83),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_80),
.Y(n_82)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_101),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_104),
.Y(n_113)
);

INVx5_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_131),
.Y(n_172)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_114),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_109),
.A2(n_110),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_114),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.C(n_119),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_201),
.B(n_207),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_153),
.B(n_200),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_143),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_127),
.B(n_143),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_136),
.C(n_139),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_128),
.A2(n_129),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_132),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_150),
.C(n_151),
.Y(n_202)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_194),
.B(n_199),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_173),
.B(n_193),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_156),
.B(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_181),
.B(n_192),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_179),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_187),
.B(n_191),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_184),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_195),
.B(n_196),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_202),
.B(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);


endmodule