module real_jpeg_7018_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_1),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_1),
.Y(n_137)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_1),
.Y(n_146)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_1),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_1),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_1),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_1),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_1),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_2),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_2),
.A2(n_120),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_2),
.A2(n_120),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_2),
.A2(n_67),
.B1(n_120),
.B2(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_3),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_3),
.A2(n_201),
.B1(n_257),
.B2(n_261),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_3),
.B(n_275),
.C(n_279),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_3),
.B(n_105),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_3),
.B(n_171),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_3),
.B(n_56),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_3),
.B(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_6),
.Y(n_171)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_6),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_6),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_6),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_6),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_7),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_7),
.A2(n_63),
.B1(n_70),
.B2(n_112),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_8),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_8),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_8),
.A2(n_51),
.B1(n_86),
.B2(n_231),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_9),
.A2(n_30),
.B1(n_51),
.B2(n_54),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_9),
.A2(n_54),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_9),
.A2(n_54),
.B1(n_356),
.B2(n_360),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_10),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_10),
.Y(n_150)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_10),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_12),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_12),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_12),
.A2(n_63),
.B1(n_133),
.B2(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_12),
.A2(n_133),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_12),
.A2(n_133),
.B1(n_190),
.B2(n_385),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_13),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_13),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_13),
.A2(n_62),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_13),
.A2(n_62),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_14),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_14),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_14),
.A2(n_159),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_14),
.A2(n_159),
.B1(n_286),
.B2(n_290),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_14),
.A2(n_159),
.B1(n_257),
.B2(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_15),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_15),
.Y(n_173)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_247),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_246),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_225),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_21),
.B(n_225),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_164),
.C(n_178),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_22),
.A2(n_23),
.B1(n_164),
.B2(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_91),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_24),
.B(n_92),
.C(n_163),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_65),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_25),
.B(n_65),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_26),
.A2(n_256),
.B(n_263),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_26),
.A2(n_55),
.B1(n_300),
.B2(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_26),
.A2(n_263),
.B(n_338),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_27),
.A2(n_56),
.B1(n_58),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_27),
.A2(n_56),
.B1(n_166),
.B2(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_27),
.B(n_264),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_31),
.Y(n_268)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_31),
.Y(n_302)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_32),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_32),
.Y(n_367)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_34),
.Y(n_278)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_39),
.A2(n_300),
.B(n_303),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_44),
.Y(n_282)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_44),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_45),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_47),
.Y(n_174)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_47),
.Y(n_209)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_50),
.A2(n_55),
.B(n_303),
.Y(n_413)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_53),
.Y(n_262)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_56),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_61),
.Y(n_232)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_73),
.B1(n_80),
.B2(n_89),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_66),
.Y(n_214)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_69),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_72),
.Y(n_311)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_73),
.B(n_295),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_73),
.A2(n_293),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_73),
.A2(n_208),
.B1(n_355),
.B2(n_390),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_76),
.Y(n_391)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_81),
.A2(n_168),
.B1(n_169),
.B2(n_172),
.Y(n_167)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_85),
.Y(n_289)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_87),
.Y(n_317)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_129),
.B1(n_162),
.B2(n_163),
.Y(n_91)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

AOI22x1_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_105),
.B1(n_116),
.B2(n_124),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_93),
.A2(n_216),
.B(n_223),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_93),
.A2(n_223),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_93),
.B(n_116),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_94),
.A2(n_125),
.B1(n_224),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_94),
.A2(n_217),
.B1(n_224),
.B2(n_384),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_105),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_97),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_100),
.Y(n_347)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_101),
.Y(n_219)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_101),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_101),
.Y(n_351)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_102),
.Y(n_373)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_105),
.Y(n_224)
);

AO22x2_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_112),
.B2(n_114),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_111),
.Y(n_341)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_117),
.B(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_118),
.Y(n_243)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_122),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_121),
.Y(n_385)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_123),
.Y(n_242)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_138),
.B1(n_151),
.B2(n_156),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_130),
.A2(n_181),
.B(n_183),
.Y(n_180)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_138),
.A2(n_156),
.B(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_184),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_139),
.A2(n_406),
.B(n_410),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_151),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.B1(n_147),
.B2(n_149),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_151),
.B(n_201),
.Y(n_388)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_164),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_165),
.B(n_167),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_170),
.B1(n_207),
.B2(n_214),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_168),
.A2(n_172),
.B(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_168),
.A2(n_285),
.B(n_292),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_168),
.A2(n_201),
.B(n_292),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_177),
.Y(n_291)
);

INVx8_ASAP7_75t_L g319 ( 
.A(n_177),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_178),
.B(n_428),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.C(n_215),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_179),
.A2(n_180),
.B1(n_215),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_182),
.B(n_184),
.Y(n_245)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_188),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_205),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_189),
.A2(n_205),
.B1(n_206),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_189),
.Y(n_399)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.A3(n_193),
.B1(n_195),
.B2(n_200),
.Y(n_189)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx6_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_SL g406 ( 
.A1(n_200),
.A2(n_201),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_SL g344 ( 
.A1(n_201),
.A2(n_345),
.B(n_348),
.Y(n_344)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_215),
.Y(n_423)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_224),
.A2(n_384),
.B(n_386),
.Y(n_383)
);

BUFx24_ASAP7_75t_SL g438 ( 
.A(n_225),
.Y(n_438)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.CI(n_237),
.CON(n_225),
.SN(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_233),
.B2(n_236),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

AOI32xp33_ASAP7_75t_L g366 ( 
.A1(n_243),
.A2(n_349),
.A3(n_367),
.B1(n_368),
.B2(n_371),
.Y(n_366)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_245),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_416),
.B(n_435),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_394),
.B(n_415),
.Y(n_249)
);

AO21x1_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_375),
.B(n_393),
.Y(n_250)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_332),
.B(n_374),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_306),
.B(n_331),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_283),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_254),
.B(n_283),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_269),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_255),
.A2(n_269),
.B1(n_270),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_255),
.Y(n_329)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

INVx5_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_282),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_297),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_298),
.C(n_305),
.Y(n_333)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_304),
.B2(n_305),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g371 ( 
.A(n_301),
.B(n_372),
.Y(n_371)
);

INVx8_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_324),
.B(n_330),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_314),
.B(n_323),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_322),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_322),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_320),
.B(n_321),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_321),
.A2(n_354),
.B(n_363),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_328),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_334),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_352),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_342),
.B2(n_343),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_342),
.C(n_352),
.Y(n_376)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_366),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_366),
.Y(n_381)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_SL g357 ( 
.A(n_358),
.Y(n_357)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_376),
.B(n_377),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_382),
.B2(n_392),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_381),
.C(n_392),
.Y(n_395)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_382),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_387),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_388),
.C(n_389),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_395),
.B(n_396),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_403),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.Y(n_397)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_398),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_400),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_401),
.C(n_403),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_405),
.B1(n_411),
.B2(n_414),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_412),
.C(n_413),
.Y(n_426)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_411),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_430),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_419),
.A2(n_436),
.B(n_437),
.Y(n_435)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_427),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_427),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_424),
.C(n_426),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_424),
.A2(n_425),
.B1(n_426),
.B2(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_426),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_432),
.Y(n_436)
);


endmodule