module fake_jpeg_2829_n_441 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_47),
.B(n_56),
.Y(n_144)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g126 ( 
.A(n_48),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_15),
.C(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_0),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_62),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_65),
.Y(n_99)
);

NOR2xp67_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_14),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_18),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_86),
.Y(n_94)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_82),
.B(n_89),
.Y(n_129)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_40),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_25),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_40),
.B1(n_46),
.B2(n_28),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_96),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_36),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_97),
.B(n_86),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_45),
.B1(n_21),
.B2(n_37),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_103),
.A2(n_109),
.B(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_108),
.B(n_122),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_21),
.B1(n_37),
.B2(n_36),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_28),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_79),
.A2(n_26),
.B1(n_42),
.B2(n_30),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_69),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_73),
.A2(n_26),
.B1(n_30),
.B2(n_42),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_49),
.A2(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_52),
.A2(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_38),
.B1(n_33),
.B2(n_31),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_74),
.A2(n_37),
.B1(n_76),
.B2(n_53),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_147),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_48),
.B(n_84),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_148),
.A2(n_156),
.B(n_167),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_38),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_192),
.Y(n_197)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_77),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g236 ( 
.A(n_153),
.B(n_190),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_155),
.B(n_161),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_72),
.B(n_33),
.Y(n_156)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_76),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_166),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_167),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_60),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_169),
.Y(n_205)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_88),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_172),
.B(n_174),
.Y(n_233)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_31),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_17),
.B(n_85),
.C(n_86),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_186),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_93),
.B1(n_59),
.B2(n_70),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_194),
.B1(n_110),
.B2(n_124),
.Y(n_225)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_182),
.Y(n_228)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_138),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_181),
.Y(n_222)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

INVx11_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_127),
.B(n_87),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_75),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_189),
.B(n_191),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_115),
.B(n_80),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_106),
.B(n_131),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_196),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_120),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_132),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_101),
.B(n_17),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_114),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_147),
.A2(n_136),
.B1(n_139),
.B2(n_146),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_200),
.A2(n_237),
.B1(n_149),
.B2(n_175),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_141),
.B1(n_133),
.B2(n_109),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_217),
.B1(n_225),
.B2(n_227),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_150),
.B(n_103),
.CI(n_124),
.CON(n_211),
.SN(n_211)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_211),
.B(n_158),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_212),
.A2(n_158),
.B(n_153),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_101),
.B(n_142),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_236),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_159),
.A2(n_121),
.B1(n_110),
.B2(n_134),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_236),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_156),
.B(n_121),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_235),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_148),
.A2(n_134),
.B1(n_114),
.B2(n_5),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_179),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_234),
.B1(n_155),
.B2(n_157),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_179),
.B(n_160),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_154),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_181),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_244),
.A2(n_247),
.B(n_266),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_158),
.B1(n_194),
.B2(n_195),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_245),
.A2(n_254),
.B1(n_267),
.B2(n_273),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_246),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_249),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_180),
.C(n_153),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_270),
.C(n_271),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_253),
.B1(n_258),
.B2(n_215),
.Y(n_289)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_198),
.A2(n_153),
.B1(n_186),
.B2(n_188),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_198),
.A2(n_178),
.B1(n_151),
.B2(n_163),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g255 ( 
.A(n_228),
.B(n_164),
.Y(n_255)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_231),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_257),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_212),
.A2(n_173),
.B1(n_192),
.B2(n_152),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_202),
.Y(n_260)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

AO22x1_ASAP7_75t_SL g262 ( 
.A1(n_225),
.A2(n_182),
.B1(n_185),
.B2(n_171),
.Y(n_262)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_162),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_276),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_264),
.A2(n_268),
.B1(n_224),
.B2(n_205),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_265),
.A2(n_211),
.B1(n_216),
.B2(n_202),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_175),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_237),
.A2(n_170),
.B1(n_166),
.B2(n_169),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_221),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_219),
.A2(n_187),
.B(n_190),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_275),
.B(n_227),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_204),
.B(n_184),
.C(n_183),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_197),
.B(n_184),
.C(n_12),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_214),
.Y(n_272)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_272),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_220),
.A2(n_184),
.B1(n_12),
.B2(n_13),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_274),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_215),
.A2(n_9),
.B(n_12),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_9),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_281),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_245),
.A2(n_215),
.B1(n_220),
.B2(n_217),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_288),
.A2(n_295),
.B1(n_297),
.B2(n_251),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_293),
.B1(n_275),
.B2(n_269),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_265),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_197),
.C(n_214),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_301),
.C(n_303),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_243),
.A2(n_234),
.B1(n_211),
.B2(n_230),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_243),
.A2(n_229),
.B1(n_230),
.B2(n_209),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_248),
.A2(n_209),
.B1(n_207),
.B2(n_205),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_207),
.C(n_221),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_309),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_210),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_242),
.Y(n_308)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_239),
.A2(n_203),
.B1(n_205),
.B2(n_218),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_296),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_319),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_294),
.A2(n_239),
.B(n_244),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_312),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_255),
.C(n_268),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_329),
.C(n_336),
.Y(n_340)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_317),
.A2(n_279),
.B1(n_309),
.B2(n_305),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_318),
.B(n_277),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_256),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_292),
.A2(n_288),
.B1(n_278),
.B2(n_295),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_320),
.A2(n_325),
.B1(n_328),
.B2(n_331),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_276),
.Y(n_321)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_255),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_315),
.Y(n_349)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_323),
.Y(n_341)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_327),
.Y(n_348)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_286),
.Y(n_326)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_326),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_297),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_292),
.A2(n_247),
.B1(n_264),
.B2(n_253),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_280),
.B(n_265),
.C(n_240),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_294),
.A2(n_306),
.B(n_281),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_332),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_278),
.A2(n_258),
.B1(n_263),
.B2(n_266),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_304),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_306),
.A2(n_270),
.B(n_254),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_333),
.A2(n_335),
.B1(n_303),
.B2(n_299),
.Y(n_352)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_334),
.A2(n_199),
.B1(n_287),
.B2(n_206),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_285),
.B(n_252),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_271),
.C(n_272),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_338),
.A2(n_343),
.B1(n_346),
.B2(n_353),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_327),
.A2(n_290),
.B1(n_279),
.B2(n_284),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_345),
.B(n_314),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_337),
.A2(n_308),
.B1(n_283),
.B2(n_300),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_322),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_354),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_337),
.A2(n_277),
.B1(n_307),
.B2(n_262),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_320),
.A2(n_267),
.B1(n_307),
.B2(n_262),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_261),
.C(n_259),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_336),
.C(n_333),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_273),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_359),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_357),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_313),
.B(n_210),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_317),
.A2(n_328),
.B1(n_331),
.B2(n_310),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_310),
.Y(n_362)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_361),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_341),
.B1(n_314),
.B2(n_351),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_319),
.Y(n_363)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_373),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_370),
.C(n_371),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_SL g366 ( 
.A(n_340),
.B(n_330),
.C(n_318),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_358),
.C(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_342),
.Y(n_369)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_312),
.C(n_335),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_321),
.C(n_332),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_355),
.C(n_356),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_375),
.C(n_346),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_334),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_380),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_324),
.C(n_323),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_377),
.A2(n_351),
.B1(n_357),
.B2(n_287),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_344),
.B(n_316),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_381),
.B(n_338),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_344),
.Y(n_385)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_391),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_358),
.C(n_339),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_387),
.B(n_389),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_395),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_348),
.C(n_353),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_393),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_378),
.A2(n_354),
.B(n_341),
.Y(n_393)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_394),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_381),
.B(n_368),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_396),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_206),
.C(n_199),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_397),
.B(n_375),
.C(n_371),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_387),
.A2(n_376),
.B1(n_373),
.B2(n_367),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_400),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_401),
.B(n_408),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_391),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_382),
.B(n_386),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_407),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_383),
.A2(n_376),
.B1(n_379),
.B2(n_370),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_388),
.A2(n_262),
.B1(n_241),
.B2(n_218),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_226),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_410),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_411),
.B(n_420),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_384),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_412),
.B(n_415),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_406),
.A2(n_397),
.B(n_392),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_413),
.A2(n_401),
.B(n_400),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_395),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_226),
.Y(n_417)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_417),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_241),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_421),
.B(n_422),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_420),
.B(n_405),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_404),
.C(n_409),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_424),
.B(n_427),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_418),
.A2(n_404),
.B1(n_408),
.B2(n_409),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_416),
.C(n_414),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_432),
.C(n_422),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_426),
.B(n_419),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_429),
.A2(n_232),
.B(n_12),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_241),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_434),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_431),
.B(n_427),
.C(n_425),
.Y(n_434)
);

OAI21xp33_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_9),
.B(n_13),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_436),
.B(n_13),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_438),
.A2(n_430),
.B(n_437),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_439),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_428),
.Y(n_441)
);


endmodule