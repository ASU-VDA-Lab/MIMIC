module fake_netlist_6_1777_n_1243 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_298, n_18, n_21, n_193, n_147, n_269, n_258, n_281, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_283, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_296, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_299, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_297, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_285, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_292, n_129, n_13, n_121, n_294, n_302, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_286, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_291, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_284, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_301, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_289, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_282, n_58, n_116, n_280, n_211, n_287, n_64, n_220, n_288, n_290, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_300, n_107, n_10, n_295, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_293, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1243);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_298;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_281;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_283;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_296;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_299;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_297;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_285;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_292;
input n_129;
input n_13;
input n_121;
input n_294;
input n_302;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_286;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_291;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_284;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_301;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_289;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_282;
input n_58;
input n_116;
input n_280;
input n_211;
input n_287;
input n_64;
input n_220;
input n_288;
input n_290;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_300;
input n_107;
input n_10;
input n_295;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_293;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1243;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_530;
wire n_618;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_304;
wire n_694;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_899;
wire n_738;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1223;
wire n_303;
wire n_511;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_848;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_380;
wire n_1190;
wire n_397;
wire n_1213;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_234),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_29),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_283),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_246),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_116),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_5),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_245),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_152),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_30),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_111),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_26),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_177),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_10),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_174),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_47),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_226),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_205),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_298),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_268),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_85),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_279),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_183),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_212),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_280),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_93),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_127),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_191),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_225),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_110),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_158),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_265),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_289),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_27),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_285),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_240),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_138),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_165),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_61),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_113),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_182),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_184),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_203),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_192),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_204),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_166),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_128),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_145),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_230),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_160),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_176),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_187),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_276),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_112),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_216),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_213),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_251),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_154),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_147),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_100),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_195),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_118),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_256),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_278),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_150),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_142),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_64),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_141),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_26),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_44),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_218),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_281),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_51),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_11),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_301),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_223),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_20),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_198),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_125),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_266),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_84),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_159),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_30),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_77),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_185),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_5),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_267),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_269),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_53),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_114),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_290),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_76),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_233),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_19),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_206),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_169),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_252),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_56),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_272),
.Y(n_405)
);

BUFx10_ASAP7_75t_L g406 ( 
.A(n_270),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_248),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_295),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_57),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_247),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_124),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_93),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_60),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_28),
.B(n_144),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_167),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_238),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_14),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_57),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_146),
.Y(n_419)
);

INVxp33_ASAP7_75t_L g420 ( 
.A(n_66),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_91),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_229),
.B(n_25),
.Y(n_422)
);

BUFx8_ASAP7_75t_SL g423 ( 
.A(n_35),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_73),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_21),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_262),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_189),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_186),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_156),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_117),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_97),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_153),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_58),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_37),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_219),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_94),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_12),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_201),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_208),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_104),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_12),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_36),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_74),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_243),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_173),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_222),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_210),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_239),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_102),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_43),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_287),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_32),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_157),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_288),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_155),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_19),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_235),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_143),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_273),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_164),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_214),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_423),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_309),
.A2(n_319),
.B1(n_379),
.B2(n_376),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_312),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_312),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_329),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_383),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_314),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_313),
.B(n_105),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_314),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_313),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_314),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_303),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_3),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_401),
.B(n_3),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_395),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_417),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_314),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_456),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_418),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_305),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_419),
.B(n_4),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_315),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_313),
.Y(n_488)
);

INVxp33_ASAP7_75t_L g489 ( 
.A(n_450),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_419),
.B(n_4),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_375),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_324),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_314),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_313),
.B(n_106),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_330),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_401),
.B(n_6),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_420),
.B(n_6),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_366),
.Y(n_499)
);

BUFx12f_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_439),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_378),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_403),
.B(n_351),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_378),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_378),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_339),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_380),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_389),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g509 ( 
.A(n_403),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_420),
.A2(n_449),
.B1(n_317),
.B2(n_412),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_378),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_329),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_318),
.B(n_328),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_344),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_390),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_439),
.B(n_7),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

CKINVDCx11_ASAP7_75t_R g519 ( 
.A(n_320),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_356),
.B(n_8),
.Y(n_521)
);

INVx6_ASAP7_75t_L g522 ( 
.A(n_451),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_356),
.B(n_9),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_373),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_437),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_333),
.B(n_10),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_447),
.B(n_11),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_441),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_436),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_442),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_452),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_351),
.B(n_13),
.Y(n_533)
);

BUFx12f_ASAP7_75t_L g534 ( 
.A(n_387),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_451),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_304),
.Y(n_536)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_348),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g539 ( 
.A(n_357),
.B(n_13),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_488),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_509),
.B(n_427),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_513),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_488),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_535),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_535),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_535),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_513),
.B(n_453),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_469),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_488),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_502),
.Y(n_550)
);

NOR2x1p5_ASAP7_75t_L g551 ( 
.A(n_503),
.B(n_398),
.Y(n_551)
);

AO21x2_ASAP7_75t_L g552 ( 
.A1(n_533),
.A2(n_422),
.B(n_414),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_482),
.B(n_404),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_536),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_519),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_469),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_485),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_487),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_502),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_505),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_489),
.A2(n_483),
.B1(n_497),
.B2(n_477),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_474),
.B(n_448),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_505),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_468),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_518),
.Y(n_565)
);

NOR3xp33_ASAP7_75t_L g566 ( 
.A(n_510),
.B(n_400),
.C(n_392),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_522),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_521),
.B(n_323),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_501),
.B(n_460),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_495),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_519),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_470),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_523),
.A2(n_368),
.B1(n_433),
.B2(n_409),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_473),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_499),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_520),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_481),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_534),
.B(n_404),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_528),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_500),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_493),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_472),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_503),
.A2(n_424),
.B1(n_434),
.B2(n_411),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_504),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_514),
.B(n_340),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_539),
.B(n_346),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_564),
.B(n_504),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_559),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_564),
.B(n_573),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_573),
.B(n_511),
.Y(n_591)
);

AOI221xp5_ASAP7_75t_L g592 ( 
.A1(n_561),
.A2(n_510),
.B1(n_498),
.B2(n_475),
.C(n_497),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_547),
.B(n_506),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_562),
.B(n_526),
.Y(n_594)
);

O2A1O1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_587),
.A2(n_477),
.B(n_533),
.C(n_475),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_586),
.B(n_491),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_541),
.A2(n_539),
.B1(n_537),
.B2(n_527),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_557),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_568),
.B(n_537),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_542),
.B(n_462),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_574),
.A2(n_537),
.B1(n_524),
.B2(n_498),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_569),
.B(n_476),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_558),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_552),
.A2(n_490),
.B1(n_517),
.B2(n_486),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_SL g605 ( 
.A(n_548),
.B(n_353),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_540),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_542),
.B(n_489),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_542),
.B(n_524),
.Y(n_608)
);

NOR2x1p5_ASAP7_75t_L g609 ( 
.A(n_581),
.B(n_496),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_585),
.B(n_517),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_585),
.B(n_397),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_571),
.Y(n_612)
);

BUFx8_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_554),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_575),
.B(n_469),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_575),
.B(n_469),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_584),
.B(n_466),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_553),
.Y(n_618)
);

NAND3xp33_ASAP7_75t_L g619 ( 
.A(n_566),
.B(n_512),
.C(n_465),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_549),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_549),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_545),
.B(n_463),
.C(n_515),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_563),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_563),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_583),
.B(n_445),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_583),
.A2(n_332),
.B(n_464),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_543),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_543),
.Y(n_628)
);

AND2x2_ASAP7_75t_SL g629 ( 
.A(n_556),
.B(n_424),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_578),
.B(n_494),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_550),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_550),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_544),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_544),
.B(n_522),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_570),
.B(n_482),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_552),
.A2(n_494),
.B1(n_411),
.B2(n_426),
.Y(n_636)
);

AND2x2_ASAP7_75t_SL g637 ( 
.A(n_556),
.B(n_353),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_540),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_L g639 ( 
.A(n_546),
.B(n_463),
.C(n_515),
.Y(n_639)
);

AND2x6_ASAP7_75t_SL g640 ( 
.A(n_579),
.B(n_507),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_567),
.B(n_471),
.Y(n_641)
);

AND2x6_ASAP7_75t_SL g642 ( 
.A(n_579),
.B(n_508),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_SL g643 ( 
.A1(n_572),
.A2(n_467),
.B1(n_494),
.B2(n_306),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_551),
.A2(n_467),
.B1(n_538),
.B2(n_479),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_560),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_552),
.B(n_478),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_540),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_565),
.B(n_480),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_579),
.A2(n_308),
.B1(n_316),
.B2(n_311),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_633),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_593),
.B(n_553),
.Y(n_651)
);

O2A1O1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_595),
.A2(n_516),
.B(n_530),
.C(n_525),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_597),
.B(n_556),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_607),
.B(n_581),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_596),
.B(n_618),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_598),
.Y(n_656)
);

BUFx8_ASAP7_75t_SL g657 ( 
.A(n_633),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_604),
.B(n_582),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_592),
.A2(n_629),
.B1(n_594),
.B2(n_637),
.Y(n_659)
);

AOI21x1_ASAP7_75t_L g660 ( 
.A1(n_615),
.A2(n_310),
.B(n_307),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_617),
.A2(n_531),
.B(n_532),
.C(n_484),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_SL g662 ( 
.A(n_601),
.B(n_555),
.C(n_572),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_611),
.B(n_636),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_625),
.B(n_321),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_599),
.A2(n_432),
.B1(n_435),
.B2(n_428),
.Y(n_665)
);

O2A1O1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_644),
.A2(n_455),
.B(n_461),
.C(n_435),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_619),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_603),
.B(n_579),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_615),
.A2(n_461),
.B(n_455),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_633),
.B(n_322),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_635),
.B(n_325),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_612),
.B(n_326),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_641),
.Y(n_673)
);

O2A1O1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_626),
.A2(n_614),
.B(n_590),
.C(n_616),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_620),
.B(n_327),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_621),
.B(n_334),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_590),
.A2(n_335),
.B(n_342),
.C(n_336),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_622),
.A2(n_345),
.B1(n_347),
.B2(n_343),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_639),
.A2(n_337),
.B1(n_338),
.B2(n_331),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_623),
.B(n_349),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_608),
.B(n_341),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_616),
.A2(n_354),
.B(n_352),
.Y(n_682)
);

OAI22x1_ASAP7_75t_L g683 ( 
.A1(n_643),
.A2(n_538),
.B1(n_360),
.B2(n_361),
.Y(n_683)
);

OAI21xp33_ASAP7_75t_L g684 ( 
.A1(n_648),
.A2(n_580),
.B(n_577),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_649),
.B(n_350),
.Y(n_685)
);

OAI321xp33_ASAP7_75t_L g686 ( 
.A1(n_634),
.A2(n_367),
.A3(n_362),
.B1(n_369),
.B2(n_363),
.C(n_355),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_624),
.B(n_371),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_609),
.B(n_492),
.Y(n_688)
);

BUFx8_ASAP7_75t_L g689 ( 
.A(n_613),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_588),
.B(n_372),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_640),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_627),
.B(n_492),
.Y(n_692)
);

CKINVDCx6p67_ASAP7_75t_R g693 ( 
.A(n_613),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_647),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_SL g695 ( 
.A(n_588),
.B(n_358),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_630),
.A2(n_393),
.B(n_391),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_630),
.A2(n_591),
.B(n_589),
.Y(n_697)
);

NOR2x1_ASAP7_75t_L g698 ( 
.A(n_606),
.B(n_394),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_628),
.A2(n_399),
.B1(n_402),
.B2(n_396),
.Y(n_699)
);

OAI21xp33_ASAP7_75t_L g700 ( 
.A1(n_632),
.A2(n_529),
.B(n_407),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_591),
.A2(n_408),
.B(n_410),
.C(n_405),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_606),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_645),
.Y(n_703)
);

A2O1A1Ixp33_ASAP7_75t_SL g704 ( 
.A1(n_605),
.A2(n_430),
.B(n_438),
.C(n_416),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_638),
.B(n_440),
.Y(n_705)
);

CKINVDCx6p67_ASAP7_75t_R g706 ( 
.A(n_642),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_638),
.B(n_454),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_598),
.B(n_457),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_592),
.A2(n_364),
.B1(n_365),
.B2(n_359),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_610),
.A2(n_374),
.B(n_370),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_604),
.B(n_377),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_598),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_598),
.Y(n_713)
);

AOI21xp33_ASAP7_75t_L g714 ( 
.A1(n_595),
.A2(n_382),
.B(n_381),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_604),
.B(n_384),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_610),
.A2(n_386),
.B(n_385),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_R g717 ( 
.A(n_594),
.B(n_388),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_618),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_602),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_593),
.B(n_415),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_633),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_593),
.B(n_429),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_610),
.A2(n_446),
.B(n_444),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_633),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_646),
.A2(n_459),
.B(n_458),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_593),
.B(n_14),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_607),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_631),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_604),
.A2(n_108),
.B1(n_109),
.B2(n_107),
.Y(n_729)
);

AO21x1_ASAP7_75t_L g730 ( 
.A1(n_595),
.A2(n_15),
.B(n_16),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_597),
.B(n_15),
.Y(n_731)
);

O2A1O1Ixp33_ASAP7_75t_SL g732 ( 
.A1(n_617),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_732)
);

CKINVDCx6p67_ASAP7_75t_R g733 ( 
.A(n_600),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_604),
.B(n_115),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_651),
.B(n_17),
.Y(n_735)
);

OA22x2_ASAP7_75t_L g736 ( 
.A1(n_709),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_736)
);

AOI31xp67_ASAP7_75t_L g737 ( 
.A1(n_653),
.A2(n_120),
.A3(n_121),
.B(n_119),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_667),
.A2(n_123),
.B1(n_126),
.B2(n_122),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_658),
.A2(n_674),
.B(n_734),
.Y(n_739)
);

O2A1O1Ixp5_ASAP7_75t_SL g740 ( 
.A1(n_665),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_655),
.B(n_22),
.Y(n_741)
);

INVx3_ASAP7_75t_SL g742 ( 
.A(n_693),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_688),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_728),
.A2(n_302),
.B(n_130),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_712),
.Y(n_745)
);

OA21x2_ASAP7_75t_L g746 ( 
.A1(n_669),
.A2(n_131),
.B(n_129),
.Y(n_746)
);

AOI221xp5_ASAP7_75t_L g747 ( 
.A1(n_726),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.C(n_27),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_711),
.A2(n_133),
.B1(n_134),
.B2(n_132),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_719),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_721),
.B(n_135),
.Y(n_750)
);

OA21x2_ASAP7_75t_L g751 ( 
.A1(n_696),
.A2(n_137),
.B(n_136),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_720),
.B(n_29),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_656),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_709),
.A2(n_725),
.B(n_685),
.C(n_722),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_715),
.A2(n_140),
.B(n_139),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_713),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_681),
.B(n_31),
.C(n_32),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_730),
.A2(n_34),
.A3(n_31),
.B(n_33),
.Y(n_758)
);

BUFx2_ASAP7_75t_SL g759 ( 
.A(n_724),
.Y(n_759)
);

NOR2x1_ASAP7_75t_SL g760 ( 
.A(n_729),
.B(n_148),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_673),
.B(n_34),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_705),
.A2(n_151),
.B(n_149),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_703),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_SL g764 ( 
.A1(n_731),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_650),
.Y(n_765)
);

INVx5_ASAP7_75t_L g766 ( 
.A(n_657),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_707),
.A2(n_299),
.B(n_161),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_718),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_708),
.Y(n_769)
);

OAI21xp33_ASAP7_75t_SL g770 ( 
.A1(n_690),
.A2(n_40),
.B(n_41),
.Y(n_770)
);

OA21x2_ASAP7_75t_L g771 ( 
.A1(n_682),
.A2(n_163),
.B(n_162),
.Y(n_771)
);

INVx6_ASAP7_75t_L g772 ( 
.A(n_689),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_666),
.A2(n_652),
.B(n_714),
.C(n_668),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_654),
.B(n_41),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_672),
.B(n_42),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_R g776 ( 
.A(n_717),
.B(n_168),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_695),
.B(n_42),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_661),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_678),
.A2(n_171),
.B1(n_175),
.B2(n_170),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_664),
.B(n_43),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_683),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_SL g782 ( 
.A(n_686),
.B(n_45),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_660),
.A2(n_297),
.B(n_178),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_675),
.B(n_676),
.Y(n_784)
);

OR2x6_ASAP7_75t_L g785 ( 
.A(n_691),
.B(n_46),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_680),
.B(n_47),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_687),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_787)
);

INVx3_ASAP7_75t_SL g788 ( 
.A(n_733),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_684),
.B(n_49),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_702),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_710),
.B(n_50),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_689),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_679),
.B(n_51),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_716),
.B(n_52),
.Y(n_794)
);

AOI21xp33_ASAP7_75t_L g795 ( 
.A1(n_671),
.A2(n_52),
.B(n_53),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_670),
.A2(n_180),
.B1(n_181),
.B2(n_179),
.Y(n_796)
);

AO22x2_ASAP7_75t_L g797 ( 
.A1(n_662),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_SL g798 ( 
.A1(n_677),
.A2(n_58),
.B(n_54),
.C(n_55),
.Y(n_798)
);

OR2x6_ASAP7_75t_L g799 ( 
.A(n_701),
.B(n_59),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_698),
.A2(n_220),
.B1(n_294),
.B2(n_293),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_SL g801 ( 
.A1(n_704),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_801)
);

OR2x6_ASAP7_75t_L g802 ( 
.A(n_700),
.B(n_62),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_723),
.B(n_63),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_694),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_699),
.B(n_64),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_732),
.B(n_65),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_706),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_657),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_651),
.B(n_67),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_719),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_651),
.B(n_67),
.Y(n_811)
);

BUFx2_ASAP7_75t_SL g812 ( 
.A(n_721),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_651),
.B(n_68),
.Y(n_813)
);

BUFx12f_ASAP7_75t_L g814 ( 
.A(n_689),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_656),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_692),
.Y(n_816)
);

O2A1O1Ixp5_ASAP7_75t_SL g817 ( 
.A1(n_665),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_817)
);

AOI21xp33_ASAP7_75t_L g818 ( 
.A1(n_685),
.A2(n_72),
.B(n_73),
.Y(n_818)
);

AO31x2_ASAP7_75t_L g819 ( 
.A1(n_730),
.A2(n_72),
.A3(n_74),
.B(n_75),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_697),
.A2(n_296),
.B(n_190),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_663),
.A2(n_193),
.B(n_188),
.Y(n_821)
);

AO22x1_ASAP7_75t_L g822 ( 
.A1(n_685),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_651),
.B(n_78),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_663),
.A2(n_196),
.B(n_194),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_688),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_651),
.B(n_78),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_659),
.A2(n_232),
.B1(n_292),
.B2(n_291),
.Y(n_827)
);

INVx6_ASAP7_75t_L g828 ( 
.A(n_689),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_663),
.A2(n_199),
.B(n_197),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_650),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_692),
.Y(n_831)
);

OAI22x1_ASAP7_75t_L g832 ( 
.A1(n_659),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_692),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_656),
.Y(n_834)
);

AO31x2_ASAP7_75t_L g835 ( 
.A1(n_730),
.A2(n_82),
.A3(n_83),
.B(n_84),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_651),
.B(n_82),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_663),
.A2(n_202),
.B(n_200),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_692),
.Y(n_838)
);

OAI21xp33_ASAP7_75t_SL g839 ( 
.A1(n_659),
.A2(n_86),
.B(n_87),
.Y(n_839)
);

AOI221xp5_ASAP7_75t_L g840 ( 
.A1(n_726),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.C(n_90),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_719),
.B(n_88),
.Y(n_841)
);

BUFx8_ASAP7_75t_SL g842 ( 
.A(n_657),
.Y(n_842)
);

AO31x2_ASAP7_75t_L g843 ( 
.A1(n_730),
.A2(n_89),
.A3(n_91),
.B(n_92),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_663),
.A2(n_237),
.B(n_286),
.Y(n_844)
);

NOR2x1_ASAP7_75t_SL g845 ( 
.A(n_729),
.B(n_207),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_727),
.B(n_92),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_650),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_SL g848 ( 
.A1(n_663),
.A2(n_236),
.B(n_282),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_692),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_651),
.B(n_94),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_754),
.B(n_784),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_759),
.B(n_95),
.Y(n_852)
);

AO31x2_ASAP7_75t_L g853 ( 
.A1(n_773),
.A2(n_95),
.A3(n_96),
.B(n_97),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_745),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_756),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_753),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_812),
.B(n_96),
.Y(n_857)
);

OA21x2_ASAP7_75t_L g858 ( 
.A1(n_824),
.A2(n_241),
.B(n_277),
.Y(n_858)
);

OA21x2_ASAP7_75t_L g859 ( 
.A1(n_755),
.A2(n_231),
.B(n_275),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_L g860 ( 
.A(n_774),
.B(n_98),
.C(n_99),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_815),
.Y(n_861)
);

OA21x2_ASAP7_75t_L g862 ( 
.A1(n_820),
.A2(n_228),
.B(n_274),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_810),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_752),
.B(n_811),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_834),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_765),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_765),
.B(n_209),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_763),
.Y(n_868)
);

BUFx12f_ASAP7_75t_L g869 ( 
.A(n_814),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_830),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_SL g871 ( 
.A1(n_793),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_871)
);

OA21x2_ASAP7_75t_L g872 ( 
.A1(n_744),
.A2(n_244),
.B(n_264),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_816),
.Y(n_873)
);

AO31x2_ASAP7_75t_L g874 ( 
.A1(n_778),
.A2(n_101),
.A3(n_102),
.B(n_103),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_831),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_842),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_833),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_768),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_783),
.A2(n_249),
.B(n_211),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_838),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_766),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_823),
.B(n_103),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_830),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_849),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_818),
.B(n_775),
.C(n_747),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_741),
.B(n_215),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_735),
.B(n_217),
.Y(n_887)
);

OA21x2_ASAP7_75t_L g888 ( 
.A1(n_821),
.A2(n_837),
.B(n_829),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_766),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_804),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_781),
.B(n_221),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_809),
.B(n_813),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_790),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_769),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_766),
.Y(n_895)
);

INVx6_ASAP7_75t_L g896 ( 
.A(n_772),
.Y(n_896)
);

CKINVDCx11_ASAP7_75t_R g897 ( 
.A(n_742),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_846),
.B(n_224),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_767),
.A2(n_227),
.B(n_250),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_789),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_841),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_847),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_805),
.B(n_253),
.Y(n_903)
);

OA21x2_ASAP7_75t_L g904 ( 
.A1(n_844),
.A2(n_254),
.B(n_255),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_761),
.B(n_257),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_826),
.A2(n_850),
.B(n_836),
.Y(n_906)
);

CKINVDCx8_ASAP7_75t_R g907 ( 
.A(n_808),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_746),
.A2(n_258),
.B(n_259),
.Y(n_908)
);

OA21x2_ASAP7_75t_L g909 ( 
.A1(n_786),
.A2(n_260),
.B(n_261),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_772),
.B(n_263),
.Y(n_910)
);

CKINVDCx11_ASAP7_75t_R g911 ( 
.A(n_788),
.Y(n_911)
);

BUFx12f_ASAP7_75t_L g912 ( 
.A(n_828),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_806),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_777),
.A2(n_795),
.B(n_780),
.C(n_839),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_750),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_750),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_791),
.A2(n_803),
.B(n_794),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_748),
.A2(n_848),
.B(n_771),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_782),
.B(n_840),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_828),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_832),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_736),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_792),
.B(n_802),
.Y(n_923)
);

AO31x2_ASAP7_75t_L g924 ( 
.A1(n_779),
.A2(n_817),
.A3(n_740),
.B(n_737),
.Y(n_924)
);

OA21x2_ASAP7_75t_L g925 ( 
.A1(n_757),
.A2(n_738),
.B(n_796),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_787),
.B(n_770),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_807),
.B(n_785),
.Y(n_927)
);

OAI21x1_ASAP7_75t_SL g928 ( 
.A1(n_751),
.A2(n_800),
.B(n_762),
.Y(n_928)
);

BUFx2_ASAP7_75t_SL g929 ( 
.A(n_762),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_764),
.B(n_822),
.Y(n_930)
);

OAI21x1_ASAP7_75t_L g931 ( 
.A1(n_776),
.A2(n_798),
.B(n_801),
.Y(n_931)
);

OAI21xp33_ASAP7_75t_SL g932 ( 
.A1(n_799),
.A2(n_785),
.B(n_797),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_819),
.A2(n_843),
.B(n_835),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_758),
.B(n_651),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_749),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_745),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_743),
.B(n_825),
.Y(n_937)
);

AO21x2_ASAP7_75t_L g938 ( 
.A1(n_739),
.A2(n_754),
.B(n_773),
.Y(n_938)
);

OAI21x1_ASAP7_75t_SL g939 ( 
.A1(n_760),
.A2(n_845),
.B(n_730),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_749),
.B(n_810),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_745),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_749),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_754),
.B(n_651),
.Y(n_943)
);

NAND2x1p5_ASAP7_75t_L g944 ( 
.A(n_765),
.B(n_830),
.Y(n_944)
);

NAND2x1p5_ASAP7_75t_L g945 ( 
.A(n_765),
.B(n_830),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_745),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_745),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_754),
.A2(n_739),
.B(n_663),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_749),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_745),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_753),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_754),
.A2(n_659),
.B(n_595),
.C(n_752),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_743),
.B(n_825),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_743),
.B(n_825),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_814),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_754),
.A2(n_659),
.B(n_595),
.C(n_752),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_745),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_753),
.Y(n_958)
);

AND2x6_ASAP7_75t_L g959 ( 
.A(n_827),
.B(n_659),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_745),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_754),
.A2(n_739),
.B(n_663),
.Y(n_961)
);

AO31x2_ASAP7_75t_L g962 ( 
.A1(n_754),
.A2(n_730),
.A3(n_773),
.B(n_739),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_936),
.Y(n_963)
);

OR2x6_ASAP7_75t_L g964 ( 
.A(n_912),
.B(n_910),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_947),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_854),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_863),
.Y(n_967)
);

NAND2x1p5_ASAP7_75t_L g968 ( 
.A(n_915),
.B(n_916),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_903),
.B(n_901),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_851),
.B(n_900),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_855),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_941),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_946),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_935),
.Y(n_974)
);

AO21x2_ASAP7_75t_L g975 ( 
.A1(n_928),
.A2(n_961),
.B(n_948),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_949),
.B(n_921),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_950),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_957),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_960),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_875),
.B(n_884),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_940),
.B(n_942),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_910),
.B(n_923),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_952),
.A2(n_956),
.B(n_943),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_892),
.B(n_864),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_900),
.B(n_913),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_870),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_873),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_922),
.B(n_923),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_959),
.B(n_906),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_938),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_877),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_880),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_878),
.B(n_894),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_868),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_856),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_861),
.B(n_865),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_951),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_958),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_883),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_959),
.B(n_919),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_885),
.A2(n_933),
.B(n_917),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_890),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_893),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_934),
.Y(n_1004)
);

AO21x2_ASAP7_75t_L g1005 ( 
.A1(n_928),
.A2(n_939),
.B(n_918),
.Y(n_1005)
);

BUFx2_ASAP7_75t_SL g1006 ( 
.A(n_907),
.Y(n_1006)
);

AOI211xp5_ASAP7_75t_L g1007 ( 
.A1(n_932),
.A2(n_860),
.B(n_914),
.C(n_891),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_870),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_870),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_962),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_896),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_898),
.B(n_905),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_944),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_871),
.B(n_937),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_896),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_866),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_959),
.B(n_886),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_902),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_937),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_959),
.B(n_926),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_945),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_882),
.B(n_953),
.Y(n_1022)
);

INVx5_ASAP7_75t_L g1023 ( 
.A(n_852),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_931),
.A2(n_908),
.B(n_887),
.Y(n_1024)
);

CKINVDCx16_ASAP7_75t_R g1025 ( 
.A(n_876),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_954),
.B(n_857),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_930),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_852),
.B(n_857),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_853),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_920),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_867),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_853),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_853),
.Y(n_1033)
);

BUFx4f_ASAP7_75t_SL g1034 ( 
.A(n_869),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_927),
.B(n_881),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_889),
.B(n_895),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_874),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_955),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_874),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_925),
.Y(n_1040)
);

INVxp33_ASAP7_75t_L g1041 ( 
.A(n_911),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_874),
.B(n_897),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_929),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_858),
.B(n_924),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_909),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_909),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_963),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_967),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_982),
.B(n_899),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_967),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_984),
.B(n_924),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_981),
.B(n_859),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_969),
.B(n_904),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1014),
.B(n_879),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_1011),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_976),
.B(n_862),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_980),
.B(n_988),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_972),
.Y(n_1058)
);

AND2x4_ASAP7_75t_SL g1059 ( 
.A(n_964),
.B(n_929),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_1011),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_974),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_974),
.B(n_872),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_1030),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_972),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_978),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1022),
.B(n_888),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1026),
.B(n_1019),
.Y(n_1067)
);

CKINVDCx14_ASAP7_75t_R g1068 ( 
.A(n_964),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_1010),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_1000),
.B(n_1020),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_1000),
.B(n_1020),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1042),
.B(n_997),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_1025),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_990),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_1034),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_1045),
.A2(n_1046),
.A3(n_1029),
.B(n_1037),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_993),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_965),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1027),
.B(n_995),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1027),
.B(n_998),
.Y(n_1080)
);

AND2x4_ASAP7_75t_SL g1081 ( 
.A(n_964),
.B(n_982),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_985),
.B(n_989),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1003),
.B(n_996),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1031),
.B(n_982),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_1008),
.B(n_1013),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_999),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_987),
.B(n_991),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_966),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_971),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_985),
.B(n_989),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_992),
.B(n_1008),
.Y(n_1091)
);

INVx2_ASAP7_75t_R g1092 ( 
.A(n_1039),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_970),
.B(n_1004),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1035),
.B(n_1017),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_973),
.B(n_977),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_979),
.B(n_994),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1002),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1007),
.B(n_1028),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_1038),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1012),
.A2(n_983),
.B1(n_1017),
.B2(n_975),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_968),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1032),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1033),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_1021),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_986),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_983),
.B(n_1012),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_1021),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1048),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1070),
.B(n_1040),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1078),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1082),
.B(n_1023),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1102),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1071),
.B(n_1040),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1051),
.B(n_975),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1103),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1066),
.B(n_1100),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1076),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1088),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1100),
.B(n_1001),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1089),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_1050),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1090),
.B(n_1023),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1097),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1053),
.B(n_1072),
.Y(n_1124)
);

AND2x4_ASAP7_75t_SL g1125 ( 
.A(n_1084),
.B(n_1036),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_1059),
.Y(n_1126)
);

INVxp67_ASAP7_75t_SL g1127 ( 
.A(n_1061),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_1055),
.B(n_1023),
.Y(n_1128)
);

INVxp67_ASAP7_75t_SL g1129 ( 
.A(n_1069),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_1069),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1094),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1058),
.Y(n_1132)
);

INVxp67_ASAP7_75t_L g1133 ( 
.A(n_1086),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1056),
.B(n_1064),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1065),
.B(n_1005),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_1060),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1077),
.B(n_1023),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1098),
.B(n_1057),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1073),
.B(n_1006),
.Y(n_1139)
);

NOR2xp67_ASAP7_75t_L g1140 ( 
.A(n_1055),
.B(n_1015),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1052),
.B(n_1044),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_1060),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1077),
.B(n_1043),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1091),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1083),
.B(n_1043),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1074),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1074),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1047),
.B(n_1005),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1112),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1115),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1124),
.B(n_1067),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1125),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1131),
.B(n_1062),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1116),
.B(n_1114),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1130),
.B(n_1049),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1124),
.B(n_1106),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1146),
.Y(n_1157)
);

AOI211xp5_ASAP7_75t_L g1158 ( 
.A1(n_1137),
.A2(n_1106),
.B(n_1041),
.C(n_1054),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1138),
.A2(n_1068),
.B1(n_1073),
.B2(n_1081),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1110),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_1130),
.B(n_1049),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1116),
.B(n_1114),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1118),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1141),
.B(n_1076),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1120),
.Y(n_1165)
);

OAI21xp33_ASAP7_75t_L g1166 ( 
.A1(n_1111),
.A2(n_1093),
.B(n_1079),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1135),
.B(n_1059),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1145),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1123),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1122),
.B(n_1093),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1119),
.B(n_1092),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1119),
.B(n_1148),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1146),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1147),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1147),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1144),
.B(n_1085),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1108),
.B(n_1080),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1132),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_1170),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1149),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1149),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1170),
.B(n_1127),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1150),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1154),
.B(n_1109),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1157),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1177),
.B(n_1109),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1156),
.B(n_1113),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1166),
.B(n_1143),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1160),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1157),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1162),
.B(n_1153),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1155),
.B(n_1117),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1168),
.B(n_1133),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1173),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1158),
.A2(n_1129),
.B(n_1024),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1162),
.B(n_1134),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1159),
.A2(n_1121),
.B1(n_1049),
.B2(n_1136),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1172),
.B(n_1176),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1172),
.B(n_1171),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1199),
.B(n_1198),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1179),
.B(n_1142),
.Y(n_1201)
);

OAI221xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1195),
.A2(n_1188),
.B1(n_1182),
.B2(n_1068),
.C(n_1161),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1180),
.Y(n_1203)
);

OAI321xp33_ASAP7_75t_L g1204 ( 
.A1(n_1188),
.A2(n_1161),
.A3(n_1155),
.B1(n_1175),
.B2(n_1174),
.C(n_1164),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1185),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1181),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1187),
.B(n_1186),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1197),
.B(n_1151),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1185),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1193),
.B(n_1192),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1190),
.Y(n_1211)
);

NOR3xp33_ASAP7_75t_L g1212 ( 
.A(n_1193),
.B(n_1139),
.C(n_1126),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1192),
.A2(n_1081),
.B(n_1041),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1202),
.A2(n_1194),
.B(n_1189),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1208),
.A2(n_1152),
.B1(n_1167),
.B2(n_1155),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1213),
.B(n_1099),
.Y(n_1216)
);

NOR3xp33_ASAP7_75t_L g1217 ( 
.A(n_1204),
.B(n_1140),
.C(n_1128),
.Y(n_1217)
);

AOI211xp5_ASAP7_75t_L g1218 ( 
.A1(n_1208),
.A2(n_1163),
.B(n_1165),
.C(n_1169),
.Y(n_1218)
);

OAI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1212),
.A2(n_1191),
.B1(n_1161),
.B2(n_1178),
.C(n_1190),
.Y(n_1219)
);

AOI211xp5_ASAP7_75t_L g1220 ( 
.A1(n_1210),
.A2(n_1192),
.B(n_1183),
.C(n_1063),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1214),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1220),
.A2(n_1218),
.B1(n_1215),
.B2(n_1219),
.Y(n_1222)
);

NAND4xp25_ASAP7_75t_SL g1223 ( 
.A(n_1217),
.B(n_1075),
.C(n_1207),
.D(n_1196),
.Y(n_1223)
);

NOR3xp33_ASAP7_75t_L g1224 ( 
.A(n_1216),
.B(n_1210),
.C(n_1201),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1214),
.B(n_1200),
.Y(n_1225)
);

AOI222xp33_ASAP7_75t_L g1226 ( 
.A1(n_1221),
.A2(n_1222),
.B1(n_1223),
.B2(n_1201),
.C1(n_1205),
.C2(n_1171),
.Y(n_1226)
);

AOI211xp5_ASAP7_75t_L g1227 ( 
.A1(n_1224),
.A2(n_1206),
.B(n_1203),
.C(n_1063),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1225),
.B(n_1199),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1224),
.B(n_1184),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1221),
.B(n_1184),
.Y(n_1230)
);

NOR2xp67_ASAP7_75t_L g1231 ( 
.A(n_1229),
.B(n_1230),
.Y(n_1231)
);

NAND4xp25_ASAP7_75t_L g1232 ( 
.A(n_1226),
.B(n_1030),
.C(n_1104),
.D(n_1107),
.Y(n_1232)
);

NAND4xp25_ASAP7_75t_L g1233 ( 
.A(n_1227),
.B(n_1104),
.C(n_1107),
.D(n_1152),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1232),
.B(n_1228),
.C(n_1101),
.Y(n_1234)
);

NAND4xp25_ASAP7_75t_L g1235 ( 
.A(n_1231),
.B(n_1087),
.C(n_1096),
.D(n_1095),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1235),
.B(n_1233),
.Y(n_1236)
);

XNOR2xp5_ASAP7_75t_L g1237 ( 
.A(n_1236),
.B(n_1075),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1237),
.B(n_1234),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_SL g1239 ( 
.A1(n_1238),
.A2(n_1034),
.B(n_1099),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1239),
.A2(n_1125),
.B1(n_1211),
.B2(n_1209),
.Y(n_1240)
);

INVxp67_ASAP7_75t_L g1241 ( 
.A(n_1240),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1241),
.A2(n_1018),
.B(n_1016),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1242),
.A2(n_1105),
.B1(n_1085),
.B2(n_1009),
.Y(n_1243)
);


endmodule