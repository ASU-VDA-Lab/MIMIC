module fake_jpeg_30805_n_314 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_10),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_28),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_55),
.B(n_60),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_24),
.B1(n_25),
.B2(n_19),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_57),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_37),
.B1(n_19),
.B2(n_20),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_58),
.A2(n_73),
.B1(n_87),
.B2(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_68),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_70),
.B(n_79),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_19),
.B1(n_21),
.B2(n_20),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_76),
.B1(n_81),
.B2(n_82),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_24),
.B1(n_25),
.B2(n_21),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_20),
.B1(n_24),
.B2(n_23),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_20),
.B1(n_38),
.B2(n_36),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_25),
.B1(n_38),
.B2(n_20),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_25),
.B1(n_38),
.B2(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_36),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_49),
.B1(n_53),
.B2(n_44),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_83),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_26),
.B1(n_32),
.B2(n_18),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_44),
.A2(n_32),
.B1(n_30),
.B2(n_25),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_34),
.B1(n_27),
.B2(n_4),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_65),
.B1(n_27),
.B2(n_39),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_12),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_14),
.Y(n_96)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g134 ( 
.A(n_99),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

HAxp5_ASAP7_75t_SL g101 ( 
.A(n_69),
.B(n_52),
.CON(n_101),
.SN(n_101)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_61),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_103),
.Y(n_142)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_27),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_127),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_33),
.B1(n_22),
.B2(n_66),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_42),
.B1(n_48),
.B2(n_51),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_128),
.B1(n_89),
.B2(n_51),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_76),
.B1(n_71),
.B2(n_64),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_126),
.B1(n_86),
.B2(n_67),
.Y(n_141)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_39),
.B(n_48),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_80),
.C(n_73),
.Y(n_130)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_122),
.Y(n_133)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_67),
.B1(n_74),
.B2(n_33),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_60),
.A2(n_70),
.B1(n_80),
.B2(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_22),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_62),
.A2(n_51),
.B1(n_48),
.B2(n_33),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_109),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_131),
.A2(n_159),
.B1(n_112),
.B2(n_108),
.Y(n_181)
);

OR2x4_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_66),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_123),
.B(n_119),
.C(n_116),
.D(n_128),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_86),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_152),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_145),
.B1(n_148),
.B2(n_103),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_115),
.B1(n_95),
.B2(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_74),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_0),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_93),
.B(n_1),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_93),
.B(n_11),
.C(n_4),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_5),
.C(n_6),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_95),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_142),
.B1(n_124),
.B2(n_150),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_119),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_163),
.B(n_165),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_121),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_164),
.B(n_167),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_119),
.C(n_118),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_166),
.A2(n_12),
.B(n_13),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_133),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_107),
.B1(n_92),
.B2(n_98),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_171),
.B1(n_177),
.B2(n_182),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_99),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_169),
.B(n_170),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_132),
.Y(n_170)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_173),
.Y(n_206)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_133),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_185),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_122),
.B1(n_120),
.B2(n_105),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_184),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_117),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_186),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_144),
.B1(n_151),
.B2(n_149),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_129),
.A2(n_130),
.B1(n_137),
.B2(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_155),
.B(n_5),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_6),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_7),
.Y(n_204)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_189),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_91),
.C(n_100),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_191),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g238 ( 
.A1(n_195),
.A2(n_203),
.B1(n_214),
.B2(n_215),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_157),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_205),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_163),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_151),
.B1(n_144),
.B2(n_143),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_204),
.B(n_207),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_143),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_135),
.B1(n_146),
.B2(n_104),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_213),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_7),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_13),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_166),
.A2(n_146),
.B1(n_8),
.B2(n_9),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_184),
.A2(n_146),
.B1(n_9),
.B2(n_11),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_161),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_194),
.B(n_172),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_222),
.B(n_223),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_165),
.C(n_162),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_242),
.C(n_199),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_236),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_232),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_161),
.B(n_162),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_239),
.B(n_240),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_172),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_237),
.Y(n_261)
);

A2O1A1O1Ixp25_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_183),
.B(n_177),
.C(n_190),
.D(n_189),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_204),
.B(n_212),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_241),
.A2(n_205),
.B(n_193),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_173),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_192),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_251),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_SL g272 ( 
.A(n_254),
.B(n_238),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_214),
.C(n_196),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_256),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_196),
.C(n_200),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_197),
.C(n_216),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_258),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_213),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_244),
.B1(n_248),
.B2(n_222),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_208),
.B1(n_193),
.B2(n_195),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_226),
.B1(n_203),
.B2(n_238),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_243),
.B(n_230),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_263),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_243),
.B(n_240),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_255),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_267),
.B1(n_270),
.B2(n_271),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_257),
.B1(n_226),
.B2(n_223),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_269),
.B(n_274),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_238),
.B1(n_237),
.B2(n_221),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_250),
.A2(n_238),
.B1(n_239),
.B2(n_227),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_260),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_254),
.A2(n_233),
.B(n_234),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_273),
.A2(n_275),
.B(n_261),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_202),
.B1(n_206),
.B2(n_201),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_261),
.A2(n_235),
.B(n_206),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_256),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_245),
.C(n_251),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_282),
.C(n_285),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_244),
.C(n_257),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_258),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_271),
.B(n_249),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_287),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_264),
.B(n_215),
.CI(n_247),
.CON(n_287),
.SN(n_287)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_269),
.B1(n_253),
.B2(n_270),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_291),
.A2(n_284),
.B1(n_283),
.B2(n_277),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_262),
.C(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_263),
.C(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_275),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_287),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_287),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_302),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_279),
.B(n_272),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_SL g303 ( 
.A(n_301),
.B(n_289),
.C(n_294),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_304),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_288),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_288),
.C(n_285),
.Y(n_305)
);

AOI31xp33_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_276),
.A3(n_174),
.B(n_16),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_308),
.A2(n_310),
.B1(n_306),
.B2(n_16),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_311),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_309),
.B1(n_14),
.B2(n_17),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_17),
.Y(n_314)
);


endmodule