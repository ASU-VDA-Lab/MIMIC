module fake_jpeg_5402_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_59),
.B1(n_71),
.B2(n_30),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

CKINVDCx6p67_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_87),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_46),
.B1(n_30),
.B2(n_36),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_86),
.B1(n_89),
.B2(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_92),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_69),
.B1(n_64),
.B2(n_74),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_28),
.B(n_20),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_94),
.CI(n_24),
.CON(n_112),
.SN(n_112)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_40),
.B1(n_28),
.B2(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_28),
.B1(n_34),
.B2(n_23),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_28),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_17),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_19),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_19),
.B1(n_34),
.B2(n_23),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_21),
.Y(n_130)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_104),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_80),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_103),
.A2(n_116),
.B1(n_118),
.B2(n_123),
.Y(n_152)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_107),
.B(n_112),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_58),
.C(n_39),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_124),
.C(n_96),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_17),
.B(n_25),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_20),
.Y(n_155)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_29),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_120),
.B1(n_129),
.B2(n_111),
.Y(n_132)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_39),
.C(n_36),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_98),
.B(n_29),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_105),
.B1(n_114),
.B2(n_116),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_69),
.B1(n_49),
.B2(n_74),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_138),
.B1(n_147),
.B2(n_154),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_49),
.B1(n_73),
.B2(n_54),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_139),
.B1(n_142),
.B2(n_126),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_95),
.B1(n_50),
.B2(n_62),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_61),
.B1(n_75),
.B2(n_90),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_61),
.B1(n_90),
.B2(n_88),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_36),
.B(n_39),
.C(n_22),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_26),
.B(n_32),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_82),
.B1(n_88),
.B2(n_77),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_77),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_106),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_32),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_96),
.B1(n_79),
.B2(n_26),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_117),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_160),
.B(n_182),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_183),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_178),
.B1(n_175),
.B2(n_176),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_133),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_156),
.C(n_157),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_112),
.B1(n_79),
.B2(n_121),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_167),
.B1(n_172),
.B2(n_24),
.Y(n_210)
);

XOR2x2_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_108),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_24),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_144),
.B1(n_142),
.B2(n_141),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_177),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_123),
.B1(n_118),
.B2(n_27),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_171),
.B(n_176),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_178),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_34),
.B(n_19),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_140),
.B(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_19),
.B1(n_26),
.B2(n_23),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_179),
.A2(n_127),
.B1(n_91),
.B2(n_32),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_184),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_131),
.B1(n_143),
.B2(n_149),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_137),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_151),
.A2(n_24),
.B(n_1),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_146),
.B(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_196),
.C(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_194),
.B(n_195),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_146),
.C(n_157),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_206),
.B(n_174),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_201),
.B(n_209),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_202),
.A2(n_213),
.B1(n_214),
.B2(n_171),
.Y(n_220)
);

AOI22x1_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_143),
.B1(n_131),
.B2(n_22),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_203),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_166),
.B1(n_161),
.B2(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_134),
.C(n_148),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_143),
.B(n_158),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_215),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

AOI22x1_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_91),
.B1(n_32),
.B2(n_22),
.Y(n_213)
);

AOI22x1_ASAP7_75t_L g214 ( 
.A1(n_161),
.A2(n_32),
.B1(n_22),
.B2(n_24),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_195),
.B(n_163),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_225),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_191),
.B(n_212),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_208),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_221),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_198),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_183),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_227),
.B(n_228),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_177),
.B(n_185),
.Y(n_227)
);

AOI21x1_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_162),
.B(n_24),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_192),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_145),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_236),
.C(n_240),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_173),
.B1(n_22),
.B2(n_145),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_237),
.B1(n_241),
.B2(n_4),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_145),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_193),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_199),
.B1(n_209),
.B2(n_194),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_189),
.B(n_0),
.C(n_2),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_255),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_230),
.A2(n_188),
.B1(n_214),
.B2(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_196),
.C(n_207),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_231),
.C(n_223),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_206),
.B(n_213),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_265),
.B(n_228),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_200),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_210),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_261),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_214),
.B1(n_211),
.B2(n_6),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_241),
.B1(n_237),
.B2(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_263),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_262),
.B1(n_260),
.B2(n_244),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_15),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_217),
.Y(n_267)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_257),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_221),
.A2(n_4),
.B(n_5),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_269),
.C(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_231),
.C(n_236),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_254),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_248),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_229),
.C(n_233),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_216),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_246),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_251),
.B1(n_8),
.B2(n_9),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_253),
.A2(n_226),
.B(n_242),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_277),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_240),
.C(n_239),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_278),
.C(n_247),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_7),
.C(n_8),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_7),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_282),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_7),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_288),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_249),
.B1(n_250),
.B2(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_290),
.A2(n_294),
.B(n_285),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_294),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_261),
.CI(n_265),
.CON(n_292),
.SN(n_292)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_292),
.B(n_297),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_7),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_8),
.C(n_10),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_8),
.Y(n_299)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_293),
.C(n_278),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_10),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_282),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_283),
.B1(n_268),
.B2(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_286),
.A2(n_275),
.B1(n_276),
.B2(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_281),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_311),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_11),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_11),
.Y(n_318)
);

INVx11_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_287),
.B1(n_279),
.B2(n_293),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_287),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_304),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_316),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_324),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_320),
.A2(n_323),
.B(n_314),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_11),
.C(n_12),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_302),
.B(n_13),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_326),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_322),
.B(n_305),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_308),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_303),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_330),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_319),
.B(n_301),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_320),
.B(n_307),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_333),
.A2(n_336),
.B(n_317),
.Y(n_338)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_321),
.B(n_306),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_339),
.B(n_334),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_337),
.B(n_313),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_335),
.B(n_331),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_304),
.C(n_331),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_13),
.B(n_14),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_14),
.B(n_331),
.Y(n_344)
);


endmodule