module fake_netlist_1_9373_n_864 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_864);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_864;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_227;
wire n_384;
wire n_617;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_695;
wire n_650;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_18), .Y(n_111) );
BUFx10_ASAP7_75t_L g112 ( .A(n_82), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_13), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_58), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_34), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_86), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_91), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_42), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_39), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_19), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_60), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_27), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_4), .Y(n_123) );
CKINVDCx14_ASAP7_75t_R g124 ( .A(n_37), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_54), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_90), .Y(n_126) );
INVxp67_ASAP7_75t_SL g127 ( .A(n_64), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_70), .Y(n_128) );
INVxp33_ASAP7_75t_SL g129 ( .A(n_6), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_5), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_100), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_101), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_88), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_77), .Y(n_134) );
BUFx10_ASAP7_75t_L g135 ( .A(n_9), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_48), .Y(n_136) );
INVxp67_ASAP7_75t_SL g137 ( .A(n_38), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_106), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_66), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_50), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_13), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_102), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_93), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g144 ( .A(n_9), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_61), .Y(n_146) );
INVx1_ASAP7_75t_SL g147 ( .A(n_22), .Y(n_147) );
INVxp33_ASAP7_75t_SL g148 ( .A(n_67), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_73), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_45), .Y(n_151) );
INVx1_ASAP7_75t_SL g152 ( .A(n_11), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_32), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_59), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_112), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_121), .B(n_0), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_120), .B(n_0), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_145), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_144), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_118), .Y(n_162) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_125), .A2(n_51), .B(n_109), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_130), .B(n_1), .Y(n_164) );
BUFx12f_ASAP7_75t_L g165 ( .A(n_112), .Y(n_165) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_116), .B(n_25), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_134), .Y(n_167) );
AND2x6_ASAP7_75t_L g168 ( .A(n_138), .B(n_26), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
AOI22xp5_ASAP7_75t_SL g170 ( .A1(n_141), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_149), .A2(n_2), .B(n_3), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_124), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_129), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_112), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_168), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_155), .B(n_117), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_168), .A2(n_148), .B1(n_135), .B2(n_111), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_173), .B(n_116), .Y(n_182) );
INVxp67_ASAP7_75t_SL g183 ( .A(n_173), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_168), .A2(n_135), .B1(n_123), .B2(n_111), .Y(n_185) );
AOI22xp33_ASAP7_75t_SL g186 ( .A1(n_170), .A2(n_123), .B1(n_114), .B2(n_135), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
INVx1_ASAP7_75t_SL g188 ( .A(n_173), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_155), .B(n_119), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_165), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_159), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_155), .B(n_119), .Y(n_195) );
BUFx10_ASAP7_75t_L g196 ( .A(n_177), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_165), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_155), .B(n_122), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_155), .B(n_122), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_176), .A2(n_113), .B1(n_147), .B2(n_152), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_162), .B(n_132), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_168), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_163), .A2(n_127), .B(n_137), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_177), .B(n_132), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_171), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_171), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_171), .Y(n_209) );
BUFx4f_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_172), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_162), .B(n_133), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_165), .B(n_133), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_176), .A2(n_154), .B1(n_153), .B2(n_146), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_172), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_172), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_169), .B(n_136), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_169), .B(n_136), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_172), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_172), .Y(n_222) );
INVx5_ASAP7_75t_L g223 ( .A(n_168), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_182), .B(n_175), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_201), .B(n_156), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_188), .A2(n_156), .B1(n_166), .B2(n_175), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_188), .B(n_157), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_201), .B(n_161), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_208), .Y(n_229) );
INVxp67_ASAP7_75t_L g230 ( .A(n_191), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_213), .A2(n_174), .B1(n_161), .B2(n_168), .Y(n_231) );
NOR3xp33_ASAP7_75t_L g232 ( .A(n_186), .B(n_157), .C(n_164), .Y(n_232) );
AOI22xp33_ASAP7_75t_SL g233 ( .A1(n_191), .A2(n_170), .B1(n_160), .B2(n_166), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_208), .Y(n_234) );
OR2x6_ASAP7_75t_SL g235 ( .A(n_197), .B(n_160), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_195), .B(n_161), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_209), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g238 ( .A(n_178), .B(n_168), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_183), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_195), .B(n_161), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_199), .B(n_164), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_178), .B(n_174), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_199), .B(n_174), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_178), .B(n_174), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_209), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_211), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_211), .A2(n_163), .B(n_167), .C(n_146), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_181), .A2(n_168), .B1(n_167), .B2(n_154), .Y(n_249) );
AND2x6_ASAP7_75t_SL g250 ( .A(n_215), .B(n_7), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_196), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_213), .A2(n_167), .B(n_139), .C(n_153), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_214), .B(n_139), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_206), .B(n_142), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_207), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_217), .A2(n_218), .B(n_222), .C(n_221), .Y(n_256) );
NOR3x1_ASAP7_75t_L g257 ( .A(n_200), .B(n_7), .C(n_8), .Y(n_257) );
OAI22xp5_ASAP7_75t_SL g258 ( .A1(n_216), .A2(n_142), .B1(n_128), .B2(n_131), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_198), .B(n_126), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_187), .Y(n_260) );
AND2x6_ASAP7_75t_SL g261 ( .A(n_200), .B(n_8), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_220), .B(n_168), .Y(n_262) );
AND2x6_ASAP7_75t_SL g263 ( .A(n_180), .B(n_10), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_217), .A2(n_57), .B(n_108), .Y(n_264) );
NOR2xp33_ASAP7_75t_SL g265 ( .A(n_178), .B(n_10), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_219), .B(n_56), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_218), .A2(n_11), .B1(n_12), .B2(n_14), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_190), .B(n_12), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_187), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_196), .B(n_63), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_203), .B(n_62), .Y(n_271) );
NOR2xp67_ASAP7_75t_L g272 ( .A(n_216), .B(n_14), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_193), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_196), .Y(n_274) );
NOR2xp33_ASAP7_75t_SL g275 ( .A(n_203), .B(n_15), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_196), .B(n_203), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_207), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_185), .B(n_15), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_203), .B(n_68), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_223), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_192), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_204), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_210), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_193), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_179), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_252), .A2(n_222), .B(n_221), .C(n_202), .Y(n_286) );
OAI21xp33_ASAP7_75t_L g287 ( .A1(n_241), .A2(n_212), .B(n_202), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_241), .B(n_204), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_225), .A2(n_210), .B1(n_212), .B2(n_223), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_251), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_256), .A2(n_210), .B(n_212), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_227), .Y(n_292) );
NOR2xp33_ASAP7_75t_R g293 ( .A(n_230), .B(n_210), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_227), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_285), .Y(n_295) );
INVx4_ASAP7_75t_L g296 ( .A(n_251), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_274), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_239), .B(n_204), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_260), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_232), .A2(n_204), .B1(n_212), .B2(n_205), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_239), .B(n_223), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_269), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_256), .A2(n_223), .B(n_192), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_274), .B(n_223), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_226), .A2(n_223), .B1(n_192), .B2(n_194), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_273), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_238), .B(n_192), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_224), .B(n_194), .Y(n_308) );
INVx5_ASAP7_75t_L g309 ( .A(n_285), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_236), .B(n_194), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
OAI21xp33_ASAP7_75t_L g312 ( .A1(n_240), .A2(n_189), .B(n_184), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_244), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_229), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_243), .A2(n_189), .B(n_184), .C(n_179), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_244), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_262), .A2(n_192), .B(n_205), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_242), .A2(n_192), .B(n_205), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_255), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_253), .B(n_189), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_228), .A2(n_184), .B(n_179), .C(n_205), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_258), .B(n_16), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_252), .B(n_17), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
OR2x6_ASAP7_75t_L g325 ( .A(n_272), .B(n_19), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_242), .A2(n_71), .B(n_107), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_245), .A2(n_69), .B(n_105), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_282), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_245), .A2(n_65), .B(n_104), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_276), .A2(n_55), .B(n_103), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_249), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_234), .B(n_20), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_SL g333 ( .A1(n_248), .A2(n_72), .B(n_99), .C(n_96), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_237), .B(n_21), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_246), .B(n_247), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_248), .A2(n_53), .B(n_95), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_281), .A2(n_52), .B(n_94), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_318), .A2(n_264), .B(n_271), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_292), .B(n_235), .Y(n_339) );
BUFx10_ASAP7_75t_L g340 ( .A(n_334), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_317), .A2(n_279), .B(n_271), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_321), .A2(n_231), .B(n_268), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_335), .A2(n_283), .B1(n_233), .B2(n_267), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_294), .B(n_235), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_300), .A2(n_291), .B(n_286), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_300), .A2(n_277), .B(n_255), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_334), .A2(n_254), .B1(n_275), .B2(n_265), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_309), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_303), .A2(n_279), .B(n_277), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_328), .B(n_263), .Y(n_350) );
BUFx2_ASAP7_75t_R g351 ( .A(n_323), .Y(n_351) );
OAI22x1_ASAP7_75t_L g352 ( .A1(n_322), .A2(n_257), .B1(n_261), .B2(n_250), .Y(n_352) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_287), .A2(n_314), .B(n_332), .C(n_302), .Y(n_353) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_290), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_288), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_287), .A2(n_278), .B(n_266), .C(n_270), .Y(n_356) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_331), .A2(n_259), .B(n_280), .C(n_24), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_296), .B(n_280), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_325), .Y(n_359) );
AOI21x1_ASAP7_75t_L g360 ( .A1(n_307), .A2(n_281), .B(n_74), .Y(n_360) );
OAI221xp5_ASAP7_75t_L g361 ( .A1(n_325), .A2(n_281), .B1(n_24), .B2(n_23), .C(n_29), .Y(n_361) );
OAI21xp33_ASAP7_75t_L g362 ( .A1(n_320), .A2(n_308), .B(n_312), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_305), .A2(n_75), .B(n_28), .Y(n_363) );
INVx3_ASAP7_75t_SL g364 ( .A(n_296), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_315), .A2(n_76), .B(n_30), .Y(n_365) );
NAND2x1_ASAP7_75t_L g366 ( .A(n_290), .B(n_78), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_336), .A2(n_49), .B(n_31), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_290), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_297), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g370 ( .A1(n_314), .A2(n_23), .B(n_33), .C(n_35), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_355), .B(n_299), .Y(n_371) );
OAI21x1_ASAP7_75t_SL g372 ( .A1(n_346), .A2(n_330), .B(n_326), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_355), .B(n_311), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_353), .Y(n_374) );
OAI21x1_ASAP7_75t_SL g375 ( .A1(n_365), .A2(n_329), .B(n_327), .Y(n_375) );
AO31x2_ASAP7_75t_L g376 ( .A1(n_356), .A2(n_306), .A3(n_337), .B(n_289), .Y(n_376) );
NOR2x1_ASAP7_75t_R g377 ( .A(n_359), .B(n_309), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_349), .Y(n_378) );
OA21x2_ASAP7_75t_L g379 ( .A1(n_345), .A2(n_295), .B(n_313), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_340), .B(n_309), .Y(n_380) );
AO31x2_ASAP7_75t_L g381 ( .A1(n_363), .A2(n_316), .A3(n_319), .B(n_310), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_369), .Y(n_382) );
OA21x2_ASAP7_75t_L g383 ( .A1(n_338), .A2(n_333), .B(n_298), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_369), .Y(n_384) );
AO21x2_ASAP7_75t_L g385 ( .A1(n_342), .A2(n_301), .B(n_293), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_362), .Y(n_386) );
NAND2x1_ASAP7_75t_L g387 ( .A(n_368), .B(n_324), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_343), .B(n_325), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_344), .B(n_328), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_370), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_340), .B(n_297), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_339), .B(n_304), .Y(n_392) );
OAI21x1_ASAP7_75t_L g393 ( .A1(n_360), .A2(n_324), .B(n_304), .Y(n_393) );
BUFx12f_ASAP7_75t_L g394 ( .A(n_348), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_341), .A2(n_324), .B(n_40), .Y(n_395) );
AO31x2_ASAP7_75t_L g396 ( .A1(n_363), .A2(n_36), .A3(n_41), .B(n_43), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_367), .A2(n_44), .B(n_46), .Y(n_397) );
AOI21x1_ASAP7_75t_L g398 ( .A1(n_367), .A2(n_47), .B(n_79), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_347), .A2(n_80), .B(n_81), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_374), .Y(n_400) );
AO21x2_ASAP7_75t_L g401 ( .A1(n_395), .A2(n_357), .B(n_361), .Y(n_401) );
NAND2xp33_ASAP7_75t_SL g402 ( .A(n_388), .B(n_364), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_388), .B(n_354), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_374), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_390), .B(n_357), .Y(n_405) );
AO21x2_ASAP7_75t_L g406 ( .A1(n_395), .A2(n_354), .B(n_358), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_372), .A2(n_358), .B(n_350), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_378), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
AO21x2_ASAP7_75t_L g410 ( .A1(n_372), .A2(n_366), .B(n_352), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_386), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_386), .Y(n_412) );
AO21x2_ASAP7_75t_L g413 ( .A1(n_375), .A2(n_390), .B(n_378), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_394), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_373), .A2(n_364), .B1(n_368), .B2(n_351), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_379), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_373), .B(n_83), .Y(n_419) );
AO21x1_ASAP7_75t_SL g420 ( .A1(n_382), .A2(n_84), .B(n_85), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_376), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_375), .A2(n_87), .B(n_89), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_396), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_396), .Y(n_425) );
AOI21xp5_ASAP7_75t_SL g426 ( .A1(n_377), .A2(n_92), .B(n_110), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_387), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_396), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_376), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_396), .B(n_381), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_377), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_387), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_382), .Y(n_433) );
OA21x2_ASAP7_75t_L g434 ( .A1(n_393), .A2(n_397), .B(n_398), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
OA21x2_ASAP7_75t_L g436 ( .A1(n_393), .A2(n_397), .B(n_398), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_381), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_381), .Y(n_439) );
BUFx12f_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_376), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_381), .B(n_376), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_437), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_403), .B(n_371), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_400), .B(n_384), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_408), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_411), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_402), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_442), .B(n_376), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_442), .B(n_376), .Y(n_450) );
NOR2x1_ASAP7_75t_SL g451 ( .A(n_420), .B(n_384), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_441), .B(n_381), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_440), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_432), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_407), .B(n_381), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_442), .B(n_383), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_407), .B(n_385), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_411), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_403), .B(n_389), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_432), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_437), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_439), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_403), .B(n_385), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_400), .B(n_385), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_432), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_432), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_402), .A2(n_392), .B1(n_394), .B2(n_391), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_403), .B(n_380), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_442), .B(n_430), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_432), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_430), .B(n_383), .Y(n_471) );
INVx2_ASAP7_75t_R g472 ( .A(n_414), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_430), .B(n_383), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_408), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_430), .B(n_383), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_441), .B(n_399), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_412), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_408), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_440), .Y(n_479) );
NAND2x1_ASAP7_75t_L g480 ( .A(n_432), .B(n_391), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_441), .B(n_435), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_441), .B(n_435), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_412), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_441), .B(n_435), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_424), .B(n_425), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_424), .B(n_425), .Y(n_486) );
NOR2xp67_ASAP7_75t_L g487 ( .A(n_424), .B(n_438), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_408), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_408), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_427), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_413), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_412), .B(n_400), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_416), .A2(n_419), .B1(n_407), .B2(n_401), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_425), .B(n_438), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_428), .B(n_438), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_428), .B(n_429), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_428), .B(n_429), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_404), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_427), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_404), .B(n_405), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_404), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_414), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_422), .B(n_429), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_414), .Y(n_504) );
BUFx3_ASAP7_75t_L g505 ( .A(n_440), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_407), .B(n_427), .Y(n_506) );
INVx3_ASAP7_75t_SL g507 ( .A(n_415), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_405), .B(n_433), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_469), .B(n_422), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_469), .B(n_422), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_467), .A2(n_416), .B1(n_440), .B2(n_415), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_446), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_444), .B(n_419), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_453), .B(n_479), .Y(n_514) );
BUFx2_ASAP7_75t_L g515 ( .A(n_448), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_444), .B(n_419), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_469), .B(n_422), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_449), .B(n_407), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_449), .B(n_407), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_443), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_449), .B(n_439), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_453), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_459), .B(n_419), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_493), .A2(n_431), .B1(n_401), .B2(n_433), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_450), .B(n_413), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_450), .B(n_413), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_459), .B(n_433), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_453), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_447), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_458), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_446), .Y(n_531) );
INVxp67_ASAP7_75t_SL g532 ( .A(n_443), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_450), .B(n_413), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_485), .B(n_433), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_481), .B(n_413), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_458), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_477), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_481), .B(n_413), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_481), .B(n_417), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_477), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_446), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_463), .B(n_417), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_485), .B(n_401), .Y(n_543) );
BUFx3_ASAP7_75t_L g544 ( .A(n_479), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_461), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_482), .B(n_484), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_482), .B(n_417), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_482), .B(n_417), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_484), .B(n_417), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_463), .B(n_421), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_485), .B(n_401), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_474), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_461), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_484), .B(n_418), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_506), .B(n_427), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_483), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_486), .B(n_401), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_486), .B(n_421), .Y(n_558) );
AND2x4_ASAP7_75t_SL g559 ( .A(n_462), .B(n_409), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_506), .B(n_410), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_486), .B(n_418), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_474), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_462), .B(n_418), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_490), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_494), .B(n_418), .Y(n_565) );
INVx4_ASAP7_75t_L g566 ( .A(n_479), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_483), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_494), .B(n_418), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_474), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_492), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_506), .B(n_410), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_506), .B(n_410), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_492), .Y(n_573) );
INVxp33_ASAP7_75t_L g574 ( .A(n_480), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_466), .B(n_410), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_502), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_502), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_478), .Y(n_578) );
BUFx3_ASAP7_75t_L g579 ( .A(n_505), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_466), .B(n_410), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_490), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_494), .B(n_401), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_495), .B(n_421), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_495), .B(n_421), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_495), .B(n_421), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_504), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_504), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_456), .B(n_473), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_456), .B(n_473), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_468), .B(n_410), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_456), .B(n_406), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_468), .B(n_423), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_466), .B(n_406), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_498), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_501), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_478), .Y(n_596) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_505), .B(n_426), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_471), .B(n_406), .Y(n_598) );
AND2x4_ASAP7_75t_SL g599 ( .A(n_454), .B(n_426), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_471), .B(n_406), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_501), .B(n_423), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_471), .B(n_406), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_496), .B(n_423), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_586), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_586), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_570), .B(n_497), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_512), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_587), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_566), .B(n_522), .Y(n_609) );
INVx2_ASAP7_75t_SL g610 ( .A(n_559), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g611 ( .A(n_566), .B(n_505), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_588), .B(n_475), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_587), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_536), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_536), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_588), .B(n_475), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_512), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_537), .Y(n_618) );
BUFx2_ASAP7_75t_L g619 ( .A(n_566), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_537), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_520), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_545), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_589), .B(n_475), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_589), .B(n_508), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_531), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_525), .B(n_473), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_573), .B(n_496), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_531), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_521), .B(n_508), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_521), .B(n_497), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_509), .B(n_497), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_546), .B(n_489), .Y(n_632) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_553), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_555), .B(n_487), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_540), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_540), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_509), .B(n_496), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_546), .B(n_478), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_510), .B(n_503), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_510), .B(n_503), .Y(n_640) );
OR2x6_ASAP7_75t_L g641 ( .A(n_514), .B(n_480), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_529), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_517), .B(n_503), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_517), .B(n_490), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_541), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_539), .B(n_499), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_544), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_541), .Y(n_648) );
BUFx2_ASAP7_75t_L g649 ( .A(n_544), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_539), .B(n_499), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_527), .B(n_500), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_534), .B(n_547), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_547), .B(n_499), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_518), .B(n_519), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_548), .B(n_452), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_549), .B(n_452), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_525), .B(n_452), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_530), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_556), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_579), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_518), .B(n_500), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_567), .Y(n_662) );
NOR2x1_ASAP7_75t_SL g663 ( .A(n_579), .B(n_420), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_526), .B(n_452), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_559), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_555), .Y(n_666) );
INVx2_ASAP7_75t_SL g667 ( .A(n_522), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_526), .B(n_452), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_552), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_519), .B(n_445), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_533), .B(n_457), .Y(n_671) );
NAND2x1p5_ASAP7_75t_L g672 ( .A(n_597), .B(n_511), .Y(n_672) );
NOR2xp67_ASAP7_75t_L g673 ( .A(n_528), .B(n_455), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_594), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_595), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_552), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_576), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_577), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_533), .B(n_457), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_532), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_558), .B(n_445), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_558), .B(n_464), .Y(n_682) );
AND2x4_ASAP7_75t_SL g683 ( .A(n_555), .B(n_465), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_535), .B(n_457), .Y(n_684) );
OAI32xp33_ASAP7_75t_L g685 ( .A1(n_514), .A2(n_507), .A3(n_465), .B1(n_454), .B2(n_460), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_561), .B(n_464), .Y(n_686) );
NAND2x1_ASAP7_75t_SL g687 ( .A(n_560), .B(n_507), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_565), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_535), .B(n_457), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_562), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_538), .B(n_455), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_568), .B(n_487), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_538), .B(n_455), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_591), .B(n_455), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_591), .B(n_472), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_568), .B(n_488), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_554), .B(n_470), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_554), .B(n_585), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_598), .B(n_472), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_612), .B(n_585), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_622), .B(n_600), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_619), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_632), .B(n_550), .Y(n_703) );
OR2x2_ASAP7_75t_L g704 ( .A(n_638), .B(n_550), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_612), .B(n_584), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_624), .B(n_542), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_616), .B(n_584), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_621), .A2(n_515), .B1(n_524), .B2(n_590), .C(n_543), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g709 ( .A1(n_672), .A2(n_574), .B(n_514), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_641), .A2(n_523), .B1(n_516), .B2(n_513), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_654), .B(n_626), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_631), .B(n_542), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_642), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_658), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_637), .B(n_652), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_659), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_649), .Y(n_717) );
OR2x2_ASAP7_75t_L g718 ( .A(n_639), .B(n_583), .Y(n_718) );
OR2x2_ASAP7_75t_L g719 ( .A(n_640), .B(n_643), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_623), .B(n_602), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_623), .B(n_602), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_698), .B(n_600), .Y(n_722) );
INVxp33_ASAP7_75t_L g723 ( .A(n_611), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_694), .B(n_515), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_662), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_661), .B(n_551), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_694), .B(n_564), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_630), .B(n_563), .Y(n_728) );
O2A1O1Ixp33_ASAP7_75t_SL g729 ( .A1(n_609), .A2(n_647), .B(n_660), .C(n_665), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_674), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_675), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_641), .A2(n_557), .B1(n_582), .B2(n_599), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_677), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_626), .B(n_629), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_678), .Y(n_735) );
NOR2x1p5_ASAP7_75t_SL g736 ( .A(n_680), .B(n_563), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_633), .B(n_601), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_611), .B(n_581), .Y(n_738) );
OAI21xp33_ASAP7_75t_L g739 ( .A1(n_672), .A2(n_560), .B(n_571), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_657), .B(n_581), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_670), .B(n_596), .Y(n_741) );
OAI21xp5_ASAP7_75t_SL g742 ( .A1(n_609), .A2(n_572), .B(n_571), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_651), .B(n_454), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_657), .B(n_560), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_664), .B(n_572), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g746 ( .A1(n_641), .A2(n_592), .B(n_470), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_688), .B(n_596), .Y(n_747) );
AND2x4_ASAP7_75t_L g748 ( .A(n_673), .B(n_571), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_682), .B(n_603), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_686), .B(n_578), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_667), .B(n_465), .Y(n_751) );
INVxp33_ASAP7_75t_L g752 ( .A(n_663), .Y(n_752) );
AO21x1_ASAP7_75t_L g753 ( .A1(n_634), .A2(n_580), .B(n_575), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_667), .Y(n_754) );
NOR3xp33_ASAP7_75t_L g755 ( .A(n_685), .B(n_460), .C(n_454), .Y(n_755) );
NOR2x1_ASAP7_75t_L g756 ( .A(n_634), .B(n_465), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_607), .Y(n_757) );
OR2x2_ASAP7_75t_L g758 ( .A(n_681), .B(n_578), .Y(n_758) );
INVx2_ASAP7_75t_SL g759 ( .A(n_610), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_664), .B(n_572), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_604), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_605), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_608), .Y(n_763) );
OAI21xp33_ASAP7_75t_L g764 ( .A1(n_687), .A2(n_593), .B(n_580), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_665), .A2(n_593), .B1(n_476), .B2(n_423), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_668), .B(n_580), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_696), .B(n_569), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_613), .Y(n_768) );
OAI21xp33_ASAP7_75t_L g769 ( .A1(n_736), .A2(n_693), .B(n_691), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_744), .B(n_671), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_729), .A2(n_699), .B(n_695), .Y(n_771) );
NAND3xp33_ASAP7_75t_SL g772 ( .A(n_709), .B(n_695), .C(n_699), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_703), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_743), .A2(n_666), .B1(n_679), .B2(n_671), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_726), .B(n_684), .Y(n_775) );
NAND3xp33_ASAP7_75t_SL g776 ( .A(n_753), .B(n_692), .C(n_644), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_704), .Y(n_777) );
INVxp67_ASAP7_75t_L g778 ( .A(n_759), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_745), .B(n_689), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_752), .B(n_634), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_715), .B(n_606), .Y(n_781) );
AOI21xp33_ASAP7_75t_SL g782 ( .A1(n_739), .A2(n_666), .B(n_646), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_757), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_701), .B(n_627), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_723), .A2(n_684), .B1(n_653), .B2(n_650), .Y(n_785) );
OAI21xp33_ASAP7_75t_L g786 ( .A1(n_739), .A2(n_656), .B(n_655), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_760), .B(n_697), .Y(n_787) );
OAI222xp33_ASAP7_75t_L g788 ( .A1(n_738), .A2(n_618), .B1(n_614), .B2(n_615), .C1(n_620), .C2(n_636), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_737), .B(n_635), .Y(n_789) );
AOI221xp5_ASAP7_75t_L g790 ( .A1(n_708), .A2(n_593), .B1(n_575), .B2(n_491), .C(n_690), .Y(n_790) );
OR2x2_ASAP7_75t_L g791 ( .A(n_734), .B(n_690), .Y(n_791) );
OAI322xp33_ASAP7_75t_L g792 ( .A1(n_749), .A2(n_628), .A3(n_625), .B1(n_617), .B2(n_607), .C1(n_676), .C2(n_669), .Y(n_792) );
NAND4xp25_ASAP7_75t_SL g793 ( .A(n_732), .B(n_683), .C(n_476), .D(n_625), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_713), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_714), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_716), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_706), .Y(n_797) );
INVx2_ASAP7_75t_SL g798 ( .A(n_717), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_728), .B(n_676), .Y(n_799) );
OAI21xp5_ASAP7_75t_SL g800 ( .A1(n_742), .A2(n_476), .B(n_648), .Y(n_800) );
NOR4xp25_ASAP7_75t_L g801 ( .A(n_742), .B(n_491), .C(n_669), .D(n_617), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_725), .Y(n_802) );
INVx1_ASAP7_75t_SL g803 ( .A(n_702), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_737), .B(n_648), .Y(n_804) );
AOI32xp33_ASAP7_75t_L g805 ( .A1(n_724), .A2(n_645), .A3(n_628), .B1(n_569), .B2(n_488), .Y(n_805) );
INVxp67_ASAP7_75t_SL g806 ( .A(n_754), .Y(n_806) );
AOI221xp5_ASAP7_75t_L g807 ( .A1(n_776), .A2(n_730), .B1(n_735), .B2(n_733), .C(n_731), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g808 ( .A1(n_800), .A2(n_782), .B1(n_771), .B2(n_772), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_786), .A2(n_769), .B1(n_785), .B2(n_778), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_775), .B(n_711), .Y(n_810) );
OAI221xp5_ASAP7_75t_SL g811 ( .A1(n_801), .A2(n_710), .B1(n_764), .B2(n_765), .C(n_732), .Y(n_811) );
AOI22xp33_ASAP7_75t_SL g812 ( .A1(n_771), .A2(n_748), .B1(n_746), .B2(n_727), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_785), .A2(n_710), .B1(n_748), .B2(n_740), .Y(n_813) );
AOI21xp33_ASAP7_75t_L g814 ( .A1(n_790), .A2(n_751), .B(n_756), .Y(n_814) );
O2A1O1Ixp33_ASAP7_75t_SL g815 ( .A1(n_780), .A2(n_788), .B(n_803), .C(n_798), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_805), .A2(n_746), .B(n_765), .C(n_755), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_789), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_775), .B(n_719), .Y(n_818) );
AOI322xp5_ASAP7_75t_L g819 ( .A1(n_781), .A2(n_720), .A3(n_721), .B1(n_722), .B2(n_700), .C1(n_705), .C2(n_707), .Y(n_819) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_792), .A2(n_768), .B1(n_763), .B2(n_762), .C(n_761), .Y(n_820) );
OAI21xp33_ASAP7_75t_L g821 ( .A1(n_774), .A2(n_750), .B(n_741), .Y(n_821) );
OAI21xp5_ASAP7_75t_L g822 ( .A1(n_793), .A2(n_747), .B(n_741), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_804), .Y(n_823) );
OAI321xp33_ASAP7_75t_L g824 ( .A1(n_804), .A2(n_766), .A3(n_758), .B1(n_712), .B2(n_767), .C(n_718), .Y(n_824) );
NOR3x1_ASAP7_75t_L g825 ( .A(n_806), .B(n_451), .C(n_420), .Y(n_825) );
BUFx12f_ASAP7_75t_L g826 ( .A(n_791), .Y(n_826) );
INVx1_ASAP7_75t_SL g827 ( .A(n_803), .Y(n_827) );
AOI221xp5_ASAP7_75t_SL g828 ( .A1(n_797), .A2(n_434), .B1(n_436), .B2(n_773), .C(n_777), .Y(n_828) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_794), .A2(n_802), .B1(n_796), .B2(n_795), .C(n_784), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g830 ( .A(n_783), .B(n_799), .C(n_787), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_770), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_779), .A2(n_619), .B1(n_663), .B2(n_566), .Y(n_832) );
OAI21xp33_ASAP7_75t_SL g833 ( .A1(n_801), .A2(n_780), .B(n_771), .Y(n_833) );
NAND4xp25_ASAP7_75t_L g834 ( .A(n_790), .B(n_511), .C(n_709), .D(n_739), .Y(n_834) );
OAI21xp5_ASAP7_75t_L g835 ( .A1(n_776), .A2(n_729), .B(n_788), .Y(n_835) );
NAND2xp33_ASAP7_75t_L g836 ( .A(n_769), .B(n_752), .Y(n_836) );
INVxp67_ASAP7_75t_L g837 ( .A(n_827), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_817), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_819), .B(n_820), .Y(n_839) );
NAND3xp33_ASAP7_75t_L g840 ( .A(n_811), .B(n_833), .C(n_835), .Y(n_840) );
NOR5xp2_ASAP7_75t_L g841 ( .A(n_811), .B(n_824), .C(n_815), .D(n_829), .E(n_816), .Y(n_841) );
AND4x1_ASAP7_75t_L g842 ( .A(n_809), .B(n_807), .C(n_825), .D(n_813), .Y(n_842) );
CKINVDCx16_ASAP7_75t_R g843 ( .A(n_826), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_821), .B(n_830), .Y(n_844) );
NOR2xp67_ASAP7_75t_SL g845 ( .A(n_843), .B(n_834), .Y(n_845) );
NOR3xp33_ASAP7_75t_L g846 ( .A(n_840), .B(n_808), .C(n_836), .Y(n_846) );
NAND4xp75_ASAP7_75t_L g847 ( .A(n_839), .B(n_828), .C(n_814), .D(n_822), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_837), .Y(n_848) );
INVx2_ASAP7_75t_SL g849 ( .A(n_842), .Y(n_849) );
NAND3x1_ASAP7_75t_L g850 ( .A(n_846), .B(n_841), .C(n_844), .Y(n_850) );
INVxp67_ASAP7_75t_L g851 ( .A(n_845), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_848), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_852), .Y(n_853) );
OA22x2_ASAP7_75t_L g854 ( .A1(n_851), .A2(n_849), .B1(n_846), .B2(n_847), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_850), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_854), .A2(n_838), .B1(n_812), .B2(n_832), .Y(n_856) );
INVx4_ASAP7_75t_L g857 ( .A(n_855), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_857), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_856), .B(n_853), .Y(n_859) );
NAND3xp33_ASAP7_75t_L g860 ( .A(n_858), .B(n_853), .C(n_832), .Y(n_860) );
INVxp67_ASAP7_75t_SL g861 ( .A(n_859), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_861), .B(n_823), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_862), .B(n_860), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_863), .A2(n_818), .B1(n_831), .B2(n_810), .Y(n_864) );
endmodule