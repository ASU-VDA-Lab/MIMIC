module fake_jpeg_2074_n_113 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_16),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_36),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_55),
.B(n_29),
.Y(n_60)
);

BUFx24_ASAP7_75t_SL g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_65),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_31),
.B1(n_30),
.B2(n_36),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_59),
.B1(n_40),
.B2(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_38),
.B1(n_33),
.B2(n_34),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_14),
.Y(n_76)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_39),
.B(n_46),
.C(n_45),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_46),
.B(n_52),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_73),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_40),
.B1(n_29),
.B2(n_2),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_60),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_0),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_85),
.B1(n_23),
.B2(n_26),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_60),
.Y(n_79)
);

AOI221xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_87),
.B1(n_89),
.B2(n_72),
.C(n_8),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_4),
.B(n_5),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_11),
.B(n_12),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_7),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_19),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_22),
.B(n_27),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_97),
.B(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_25),
.C(n_17),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_80),
.B1(n_83),
.B2(n_12),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_96),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_97),
.C(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_103),
.B1(n_100),
.B2(n_106),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_94),
.Y(n_109)
);

OAI21x1_ASAP7_75t_SL g110 ( 
.A1(n_109),
.A2(n_101),
.B(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_104),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_92),
.C(n_28),
.Y(n_113)
);


endmodule