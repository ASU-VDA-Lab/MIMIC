module fake_jpeg_5437_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_265;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_26),
.B1(n_19),
.B2(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_14),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_20),
.B1(n_21),
.B2(n_41),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_44),
.B1(n_54),
.B2(n_58),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_20),
.B1(n_21),
.B2(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_30),
.B(n_22),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_33),
.Y(n_73)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_21),
.B1(n_29),
.B2(n_16),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_62),
.B1(n_17),
.B2(n_18),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_60),
.Y(n_81)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_33),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_37),
.C(n_35),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_80),
.Y(n_96)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_56),
.B1(n_49),
.B2(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_54),
.B1(n_17),
.B2(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_43),
.Y(n_90)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_35),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_15),
.B(n_28),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_47),
.B(n_46),
.C(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_84),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_54),
.B1(n_48),
.B2(n_57),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_101),
.B1(n_75),
.B2(n_64),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_82),
.B(n_79),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_69),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_49),
.B1(n_46),
.B2(n_55),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_71),
.B1(n_84),
.B2(n_78),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_57),
.B1(n_44),
.B2(n_60),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_22),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_68),
.B1(n_82),
.B2(n_74),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_88),
.B1(n_101),
.B2(n_91),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_115),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_66),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_127),
.C(n_125),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_65),
.B(n_99),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_120),
.B1(n_89),
.B2(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_121),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_73),
.B1(n_66),
.B2(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_124),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_67),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_73),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_127),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_93),
.B(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_72),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_129),
.A2(n_94),
.B(n_105),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_140),
.B1(n_130),
.B2(n_121),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_115),
.C(n_120),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_134),
.C(n_142),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_91),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_148),
.B(n_151),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_139),
.B1(n_114),
.B2(n_117),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_107),
.B(n_119),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_87),
.B(n_86),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_78),
.B(n_84),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_74),
.B1(n_90),
.B2(n_105),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_101),
.B1(n_91),
.B2(n_86),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_106),
.C(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_119),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_122),
.C(n_124),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_147),
.B(n_113),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_99),
.B(n_76),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_76),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_109),
.A2(n_85),
.B(n_81),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_38),
.C(n_83),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_111),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_159),
.A2(n_163),
.B1(n_168),
.B2(n_172),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_164),
.B(n_169),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_136),
.B1(n_180),
.B2(n_170),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_107),
.B1(n_126),
.B2(n_110),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_165),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_116),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_176),
.B1(n_180),
.B2(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_123),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_171),
.B(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_146),
.Y(n_174)
);

NAND4xp25_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_103),
.C(n_97),
.D(n_152),
.Y(n_186)
);

AO22x1_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_83),
.B1(n_31),
.B2(n_34),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_38),
.B(n_116),
.C(n_22),
.D(n_30),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_181),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_38),
.Y(n_181)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_188),
.A2(n_193),
.B1(n_195),
.B2(n_202),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_154),
.B1(n_145),
.B2(n_131),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_197),
.B1(n_199),
.B2(n_201),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_135),
.B1(n_176),
.B2(n_161),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_194),
.B1(n_203),
.B2(n_169),
.Y(n_214)
);

OAI21x1_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_148),
.B(n_137),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_140),
.B1(n_149),
.B2(n_155),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_159),
.A2(n_149),
.B1(n_144),
.B2(n_134),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_142),
.C(n_150),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_179),
.C(n_195),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_103),
.B1(n_97),
.B2(n_19),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_97),
.B1(n_26),
.B2(n_34),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_34),
.B1(n_32),
.B2(n_27),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_32),
.B1(n_27),
.B2(n_25),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_150),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_30),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_175),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_215),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_213),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_181),
.C(n_166),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_210),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_169),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_187),
.B(n_184),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_166),
.C(n_178),
.Y(n_210)
);

NOR4xp25_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_158),
.C(n_157),
.D(n_174),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_25),
.Y(n_241)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_222),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_32),
.C(n_30),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_220),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_30),
.C(n_27),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_30),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_0),
.Y(n_244)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_27),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_25),
.B1(n_23),
.B2(n_2),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_203),
.B1(n_202),
.B2(n_201),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_0),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_205),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_230),
.A2(n_231),
.B(n_232),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_187),
.B(n_184),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_189),
.B(n_182),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_209),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_199),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_239),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_214),
.A2(n_182),
.B1(n_189),
.B2(n_224),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_241),
.B1(n_219),
.B2(n_216),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_25),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_5),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_221),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_0),
.C(n_1),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_245),
.A2(n_14),
.B(n_7),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_208),
.C(n_207),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_248),
.C(n_240),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_210),
.C(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_254),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_209),
.B(n_2),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_6),
.B(n_7),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_260),
.B(n_6),
.Y(n_270)
);

OAI321xp33_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_4),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_237),
.B(n_5),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_258),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_5),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_262),
.B(n_266),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_252),
.A2(n_227),
.B1(n_233),
.B2(n_238),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_255),
.B1(n_248),
.B2(n_247),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_243),
.B(n_245),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_271),
.B(n_273),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_235),
.C(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_9),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_243),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_253),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_284),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_265),
.B(n_10),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_235),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_282),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_7),
.B(n_8),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_281),
.A2(n_9),
.B(n_11),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_8),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_8),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_277),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_272),
.A3(n_267),
.B1(n_268),
.B2(n_265),
.C1(n_273),
.C2(n_270),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_289),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_12),
.C(n_13),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_291),
.C(n_283),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_290),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.C(n_296),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_285),
.A2(n_278),
.B(n_275),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_285),
.C(n_13),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_295),
.C(n_13),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_298),
.Y(n_300)
);


endmodule