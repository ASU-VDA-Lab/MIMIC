module fake_jpeg_26800_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_62),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_0),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_47),
.B1(n_56),
.B2(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_71),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_47),
.B1(n_54),
.B2(n_45),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_76),
.B1(n_1),
.B2(n_2),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_49),
.B1(n_41),
.B2(n_46),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_76),
.B1(n_69),
.B2(n_77),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_75),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_57),
.B1(n_49),
.B2(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_50),
.B1(n_48),
.B2(n_42),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_94),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_18),
.B(n_38),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_100),
.B1(n_86),
.B2(n_87),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_103),
.B(n_8),
.C(n_9),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_6),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_26),
.B(n_33),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_107),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_110),
.B(n_111),
.Y(n_114)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_101),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_109),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_8),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_103),
.B(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_116),
.B1(n_91),
.B2(n_102),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_114),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_117),
.Y(n_121)
);

AOI31xp67_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_122),
.A3(n_115),
.B(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_121),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_9),
.B(n_10),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_10),
.B(n_11),
.C(n_13),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_19),
.C(n_24),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_102),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_28),
.B(n_29),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_31),
.Y(n_131)
);


endmodule