module fake_jpeg_30451_n_155 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_13),
.B(n_4),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_68),
.Y(n_76)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_1),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_54),
.B1(n_57),
.B2(n_46),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_84),
.B1(n_86),
.B2(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_79),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_59),
.B1(n_55),
.B2(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_58),
.B1(n_51),
.B2(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_45),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_59),
.B1(n_45),
.B2(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_62),
.B1(n_47),
.B2(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_95),
.B1(n_96),
.B2(n_101),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_18),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_11),
.C(n_12),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_6),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_44),
.B1(n_25),
.B2(n_26),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_7),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_20),
.B1(n_39),
.B2(n_37),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_8),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_10),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_10),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_114),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_116),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_28),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_99),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_11),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_43),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_14),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_88),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_36),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_128),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_132),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_15),
.C(n_16),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_17),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_27),
.C(n_33),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_112),
.B1(n_109),
.B2(n_115),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_126),
.C(n_130),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_106),
.B(n_118),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_133),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_141),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_134),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_137),
.B(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_129),
.B1(n_143),
.B2(n_138),
.Y(n_153)
);

OAI321xp33_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_145),
.A3(n_131),
.B1(n_115),
.B2(n_113),
.C(n_140),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_142),
.Y(n_155)
);


endmodule