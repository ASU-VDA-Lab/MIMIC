module fake_netlist_1_12353_n_28 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
NAND3xp33_ASAP7_75t_L g11 ( .A(n_10), .B(n_6), .C(n_9), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
INVx5_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
NOR2xp33_ASAP7_75t_R g14 ( .A(n_2), .B(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
AND3x1_ASAP7_75t_L g18 ( .A(n_12), .B(n_0), .C(n_2), .Y(n_18) );
OAI22xp5_ASAP7_75t_SL g19 ( .A1(n_18), .A2(n_16), .B1(n_13), .B2(n_11), .Y(n_19) );
NAND2xp33_ASAP7_75t_R g20 ( .A(n_17), .B(n_14), .Y(n_20) );
AOI221xp5_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_17), .B1(n_14), .B2(n_13), .C(n_3), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_13), .Y(n_22) );
AOI31xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_20), .A3(n_5), .B(n_4), .Y(n_23) );
NAND2xp33_ASAP7_75t_R g24 ( .A(n_23), .B(n_22), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_13), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AOI22xp33_ASAP7_75t_R g27 ( .A1(n_26), .A2(n_24), .B1(n_7), .B2(n_8), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
endmodule