module real_jpeg_23347_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_3),
.A2(n_31),
.B1(n_36),
.B2(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_3),
.A2(n_31),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_3),
.A2(n_31),
.B1(n_51),
.B2(n_52),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_5),
.A2(n_51),
.B1(n_52),
.B2(n_66),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_5),
.A2(n_36),
.B1(n_40),
.B2(n_66),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_66),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_24),
.B1(n_36),
.B2(n_40),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_10),
.A2(n_36),
.B1(n_40),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_10),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_43),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_10),
.A2(n_43),
.B1(n_64),
.B2(n_65),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_10),
.A2(n_62),
.B(n_125),
.C(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_10),
.B(n_60),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_10),
.A2(n_49),
.B(n_51),
.C(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_10),
.B(n_23),
.C(n_39),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_10),
.B(n_147),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_10),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_10),
.B(n_41),
.Y(n_221)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_11),
.B(n_204),
.Y(n_209)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_11),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_130),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_129),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_107),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_16),
.B(n_107),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_74),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_46),
.C(n_58),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_18),
.A2(n_19),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_20),
.B(n_32),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_27),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_21),
.A2(n_29),
.B(n_82),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_22),
.A2(n_23),
.B1(n_38),
.B2(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_23),
.B(n_215),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_25),
.B(n_30),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_25),
.A2(n_81),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_25),
.B(n_81),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_25),
.B(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_28),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_28),
.B(n_202),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_44),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_33),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_42),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_34),
.B(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_34),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_41),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_35)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_40),
.B1(n_49),
.B2(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_36),
.B(n_192),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_40),
.A2(n_43),
.B(n_54),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_41),
.B(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_42),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_43),
.A2(n_51),
.B(n_61),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_44),
.A2(n_85),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_44),
.B(n_178),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_46),
.A2(n_58),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_46),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_55),
.B(n_56),
.Y(n_46)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_47),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_47),
.B(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_55),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_48)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_52),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_55),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_55),
.B(n_56),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_55),
.Y(n_147)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_57),
.B(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_58),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_59),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_71),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_68),
.Y(n_92)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_68),
.B(n_91),
.Y(n_139)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_100),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_87),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_78),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_82),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_84),
.A2(n_105),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_84),
.B(n_142),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_86),
.B(n_189),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_119),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_98),
.B(n_146),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_101),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_101),
.A2(n_106),
.B1(n_173),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_114),
.C(n_128),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_108),
.A2(n_109),
.B1(n_128),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_114),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_123),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_127),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_128),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_166),
.B(n_242),
.C(n_247),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_154),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_132),
.B(n_154),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_150),
.B2(n_153),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_148),
.B2(n_149),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_135),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_135),
.B(n_149),
.C(n_153),
.Y(n_243)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_143),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_138),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.C(n_161),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_156),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_161),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_164),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_241),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_183),
.B(n_240),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_180),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_169),
.B(n_180),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_175),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_170),
.B(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_172),
.B(n_175),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_173),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_235),
.B(n_239),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_226),
.B(n_234),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_206),
.B(n_225),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_187),
.B(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_190),
.B1(n_191),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_200),
.B2(n_205),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_199),
.C(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_200),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_212),
.B(n_224),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_210),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_209),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_220),
.B(n_223),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_231),
.C(n_232),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_236),
.B(n_237),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);


endmodule