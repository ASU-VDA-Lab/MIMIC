module fake_ariane_1852_n_617 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_617);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_617;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_588;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_616;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_544;
wire n_216;
wire n_540;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_337;
wire n_437;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_292;
wire n_156;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_52),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_50),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_30),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_107),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_58),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_39),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_87),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_7),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_2),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_47),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_88),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_5),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_1),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_31),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_98),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_77),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_114),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_64),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_18),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_59),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_48),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_43),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_14),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_78),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_10),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_34),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_32),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_19),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_20),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_91),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_4),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_42),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_55),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_41),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_4),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_61),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_79),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_69),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_38),
.B(n_7),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_118),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_102),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_131),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_1),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_9),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_15),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_70),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_33),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_40),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_3),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_71),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_80),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_27),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_82),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_21),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_94),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_106),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

OAI21x1_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_73),
.B(n_134),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

OA21x2_ASAP7_75t_L g209 ( 
.A1(n_137),
.A2(n_0),
.B(n_2),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_138),
.A2(n_0),
.B(n_3),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_12),
.Y(n_212)
);

OAI22x1_ASAP7_75t_R g213 ( 
.A1(n_169),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_141),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_153),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

OAI22x1_ASAP7_75t_R g226 ( 
.A1(n_189),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_226)
);

AOI22x1_ASAP7_75t_SL g227 ( 
.A1(n_145),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_164),
.B(n_11),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_168),
.B(n_16),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_170),
.B(n_17),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_22),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_146),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_158),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_136),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_182),
.B(n_26),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_161),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_143),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

INVxp33_ASAP7_75t_SL g246 ( 
.A(n_185),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_196),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_223),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_238),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_238),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_178),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_228),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_242),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_242),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_221),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_216),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_239),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_221),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_225),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_R g263 ( 
.A(n_212),
.B(n_140),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_218),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_206),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_220),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_206),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_220),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_223),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_204),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_223),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_223),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_224),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_224),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_224),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_233),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_245),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_237),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_227),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_204),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_214),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_R g292 ( 
.A(n_234),
.B(n_144),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_204),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_268),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_251),
.B(n_235),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_230),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_270),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_263),
.A2(n_210),
.B1(n_209),
.B2(n_241),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_231),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_282),
.B(n_240),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_232),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_207),
.B(n_244),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

BUFx8_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_214),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_247),
.B(n_197),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_285),
.B(n_292),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_258),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_262),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_199),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_267),
.Y(n_318)
);

NAND2xp33_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_278),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_248),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_271),
.B(n_203),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_293),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_273),
.B(n_275),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_209),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_280),
.B(n_290),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_209),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_252),
.B(n_147),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_210),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_283),
.B(n_210),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_265),
.B(n_217),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_253),
.B(n_211),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_254),
.B(n_211),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_SL g338 ( 
.A(n_256),
.B(n_150),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_259),
.B(n_217),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_L g340 ( 
.A(n_249),
.B(n_213),
.C(n_226),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_289),
.B(n_151),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_269),
.B(n_217),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_250),
.B(n_217),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_251),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_283),
.Y(n_345)
);

A2O1A1Ixp33_ASAP7_75t_L g346 ( 
.A1(n_251),
.A2(n_243),
.B(n_179),
.C(n_202),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_268),
.B(n_219),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_284),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_291),
.B(n_219),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_284),
.Y(n_350)
);

NOR3xp33_ASAP7_75t_L g351 ( 
.A(n_251),
.B(n_173),
.C(n_200),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_261),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_L g353 ( 
.A(n_251),
.B(n_171),
.C(n_198),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_291),
.B(n_219),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_297),
.B(n_152),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_306),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_294),
.B(n_156),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_336),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_295),
.A2(n_174),
.B1(n_192),
.B2(n_191),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_296),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_167),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_302),
.A2(n_162),
.B1(n_188),
.B2(n_187),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_315),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_300),
.A2(n_219),
.B1(n_155),
.B2(n_184),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_313),
.A2(n_186),
.B(n_160),
.C(n_159),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_316),
.B(n_157),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_301),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

BUFx12f_ASAP7_75t_SL g370 ( 
.A(n_347),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_305),
.B(n_155),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_309),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_299),
.B(n_155),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_334),
.Y(n_375)
);

NOR3xp33_ASAP7_75t_SL g376 ( 
.A(n_353),
.B(n_45),
.C(n_46),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_310),
.B(n_135),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_335),
.B(n_49),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_351),
.B(n_51),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_323),
.B(n_53),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_314),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_307),
.A2(n_54),
.B(n_56),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_304),
.B(n_57),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_346),
.B(n_60),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_343),
.B(n_62),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_322),
.B(n_63),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_303),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_317),
.A2(n_66),
.B(n_67),
.C(n_72),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_338),
.B(n_74),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_298),
.B(n_133),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_326),
.B(n_75),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_331),
.B(n_76),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_312),
.B(n_83),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_328),
.A2(n_84),
.B1(n_85),
.B2(n_89),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_340),
.B(n_90),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_308),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_307),
.A2(n_92),
.B(n_93),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_308),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_311),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

AND2x4_ASAP7_75t_SL g411 ( 
.A(n_325),
.B(n_95),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_329),
.B(n_96),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_349),
.B(n_132),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_317),
.B(n_97),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_410),
.Y(n_416)
);

O2A1O1Ixp33_ASAP7_75t_SL g417 ( 
.A1(n_382),
.A2(n_330),
.B(n_333),
.C(n_332),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_364),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_359),
.A2(n_328),
.B1(n_332),
.B2(n_333),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_361),
.B(n_354),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_329),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_413),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_375),
.B(n_327),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_359),
.A2(n_330),
.B1(n_341),
.B2(n_345),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_363),
.A2(n_345),
.B1(n_100),
.B2(n_101),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_365),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_369),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_358),
.B(n_108),
.Y(n_428)
);

A2O1A1Ixp33_ASAP7_75t_L g429 ( 
.A1(n_382),
.A2(n_407),
.B(n_378),
.C(n_380),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_371),
.A2(n_111),
.B(n_113),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_356),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_377),
.A2(n_120),
.B(n_122),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_374),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_358),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_L g436 ( 
.A1(n_412),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_355),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_401),
.A2(n_414),
.B(n_398),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_384),
.B(n_394),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_357),
.B(n_381),
.Y(n_441)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_357),
.B(n_381),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_399),
.A2(n_368),
.B1(n_372),
.B2(n_388),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_374),
.A2(n_399),
.B1(n_362),
.B2(n_387),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_385),
.A2(n_389),
.B(n_402),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_374),
.Y(n_448)
);

NOR3xp33_ASAP7_75t_L g449 ( 
.A(n_367),
.B(n_379),
.C(n_366),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_397),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_402),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_386),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_L g455 ( 
.A1(n_376),
.A2(n_391),
.B(n_383),
.C(n_403),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_415),
.B(n_395),
.Y(n_456)
);

AO21x2_ASAP7_75t_L g457 ( 
.A1(n_429),
.A2(n_400),
.B(n_392),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_404),
.Y(n_458)
);

AOI22x1_ASAP7_75t_L g459 ( 
.A1(n_446),
.A2(n_409),
.B1(n_408),
.B2(n_386),
.Y(n_459)
);

INVx3_ASAP7_75t_SL g460 ( 
.A(n_442),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_419),
.A2(n_406),
.B(n_386),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_450),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_408),
.Y(n_463)
);

AO21x2_ASAP7_75t_L g464 ( 
.A1(n_417),
.A2(n_408),
.B(n_406),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_418),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_435),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_439),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_422),
.Y(n_471)
);

INVx6_ASAP7_75t_SL g472 ( 
.A(n_454),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_437),
.B(n_406),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_419),
.A2(n_430),
.B(n_433),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_427),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

OR3x4_ASAP7_75t_SL g479 ( 
.A(n_447),
.B(n_425),
.C(n_443),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_423),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_441),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_448),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_421),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_454),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_462),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_460),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_460),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_472),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

INVx8_ASAP7_75t_L g491 ( 
.A(n_484),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_469),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_461),
.A2(n_455),
.B(n_445),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_462),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_458),
.A2(n_420),
.B1(n_434),
.B2(n_449),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_472),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_465),
.Y(n_497)
);

AO21x2_ASAP7_75t_L g498 ( 
.A1(n_475),
.A2(n_424),
.B(n_428),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_471),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_465),
.Y(n_500)
);

BUFx2_ASAP7_75t_R g501 ( 
.A(n_477),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_458),
.A2(n_476),
.B1(n_434),
.B2(n_473),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_470),
.A2(n_426),
.B1(n_424),
.B2(n_431),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_477),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_475),
.A2(n_426),
.B(n_436),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_471),
.Y(n_508)
);

BUFx2_ASAP7_75t_R g509 ( 
.A(n_467),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_485),
.B(n_463),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_487),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_499),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_506),
.A2(n_457),
.B(n_456),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_463),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_497),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_464),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_486),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_492),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_495),
.A2(n_479),
.B(n_481),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_504),
.B(n_480),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_505),
.Y(n_523)
);

AND2x4_ASAP7_75t_SL g524 ( 
.A(n_487),
.B(n_468),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_487),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_498),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_507),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_505),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_493),
.B(n_502),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_488),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_R g531 ( 
.A(n_489),
.B(n_474),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_500),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_478),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_495),
.B(n_478),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_509),
.B(n_468),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_509),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_501),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_503),
.A2(n_470),
.B1(n_482),
.B2(n_457),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_R g539 ( 
.A(n_489),
.B(n_490),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_491),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_529),
.B(n_498),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_510),
.B(n_507),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_532),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_513),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_518),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_511),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_506),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_519),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_517),
.B(n_464),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_515),
.B(n_464),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_538),
.A2(n_482),
.B1(n_491),
.B2(n_484),
.Y(n_551)
);

AO21x2_ASAP7_75t_L g552 ( 
.A1(n_514),
.A2(n_456),
.B(n_459),
.Y(n_552)
);

AOI221xp5_ASAP7_75t_L g553 ( 
.A1(n_521),
.A2(n_490),
.B1(n_491),
.B2(n_496),
.C(n_522),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_496),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_510),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_533),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_534),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_534),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_528),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_547),
.B(n_512),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_559),
.B(n_536),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_544),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_547),
.B(n_526),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_546),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_532),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_545),
.B(n_520),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_556),
.B(n_523),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_558),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_542),
.B(n_543),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_543),
.B(n_535),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_548),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_555),
.B(n_525),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_554),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_557),
.B(n_527),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_569),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_566),
.B(n_549),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_569),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_563),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_564),
.B(n_541),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_574),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_570),
.B(n_541),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_564),
.A2(n_551),
.B(n_553),
.Y(n_583)
);

AOI322xp5_ASAP7_75t_L g584 ( 
.A1(n_582),
.A2(n_551),
.A3(n_537),
.B1(n_561),
.B2(n_555),
.C1(n_572),
.C2(n_571),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_576),
.B(n_562),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_580),
.B(n_567),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_578),
.B(n_568),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_579),
.Y(n_588)
);

NOR2x1p5_ASAP7_75t_SL g589 ( 
.A(n_581),
.B(n_565),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_581),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_588),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_585),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_586),
.B(n_575),
.Y(n_593)
);

AOI211xp5_ASAP7_75t_L g594 ( 
.A1(n_587),
.A2(n_583),
.B(n_573),
.C(n_575),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_590),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_591),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_594),
.A2(n_592),
.B(n_595),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_593),
.Y(n_598)
);

AOI21xp33_ASAP7_75t_L g599 ( 
.A1(n_594),
.A2(n_539),
.B(n_583),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_L g600 ( 
.A1(n_592),
.A2(n_531),
.B1(n_584),
.B2(n_537),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_596),
.B(n_516),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_600),
.A2(n_566),
.B1(n_525),
.B2(n_530),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_598),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_603),
.Y(n_604)
);

A2O1A1Ixp33_ASAP7_75t_SL g605 ( 
.A1(n_601),
.A2(n_597),
.B(n_599),
.C(n_530),
.Y(n_605)
);

AOI221xp5_ASAP7_75t_L g606 ( 
.A1(n_604),
.A2(n_602),
.B1(n_584),
.B2(n_516),
.C(n_550),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_606),
.Y(n_607)
);

NOR2x1p5_ASAP7_75t_L g608 ( 
.A(n_607),
.B(n_605),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_608),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_609),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_610),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_524),
.Y(n_612)
);

OAI22xp33_ASAP7_75t_L g613 ( 
.A1(n_612),
.A2(n_560),
.B1(n_540),
.B2(n_589),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_613),
.B(n_524),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_614),
.A2(n_540),
.B1(n_560),
.B2(n_577),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_615),
.B(n_540),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_616),
.A2(n_552),
.B1(n_560),
.B2(n_577),
.Y(n_617)
);


endmodule