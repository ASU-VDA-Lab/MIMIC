module fake_netlist_5_2537_n_1858 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1858);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1858;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_14),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_28),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_3),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_105),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_135),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_88),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_96),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_51),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_73),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_17),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_45),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_118),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_104),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_155),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_61),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_147),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_67),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_27),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_20),
.Y(n_216)
);

CKINVDCx11_ASAP7_75t_R g217 ( 
.A(n_81),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_129),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_86),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_66),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_8),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_156),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_101),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_98),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_112),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_95),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_57),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_65),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_61),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_119),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_149),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_128),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_41),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_27),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_79),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_97),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_70),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_110),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_66),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_43),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_74),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_13),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_141),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_60),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_109),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_25),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_76),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_148),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_7),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_49),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_10),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_94),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_50),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_180),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_92),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_16),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_122),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_158),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_166),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_64),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_138),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_100),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_0),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_62),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_35),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_126),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_165),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_33),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_31),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_4),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_91),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_115),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_21),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_49),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_42),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_24),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_93),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_181),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_174),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_78),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_71),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_134),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_19),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_130),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_28),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_9),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_143),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_32),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_176),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_45),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_56),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_120),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_15),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_21),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_72),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_32),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_107),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_41),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_58),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_15),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_154),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_132),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_69),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_2),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_24),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_4),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_177),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_85),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_14),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_64),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_182),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_26),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_39),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_157),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_5),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_43),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_53),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_29),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_31),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_39),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_42),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_6),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_77),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_58),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_29),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_103),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_17),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_178),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_22),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_84),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_0),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_51),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_127),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_152),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_8),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_7),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_136),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_131),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_37),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_40),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_1),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_153),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_167),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_16),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_160),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_90),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_102),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_133),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_151),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_123),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_59),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_10),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_80),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_55),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_56),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_6),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_252),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_R g366 ( 
.A(n_204),
.B(n_183),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_252),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_197),
.B(n_1),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_305),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_268),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_217),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_214),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_268),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_218),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_277),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_254),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_321),
.B(n_2),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_277),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_185),
.B(n_3),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_245),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_260),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_329),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_189),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_184),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_184),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_193),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_214),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_187),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_187),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_191),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_191),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_205),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_208),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_288),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_199),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_202),
.B(n_5),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_212),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_231),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_239),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_240),
.Y(n_401)
);

INVxp33_ASAP7_75t_SL g402 ( 
.A(n_186),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_199),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_216),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_254),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_216),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_185),
.B(n_9),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_222),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_315),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_222),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_319),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_188),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_227),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_227),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_235),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_196),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_243),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_244),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_235),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_249),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_251),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_237),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g423 ( 
.A(n_237),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_253),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_256),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_261),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_262),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_261),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_273),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_346),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_273),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_276),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_276),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_278),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_353),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_225),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_263),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_196),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_188),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_265),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_266),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_267),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_278),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_274),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_275),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_203),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_291),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_309),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_225),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_291),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_279),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_215),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_280),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_285),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_299),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_223),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_384),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_387),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_286),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_367),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_367),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_412),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_416),
.B(n_204),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_439),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_393),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_394),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_385),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_386),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_398),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_436),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_376),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_438),
.B(n_287),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_448),
.B(n_204),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_390),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_SL g483 ( 
.A(n_366),
.B(n_259),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_438),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_372),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_365),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_374),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_391),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_380),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_399),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_391),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_R g492 ( 
.A(n_371),
.B(n_289),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_392),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_396),
.B(n_309),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_206),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_400),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_370),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_370),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_401),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_403),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_404),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_406),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_417),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_373),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_372),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_379),
.B(n_407),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_388),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_406),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_408),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_408),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_410),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_418),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_388),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_410),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_373),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_446),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_413),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_413),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_375),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_446),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_420),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_421),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_375),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_382),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_414),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_395),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_378),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_424),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_415),
.A2(n_233),
.B(n_206),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_485),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_465),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_459),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_459),
.Y(n_539)
);

BUFx4f_ASAP7_75t_L g540 ( 
.A(n_466),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_510),
.B(n_449),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_465),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_464),
.B(n_233),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_459),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_457),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_509),
.B(n_259),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_510),
.B(n_516),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_509),
.B(n_402),
.Y(n_548)
);

AND2x6_ASAP7_75t_L g549 ( 
.A(n_464),
.B(n_190),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_485),
.B(n_456),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g551 ( 
.A(n_523),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_470),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_508),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_484),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_484),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_463),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_470),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_472),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_463),
.Y(n_560)
);

AND2x6_ASAP7_75t_L g561 ( 
.A(n_464),
.B(n_190),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_479),
.A2(n_377),
.B1(n_369),
.B2(n_368),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_479),
.B(n_194),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_516),
.B(n_449),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_479),
.B(n_378),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_495),
.B(n_381),
.Y(n_566)
);

BUFx4f_ASAP7_75t_L g567 ( 
.A(n_466),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_484),
.B(n_230),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_466),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_472),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_468),
.B(n_425),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_475),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_469),
.B(n_427),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_463),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_483),
.A2(n_453),
.B1(n_454),
.B2(n_440),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_527),
.Y(n_576)
);

BUFx4f_ASAP7_75t_L g577 ( 
.A(n_466),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_484),
.B(n_230),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_508),
.B(n_452),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_473),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_484),
.Y(n_581)
);

NOR3xp33_ASAP7_75t_L g582 ( 
.A(n_519),
.B(n_405),
.C(n_347),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_527),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_475),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_527),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_460),
.B(n_230),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_490),
.B(n_437),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_466),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_478),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_L g590 ( 
.A1(n_519),
.A2(n_405),
.B1(n_423),
.B2(n_234),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_476),
.A2(n_508),
.B1(n_500),
.B2(n_506),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_460),
.B(n_441),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_477),
.B(n_442),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_478),
.Y(n_594)
);

BUFx4f_ASAP7_75t_L g595 ( 
.A(n_466),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_477),
.B(n_230),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_495),
.B(n_444),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_458),
.B(n_230),
.Y(n_598)
);

INVx6_ASAP7_75t_L g599 ( 
.A(n_495),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_527),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_497),
.B(n_445),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_495),
.B(n_451),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_467),
.B(n_246),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_496),
.B(n_194),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_527),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_466),
.B(n_195),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_527),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_L g608 ( 
.A1(n_476),
.A2(n_284),
.B1(n_224),
.B2(n_364),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_SL g609 ( 
.A(n_474),
.B(n_397),
.Y(n_609)
);

AND2x2_ASAP7_75t_SL g610 ( 
.A(n_496),
.B(n_195),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_458),
.B(n_198),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_523),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_467),
.B(n_341),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_480),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_458),
.B(n_452),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_474),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_515),
.A2(n_435),
.B1(n_430),
.B2(n_411),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_524),
.A2(n_282),
.B1(n_363),
.B2(n_362),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_527),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_480),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_467),
.B(n_358),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_467),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_496),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_458),
.B(n_198),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_458),
.B(n_200),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_492),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_496),
.B(n_200),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_471),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_496),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_471),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_461),
.B(n_290),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_471),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_461),
.B(n_295),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_526),
.B(n_409),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_471),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_461),
.B(n_297),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_487),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_461),
.B(n_300),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_486),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_533),
.B(n_201),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_532),
.B(n_455),
.C(n_242),
.Y(n_641)
);

OAI21xp33_ASAP7_75t_L g642 ( 
.A1(n_481),
.A2(n_488),
.B(n_482),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_481),
.B(n_381),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_533),
.B(n_301),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_489),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_482),
.B(n_301),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_533),
.B(n_201),
.Y(n_647)
);

AND2x2_ASAP7_75t_SL g648 ( 
.A(n_488),
.B(n_207),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_492),
.B(n_207),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_491),
.B(n_210),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_491),
.B(n_210),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_486),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_493),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_493),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_494),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_494),
.B(n_303),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_501),
.B(n_211),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_501),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_486),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_486),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_502),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_502),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_503),
.B(n_211),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_528),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_503),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_504),
.A2(n_352),
.B1(n_313),
.B2(n_328),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_504),
.B(n_213),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_505),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_530),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_505),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_499),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_511),
.B(n_213),
.Y(n_672)
);

BUFx4f_ASAP7_75t_L g673 ( 
.A(n_511),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_499),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_512),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_512),
.B(n_310),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_513),
.B(n_219),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_513),
.B(n_419),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_499),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_499),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_514),
.A2(n_317),
.B1(n_271),
.B2(n_360),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_514),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_517),
.B(n_219),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_498),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_535),
.B(n_422),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_517),
.A2(n_352),
.B1(n_299),
.B2(n_313),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_498),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_520),
.B(n_422),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_538),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_538),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_548),
.B(n_241),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_565),
.A2(n_324),
.B(n_320),
.C(n_323),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_552),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_648),
.B(n_220),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_629),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_592),
.B(n_247),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_549),
.A2(n_331),
.B1(n_361),
.B2(n_311),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_566),
.Y(n_698)
);

OAI22x1_ASAP7_75t_L g699 ( 
.A1(n_612),
.A2(n_397),
.B1(n_326),
.B2(n_325),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_610),
.B(n_316),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_539),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_566),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_610),
.B(n_322),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_648),
.B(n_334),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_550),
.B(n_520),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_673),
.B(n_338),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_552),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_549),
.A2(n_350),
.B1(n_354),
.B2(n_356),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_593),
.B(n_220),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_673),
.B(n_221),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_673),
.B(n_221),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_555),
.B(n_556),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_549),
.A2(n_342),
.B1(n_229),
.B2(n_232),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_555),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_536),
.B(n_521),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_555),
.B(n_226),
.Y(n_716)
);

AND3x1_ASAP7_75t_L g717 ( 
.A(n_582),
.B(n_320),
.C(n_323),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_SL g718 ( 
.A(n_626),
.B(n_545),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_643),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_612),
.B(n_521),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_539),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_549),
.A2(n_336),
.B1(n_226),
.B2(n_229),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_599),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_565),
.B(n_232),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_556),
.B(n_238),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_623),
.B(n_238),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_615),
.A2(n_343),
.B1(n_257),
.B2(n_314),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_544),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_643),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_556),
.B(n_255),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_678),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_623),
.B(n_255),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_549),
.B(n_561),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_581),
.B(n_269),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_549),
.B(n_269),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_561),
.B(n_563),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_579),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_561),
.B(n_270),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_561),
.B(n_270),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_562),
.A2(n_357),
.B1(n_342),
.B2(n_336),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_547),
.B(n_525),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_544),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_557),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_561),
.B(n_292),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_561),
.B(n_292),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_563),
.B(n_345),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_546),
.B(n_525),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_563),
.B(n_345),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_563),
.B(n_351),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_557),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_599),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_581),
.B(n_351),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_571),
.B(n_248),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_546),
.A2(n_357),
.B1(n_355),
.B2(n_272),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_685),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_563),
.B(n_639),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_563),
.B(n_355),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_573),
.B(n_250),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_599),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_581),
.B(n_192),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_639),
.B(n_529),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_639),
.B(n_529),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_597),
.A2(n_518),
.B(n_531),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_680),
.B(n_534),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_560),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_688),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_543),
.A2(n_535),
.B1(n_534),
.B2(n_264),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_560),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_630),
.B(n_192),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_680),
.B(n_498),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_551),
.B(n_209),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_602),
.A2(n_567),
.B(n_540),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_630),
.B(n_192),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_630),
.B(n_192),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_574),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_537),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_587),
.B(n_258),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_543),
.A2(n_324),
.B1(n_337),
.B2(n_328),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_680),
.B(n_507),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_574),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_542),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_628),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_652),
.B(n_228),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_553),
.B(n_558),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_652),
.B(n_671),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_559),
.B(n_507),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_570),
.B(n_507),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_657),
.A2(n_337),
.B(n_327),
.C(n_339),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_652),
.B(n_228),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_671),
.B(n_228),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_572),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_671),
.B(n_228),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_551),
.B(n_209),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_541),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_628),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_554),
.B(n_531),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_584),
.B(n_518),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_601),
.B(n_281),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_554),
.B(n_283),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_589),
.B(n_518),
.Y(n_800)
);

INVx8_ASAP7_75t_L g801 ( 
.A(n_543),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_SL g802 ( 
.A1(n_564),
.A2(n_308),
.B1(n_209),
.B2(n_236),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_594),
.B(n_522),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_L g804 ( 
.A(n_543),
.B(n_293),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_543),
.A2(n_327),
.B1(n_339),
.B2(n_531),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_650),
.Y(n_806)
);

AOI221xp5_ASAP7_75t_L g807 ( 
.A1(n_590),
.A2(n_344),
.B1(n_296),
.B2(n_298),
.C(n_302),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_618),
.B(n_611),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_611),
.B(n_294),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_543),
.A2(n_625),
.B1(n_624),
.B2(n_598),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_632),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_624),
.B(n_304),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_625),
.A2(n_462),
.B1(n_522),
.B2(n_359),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_622),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_614),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_626),
.B(n_641),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_620),
.B(n_522),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_640),
.B(n_462),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_540),
.A2(n_383),
.B(n_447),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_653),
.B(n_426),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_598),
.A2(n_348),
.B1(n_306),
.B2(n_307),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_654),
.B(n_426),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_655),
.B(n_658),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_540),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_632),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_546),
.B(n_209),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_546),
.B(n_236),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_575),
.B(n_312),
.Y(n_828)
);

NOR2xp67_ASAP7_75t_L g829 ( 
.A(n_617),
.B(n_616),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_L g830 ( 
.A1(n_661),
.A2(n_665),
.B1(n_668),
.B2(n_670),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_662),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_640),
.B(n_318),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_591),
.B(n_75),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_640),
.B(n_330),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_675),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_647),
.B(n_635),
.Y(n_836)
);

OAI22x1_ASAP7_75t_SL g837 ( 
.A1(n_637),
.A2(n_332),
.B1(n_333),
.B2(n_335),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_682),
.A2(n_340),
.B1(n_349),
.B2(n_443),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_649),
.B(n_656),
.Y(n_839)
);

NAND2x1p5_ASAP7_75t_L g840 ( 
.A(n_647),
.B(n_450),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_676),
.B(n_450),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_603),
.B(n_447),
.Y(n_842)
);

INVxp33_ASAP7_75t_L g843 ( 
.A(n_634),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_647),
.B(n_236),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_635),
.B(n_236),
.Y(n_845)
);

OAI22x1_ASAP7_75t_SL g846 ( 
.A1(n_645),
.A2(n_443),
.B1(n_434),
.B2(n_433),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_613),
.B(n_434),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_642),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_644),
.A2(n_433),
.B1(n_432),
.B2(n_431),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_545),
.B(n_432),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_644),
.A2(n_431),
.B1(n_429),
.B2(n_428),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_649),
.B(n_608),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_621),
.B(n_429),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_622),
.B(n_428),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_664),
.B(n_383),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_604),
.A2(n_173),
.B1(n_169),
.B2(n_168),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_646),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_622),
.B(n_164),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_659),
.B(n_660),
.Y(n_859)
);

NOR2xp67_ASAP7_75t_L g860 ( 
.A(n_631),
.B(n_162),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_785),
.A2(n_567),
.B(n_595),
.Y(n_861)
);

AO21x1_ASAP7_75t_L g862 ( 
.A1(n_808),
.A2(n_596),
.B(n_586),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_836),
.A2(n_586),
.B(n_596),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_785),
.A2(n_567),
.B(n_577),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_691),
.B(n_669),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_852),
.A2(n_667),
.B(n_650),
.C(n_660),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_712),
.A2(n_577),
.B(n_595),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_840),
.Y(n_868)
);

AOI22x1_ASAP7_75t_L g869 ( 
.A1(n_814),
.A2(n_674),
.B1(n_679),
.B2(n_650),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_L g870 ( 
.A(n_801),
.B(n_604),
.Y(n_870)
);

NOR2x1_ASAP7_75t_L g871 ( 
.A(n_816),
.B(n_681),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_794),
.B(n_857),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_740),
.A2(n_657),
.B(n_677),
.C(n_672),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_712),
.A2(n_595),
.B(n_577),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_843),
.B(n_580),
.Y(n_875)
);

AO21x1_ASAP7_75t_L g876 ( 
.A1(n_694),
.A2(n_568),
.B(n_578),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_696),
.B(n_580),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_836),
.A2(n_644),
.B(n_568),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_756),
.A2(n_644),
.B(n_578),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_824),
.A2(n_636),
.B(n_633),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_839),
.B(n_667),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_824),
.A2(n_638),
.B(n_576),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_843),
.B(n_580),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_753),
.B(n_667),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_710),
.A2(n_672),
.B(n_683),
.C(n_677),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_824),
.A2(n_619),
.B(n_576),
.Y(n_886)
);

BUFx4f_ASAP7_75t_L g887 ( 
.A(n_855),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_818),
.A2(n_619),
.B(n_583),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_698),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_709),
.B(n_651),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_818),
.A2(n_607),
.B(n_583),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_741),
.B(n_674),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_SL g893 ( 
.A1(n_716),
.A2(n_683),
.B(n_679),
.C(n_607),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_810),
.A2(n_686),
.B1(n_666),
.B2(n_588),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_704),
.A2(n_606),
.B(n_684),
.C(n_687),
.Y(n_895)
);

INVx11_ASAP7_75t_L g896 ( 
.A(n_718),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_714),
.A2(n_585),
.B(n_600),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_714),
.A2(n_585),
.B(n_600),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_737),
.B(n_609),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_714),
.A2(n_605),
.B(n_569),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_763),
.A2(n_605),
.B(n_588),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_841),
.B(n_663),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_772),
.A2(n_569),
.B(n_588),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_758),
.B(n_663),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_767),
.A2(n_569),
.B1(n_684),
.B2(n_687),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_715),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_733),
.A2(n_736),
.B1(n_806),
.B2(n_848),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_801),
.A2(n_859),
.B(n_762),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_777),
.B(n_663),
.Y(n_909)
);

BUFx12f_ASAP7_75t_L g910 ( 
.A(n_705),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_693),
.B(n_687),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_R g912 ( 
.A(n_804),
.B(n_604),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_L g913 ( 
.A(n_828),
.B(n_606),
.C(n_684),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_795),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_702),
.A2(n_725),
.B(n_716),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_798),
.B(n_663),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_801),
.A2(n_627),
.B(n_604),
.Y(n_917)
);

CKINVDCx8_ASAP7_75t_R g918 ( 
.A(n_809),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_725),
.A2(n_627),
.B(n_604),
.Y(n_919)
);

AO22x1_ASAP7_75t_L g920 ( 
.A1(n_812),
.A2(n_663),
.B1(n_651),
.B2(n_627),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_811),
.Y(n_921)
);

AOI21x1_ASAP7_75t_L g922 ( 
.A1(n_796),
.A2(n_627),
.B(n_604),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_842),
.B(n_651),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_799),
.A2(n_663),
.B(n_651),
.C(n_627),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_719),
.A2(n_651),
.B1(n_627),
.B2(n_18),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_761),
.A2(n_651),
.B(n_161),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_720),
.B(n_695),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_704),
.A2(n_11),
.B(n_12),
.C(n_19),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_825),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_730),
.A2(n_140),
.B(n_139),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_707),
.A2(n_125),
.B1(n_124),
.B2(n_121),
.Y(n_931)
);

NAND2x1_ASAP7_75t_L g932 ( 
.A(n_723),
.B(n_113),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_764),
.A2(n_108),
.B(n_106),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_844),
.B(n_11),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_844),
.B(n_12),
.Y(n_935)
);

O2A1O1Ixp5_ASAP7_75t_L g936 ( 
.A1(n_710),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_693),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_693),
.A2(n_99),
.B1(n_83),
.B2(n_82),
.Y(n_938)
);

O2A1O1Ixp5_ASAP7_75t_SL g939 ( 
.A1(n_711),
.A2(n_23),
.B(n_25),
.C(n_26),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_730),
.A2(n_752),
.B(n_734),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_825),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_734),
.A2(n_30),
.B(n_33),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_752),
.A2(n_30),
.B(n_34),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_L g944 ( 
.A(n_754),
.B(n_34),
.C(n_35),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_770),
.A2(n_36),
.B(n_37),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_779),
.A2(n_796),
.B(n_823),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_784),
.A2(n_38),
.B(n_40),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_846),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_769),
.A2(n_38),
.B(n_44),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_769),
.A2(n_44),
.B(n_46),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_773),
.A2(n_46),
.B(n_47),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_692),
.A2(n_832),
.B(n_834),
.C(n_703),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_771),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_751),
.A2(n_68),
.B1(n_48),
.B2(n_52),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_689),
.Y(n_955)
);

OAI321xp33_ASAP7_75t_L g956 ( 
.A1(n_807),
.A2(n_47),
.A3(n_48),
.B1(n_52),
.B2(n_54),
.C(n_55),
.Y(n_956)
);

NAND3xp33_ASAP7_75t_SL g957 ( 
.A(n_802),
.B(n_54),
.C(n_57),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_689),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_773),
.A2(n_59),
.B(n_60),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_774),
.A2(n_62),
.B(n_63),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_793),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_729),
.B(n_63),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_774),
.A2(n_65),
.B(n_67),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_723),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_751),
.A2(n_68),
.B1(n_759),
.B2(n_722),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_L g966 ( 
.A(n_727),
.B(n_829),
.C(n_834),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_832),
.A2(n_833),
.B(n_747),
.C(n_724),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_847),
.B(n_853),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_735),
.A2(n_745),
.B(n_757),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_783),
.A2(n_792),
.B(n_789),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_783),
.A2(n_792),
.B(n_789),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_776),
.B(n_781),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_791),
.B(n_815),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_831),
.B(n_835),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_778),
.A2(n_711),
.B1(n_703),
.B2(n_700),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_731),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_830),
.B(n_759),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_854),
.B(n_766),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_755),
.B(n_723),
.Y(n_979)
);

NOR2xp67_ASAP7_75t_SL g980 ( 
.A(n_723),
.B(n_790),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_738),
.A2(n_749),
.B(n_746),
.C(n_748),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_726),
.B(n_732),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_790),
.A2(n_760),
.B(n_706),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_760),
.B(n_700),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_739),
.A2(n_744),
.B(n_690),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_820),
.B(n_822),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_706),
.A2(n_797),
.B(n_803),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_805),
.A2(n_708),
.B1(n_697),
.B2(n_713),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_826),
.B(n_827),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_786),
.B(n_787),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_800),
.A2(n_817),
.B(n_858),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_690),
.B(n_780),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_701),
.A2(n_780),
.B(n_775),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_701),
.A2(n_743),
.B(n_768),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_845),
.B(n_821),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_849),
.A2(n_851),
.B1(n_717),
.B2(n_845),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_837),
.B(n_838),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_721),
.B(n_768),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_692),
.A2(n_788),
.B(n_819),
.C(n_742),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_813),
.A2(n_860),
.B(n_728),
.C(n_742),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_728),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_743),
.B(n_750),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_699),
.B(n_750),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_765),
.A2(n_775),
.B(n_856),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_765),
.B(n_548),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_740),
.A2(n_509),
.B(n_694),
.C(n_852),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_801),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_691),
.B(n_548),
.Y(n_1008)
);

OA22x2_ASAP7_75t_L g1009 ( 
.A1(n_740),
.A2(n_546),
.B1(n_794),
.B2(n_699),
.Y(n_1009)
);

AOI22x1_ASAP7_75t_L g1010 ( 
.A1(n_814),
.A2(n_848),
.B1(n_782),
.B2(n_811),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_850),
.B(n_548),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_808),
.A2(n_839),
.B1(n_691),
.B2(n_852),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_850),
.B(n_548),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_850),
.B(n_548),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_691),
.B(n_548),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1017)
);

NOR2xp67_ASAP7_75t_SL g1018 ( 
.A(n_824),
.B(n_714),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_L g1019 ( 
.A(n_801),
.B(n_543),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_808),
.A2(n_839),
.B1(n_691),
.B2(n_852),
.Y(n_1020)
);

NOR2x1_ASAP7_75t_L g1021 ( 
.A(n_816),
.B(n_591),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_715),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_691),
.A2(n_548),
.B(n_852),
.C(n_808),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_691),
.B(n_548),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_SL g1030 ( 
.A(n_731),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_836),
.A2(n_818),
.B(n_796),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_808),
.A2(n_839),
.B1(n_691),
.B2(n_852),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_691),
.B(n_548),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1035)
);

AO32x1_ASAP7_75t_L g1036 ( 
.A1(n_740),
.A2(n_851),
.A3(n_849),
.B1(n_791),
.B2(n_815),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_SL g1037 ( 
.A(n_718),
.B(n_545),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_840),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_785),
.A2(n_712),
.B(n_556),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_691),
.B(n_548),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1016),
.B(n_1013),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_921),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1012),
.A2(n_1022),
.B(n_1017),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_906),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1026),
.A2(n_1028),
.B(n_1027),
.Y(n_1046)
);

NOR2x1_ASAP7_75t_L g1047 ( 
.A(n_877),
.B(n_1011),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1029),
.A2(n_1035),
.B(n_1033),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_1020),
.A2(n_1032),
.B(n_1024),
.C(n_1016),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_964),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1039),
.A2(n_1040),
.B(n_1019),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_872),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1008),
.B(n_1025),
.Y(n_1054)
);

AOI221xp5_ASAP7_75t_SL g1055 ( 
.A1(n_1006),
.A2(n_1041),
.B1(n_1034),
.B2(n_953),
.C(n_935),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_884),
.B(n_881),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_879),
.A2(n_878),
.B(n_864),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_869),
.A2(n_861),
.B(n_1004),
.Y(n_1059)
);

INVx6_ASAP7_75t_L g1060 ( 
.A(n_910),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1005),
.B(n_968),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_1031),
.A2(n_882),
.B(n_874),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_969),
.A2(n_867),
.B(n_908),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1005),
.B(n_986),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_948),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_SL g1066 ( 
.A1(n_930),
.A2(n_952),
.B(n_950),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_978),
.B(n_872),
.Y(n_1067)
);

AOI211x1_ASAP7_75t_L g1068 ( 
.A1(n_957),
.A2(n_1003),
.B(n_972),
.C(n_973),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_941),
.Y(n_1069)
);

AOI21x1_ASAP7_75t_L g1070 ( 
.A1(n_984),
.A2(n_980),
.B(n_987),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_927),
.B(n_953),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_904),
.A2(n_916),
.B(n_909),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_885),
.A2(n_940),
.B(n_866),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_927),
.B(n_990),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_934),
.A2(n_935),
.B(n_995),
.C(n_956),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_961),
.B(n_962),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_991),
.A2(n_922),
.B(n_891),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_966),
.A2(n_1021),
.B1(n_871),
.B2(n_865),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_888),
.A2(n_907),
.B(n_880),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_889),
.B(n_974),
.Y(n_1080)
);

AOI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_906),
.A2(n_1023),
.B(n_887),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_946),
.A2(n_886),
.B(n_900),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_982),
.B(n_1023),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_899),
.B(n_976),
.Y(n_1084)
);

OAI22x1_ASAP7_75t_L g1085 ( 
.A1(n_997),
.A2(n_934),
.B1(n_875),
.B2(n_883),
.Y(n_1085)
);

AO21x1_ASAP7_75t_L g1086 ( 
.A1(n_928),
.A2(n_913),
.B(n_988),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_981),
.A2(n_870),
.B(n_985),
.Y(n_1087)
);

CKINVDCx8_ASAP7_75t_R g1088 ( 
.A(n_962),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_890),
.A2(n_863),
.B(n_902),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_955),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_885),
.A2(n_967),
.B(n_915),
.Y(n_1091)
);

NAND2x1p5_ASAP7_75t_L g1092 ( 
.A(n_937),
.B(n_1007),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_897),
.A2(n_898),
.B(n_994),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_993),
.A2(n_895),
.B(n_905),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_999),
.A2(n_917),
.B(n_926),
.Y(n_1095)
);

NOR2x1_ASAP7_75t_SL g1096 ( 
.A(n_1007),
.B(n_937),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_887),
.B(n_875),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_SL g1098 ( 
.A1(n_1037),
.A2(n_997),
.B1(n_1009),
.B2(n_996),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_977),
.B(n_979),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_919),
.A2(n_923),
.B(n_924),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_937),
.Y(n_1101)
);

CKINVDCx11_ASAP7_75t_R g1102 ( 
.A(n_918),
.Y(n_1102)
);

INVx5_ASAP7_75t_L g1103 ( 
.A(n_964),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1018),
.A2(n_911),
.B(n_1002),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_SL g1105 ( 
.A1(n_949),
.A2(n_963),
.B(n_960),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_966),
.B(n_989),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_992),
.A2(n_876),
.B(n_862),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_L g1108 ( 
.A1(n_1000),
.A2(n_920),
.B(n_959),
.C(n_951),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_892),
.B(n_1038),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_975),
.A2(n_873),
.B(n_894),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_958),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_964),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1007),
.A2(n_937),
.B(n_998),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_914),
.A2(n_929),
.B(n_932),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_964),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1001),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1007),
.A2(n_998),
.B(n_893),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_925),
.B(n_975),
.Y(n_1118)
);

AOI221xp5_ASAP7_75t_L g1119 ( 
.A1(n_957),
.A2(n_944),
.B1(n_954),
.B2(n_965),
.C(n_1030),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1001),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_868),
.A2(n_933),
.B(n_1009),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_925),
.A2(n_944),
.B(n_936),
.C(n_942),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1001),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_931),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_913),
.B(n_947),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_943),
.B(n_945),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_939),
.B(n_912),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_938),
.A2(n_1036),
.B(n_896),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1036),
.A2(n_1024),
.B(n_1020),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_1036),
.A2(n_1024),
.B(n_983),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_1030),
.A2(n_862),
.A3(n_876),
.B(n_1024),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_921),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1135)
);

BUFx4f_ASAP7_75t_SL g1136 ( 
.A(n_910),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1024),
.A2(n_1020),
.B(n_1013),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_SL g1139 ( 
.A1(n_930),
.A2(n_952),
.B(n_970),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_862),
.A2(n_876),
.A3(n_1024),
.B(n_866),
.Y(n_1141)
);

NOR2xp67_ASAP7_75t_L g1142 ( 
.A(n_953),
.B(n_961),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_SL g1144 ( 
.A1(n_977),
.A2(n_1025),
.B(n_1008),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1024),
.A2(n_1016),
.B(n_1025),
.C(n_1008),
.Y(n_1145)
);

AOI221x1_ASAP7_75t_L g1146 ( 
.A1(n_1024),
.A2(n_1016),
.B1(n_1008),
.B2(n_1025),
.C(n_1034),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1013),
.A2(n_1020),
.B1(n_1032),
.B2(n_1024),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_921),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_948),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_937),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1013),
.A2(n_1020),
.B1(n_1032),
.B2(n_1024),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1013),
.A2(n_1020),
.B(n_1032),
.C(n_1024),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1013),
.B(n_1020),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1016),
.B(n_1013),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1024),
.A2(n_1020),
.B(n_1013),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1016),
.B(n_1013),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1016),
.B(n_1013),
.Y(n_1165)
);

AOI21xp33_ASAP7_75t_L g1166 ( 
.A1(n_1016),
.A2(n_1025),
.B(n_1008),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_862),
.A2(n_876),
.A3(n_1024),
.B(n_866),
.Y(n_1167)
);

AOI21xp33_ASAP7_75t_L g1168 ( 
.A1(n_1016),
.A2(n_1025),
.B(n_1008),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1169)
);

AOI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_1016),
.A2(n_1025),
.B(n_1008),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_887),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1024),
.A2(n_1020),
.B(n_1013),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_872),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_970),
.A2(n_971),
.B(n_983),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1013),
.A2(n_1020),
.B1(n_1032),
.B2(n_1024),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_910),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1016),
.B(n_1013),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_937),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_903),
.A2(n_1010),
.B(n_901),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1013),
.A2(n_1020),
.B1(n_1032),
.B2(n_1024),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_887),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1012),
.A2(n_785),
.B(n_712),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_887),
.Y(n_1194)
);

OA22x2_ASAP7_75t_L g1195 ( 
.A1(n_1013),
.A2(n_1032),
.B1(n_1020),
.B2(n_1025),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_964),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1061),
.B(n_1064),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1042),
.B(n_1157),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1076),
.B(n_1171),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1076),
.B(n_1192),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1084),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1163),
.A2(n_1187),
.B1(n_1165),
.B2(n_1075),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1166),
.B(n_1168),
.Y(n_1203)
);

BUFx4_ASAP7_75t_SL g1204 ( 
.A(n_1065),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1058),
.A2(n_1063),
.B(n_1072),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1090),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1054),
.B(n_1146),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1074),
.B(n_1145),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_SL g1209 ( 
.A(n_1136),
.B(n_1088),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1060),
.Y(n_1210)
);

NAND2xp33_ASAP7_75t_L g1211 ( 
.A(n_1075),
.B(n_1050),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1067),
.B(n_1049),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1045),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1153),
.B(n_1180),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1156),
.B(n_1170),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1150),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1069),
.Y(n_1217)
);

INVx4_ASAP7_75t_L g1218 ( 
.A(n_1188),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_SL g1219 ( 
.A1(n_1110),
.A2(n_1137),
.B(n_1162),
.C(n_1172),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1133),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1076),
.B(n_1194),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1059),
.A2(n_1077),
.B(n_1052),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1142),
.B(n_1106),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1045),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1148),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1059),
.A2(n_1077),
.B(n_1062),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1087),
.A2(n_1044),
.B(n_1046),
.Y(n_1227)
);

INVx3_ASAP7_75t_SL g1228 ( 
.A(n_1060),
.Y(n_1228)
);

OR2x6_ASAP7_75t_L g1229 ( 
.A(n_1060),
.B(n_1150),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1186),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1118),
.A2(n_1050),
.B1(n_1152),
.B2(n_1195),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1097),
.B(n_1185),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1156),
.B(n_1152),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1078),
.A2(n_1147),
.B(n_1182),
.C(n_1151),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1048),
.A2(n_1181),
.B(n_1173),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1190),
.B(n_1083),
.Y(n_1236)
);

O2A1O1Ixp5_ASAP7_75t_L g1237 ( 
.A1(n_1086),
.A2(n_1129),
.B(n_1118),
.C(n_1191),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1135),
.A2(n_1161),
.B(n_1169),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1053),
.B(n_1175),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1150),
.B(n_1103),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1188),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1195),
.B(n_1098),
.Y(n_1242)
);

OR2x6_ASAP7_75t_SL g1243 ( 
.A(n_1071),
.B(n_1099),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1138),
.A2(n_1193),
.B(n_1155),
.Y(n_1244)
);

AOI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1055),
.A2(n_1085),
.B(n_1057),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1115),
.B(n_1047),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1188),
.B(n_1092),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1154),
.A2(n_1183),
.B(n_1177),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1136),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1081),
.B(n_1080),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1057),
.B(n_1068),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1123),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1125),
.B(n_1123),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1119),
.B(n_1109),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1111),
.B(n_1131),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1102),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1139),
.A2(n_1073),
.B(n_1091),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1102),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1103),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1125),
.B(n_1131),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1120),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1100),
.A2(n_1089),
.B(n_1107),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1065),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1122),
.A2(n_1124),
.B1(n_1127),
.B2(n_1125),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1149),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1115),
.B(n_1103),
.Y(n_1266)
);

NAND2xp33_ASAP7_75t_L g1267 ( 
.A(n_1092),
.B(n_1122),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1149),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1131),
.B(n_1051),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1131),
.B(n_1116),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1116),
.B(n_1167),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1066),
.A2(n_1117),
.B(n_1126),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1062),
.A2(n_1093),
.B(n_1082),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1112),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1101),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1107),
.A2(n_1108),
.B(n_1128),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1121),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1196),
.A2(n_1113),
.B1(n_1101),
.B2(n_1070),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1128),
.A2(n_1130),
.B1(n_1095),
.B2(n_1114),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1114),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1141),
.B(n_1167),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1105),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1141),
.B(n_1167),
.Y(n_1283)
);

OR2x6_ASAP7_75t_L g1284 ( 
.A(n_1095),
.B(n_1094),
.Y(n_1284)
);

CKINVDCx6p67_ASAP7_75t_R g1285 ( 
.A(n_1144),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1141),
.B(n_1167),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1141),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1056),
.A2(n_1158),
.B(n_1189),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1130),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1178),
.A2(n_1104),
.B1(n_1096),
.B2(n_1094),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1132),
.A2(n_1160),
.B(n_1189),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1079),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1079),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1134),
.A2(n_1160),
.B(n_1184),
.C(n_1140),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1143),
.B(n_1184),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1082),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1159),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1164),
.B(n_1174),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1179),
.B(n_1176),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1093),
.A2(n_1020),
.B1(n_1032),
.B2(n_1013),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1102),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1061),
.B(n_1013),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1076),
.B(n_1171),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1061),
.B(n_1013),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1058),
.A2(n_1063),
.B(n_1024),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1188),
.Y(n_1308)
);

AND2x6_ASAP7_75t_L g1309 ( 
.A(n_1125),
.B(n_1013),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1076),
.B(n_1171),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1084),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1076),
.B(n_1171),
.Y(n_1312)
);

AO32x1_ASAP7_75t_L g1313 ( 
.A1(n_1147),
.A2(n_1151),
.A3(n_1191),
.B1(n_1182),
.B2(n_740),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1076),
.B(n_1171),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_SL g1316 ( 
.A(n_1136),
.B(n_487),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1075),
.A2(n_1024),
.B(n_1016),
.C(n_1008),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1058),
.A2(n_1063),
.B(n_1024),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1045),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1076),
.B(n_1171),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1061),
.B(n_1013),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1058),
.A2(n_1063),
.B(n_1024),
.Y(n_1322)
);

BUFx12f_ASAP7_75t_L g1323 ( 
.A(n_1102),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1059),
.A2(n_1077),
.B(n_1052),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1090),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1043),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1150),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1061),
.B(n_1013),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1058),
.A2(n_1063),
.B(n_1024),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1188),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1058),
.A2(n_1063),
.B(n_1024),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_SL g1332 ( 
.A1(n_1075),
.A2(n_1024),
.B(n_1050),
.C(n_1152),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1078),
.B(n_887),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1042),
.A2(n_1020),
.B1(n_1032),
.B2(n_1013),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1058),
.A2(n_1063),
.B(n_1024),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1058),
.A2(n_1063),
.B(n_1024),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1206),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1197),
.A2(n_1234),
.B1(n_1243),
.B2(n_1198),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1213),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1240),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1302),
.B(n_1305),
.Y(n_1343)
);

OR2x6_ASAP7_75t_L g1344 ( 
.A(n_1231),
.B(n_1253),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1272),
.A2(n_1276),
.B(n_1262),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1335),
.A2(n_1211),
.B1(n_1203),
.B2(n_1202),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1239),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1302),
.B(n_1305),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1217),
.Y(n_1349)
);

BUFx8_ASAP7_75t_L g1350 ( 
.A(n_1323),
.Y(n_1350)
);

NOR2x1_ASAP7_75t_R g1351 ( 
.A(n_1258),
.B(n_1265),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1214),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1220),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1225),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1321),
.B(n_1328),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1197),
.A2(n_1212),
.B1(n_1321),
.B2(n_1328),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1335),
.A2(n_1242),
.B1(n_1309),
.B2(n_1231),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1272),
.A2(n_1276),
.B(n_1262),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1226),
.A2(n_1273),
.B(n_1222),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1202),
.A2(n_1233),
.B1(n_1309),
.B2(n_1254),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1233),
.A2(n_1309),
.B1(n_1215),
.B2(n_1300),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1228),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1333),
.A2(n_1215),
.B1(n_1208),
.B2(n_1251),
.Y(n_1363)
);

AO21x1_ASAP7_75t_L g1364 ( 
.A1(n_1317),
.A2(n_1208),
.B(n_1300),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_1301),
.Y(n_1365)
);

INVx4_ASAP7_75t_SL g1366 ( 
.A(n_1309),
.Y(n_1366)
);

INVx11_ASAP7_75t_L g1367 ( 
.A(n_1309),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1223),
.B(n_1246),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1326),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1236),
.A2(n_1223),
.B1(n_1201),
.B2(n_1311),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1317),
.A2(n_1219),
.B(n_1237),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1224),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1250),
.A2(n_1232),
.B1(n_1334),
.B2(n_1315),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1319),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1232),
.A2(n_1338),
.B1(n_1306),
.B2(n_1303),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1316),
.A2(n_1264),
.B1(n_1209),
.B2(n_1267),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1252),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1199),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1325),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1275),
.Y(n_1380)
);

INVx6_ASAP7_75t_L g1381 ( 
.A(n_1229),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1264),
.A2(n_1245),
.B1(n_1257),
.B2(n_1251),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_SL g1383 ( 
.A(n_1256),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1245),
.A2(n_1257),
.B1(n_1207),
.B2(n_1318),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1266),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1261),
.Y(n_1386)
);

BUFx12f_ASAP7_75t_L g1387 ( 
.A(n_1249),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1210),
.Y(n_1388)
);

INVx5_ASAP7_75t_L g1389 ( 
.A(n_1259),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1253),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1255),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1246),
.B(n_1229),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1199),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1230),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1332),
.B(n_1207),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1263),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1240),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1271),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1271),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1241),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1229),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1270),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1270),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1200),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1307),
.A2(n_1337),
.B1(n_1336),
.B2(n_1331),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1307),
.A2(n_1337),
.B1(n_1336),
.B2(n_1331),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1274),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1241),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1269),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1200),
.A2(n_1310),
.B1(n_1314),
.B2(n_1320),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1260),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1290),
.A2(n_1238),
.B(n_1244),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1260),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1221),
.B(n_1304),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1241),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1221),
.A2(n_1314),
.B1(n_1310),
.B2(n_1320),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1237),
.A2(n_1318),
.B(n_1329),
.Y(n_1417)
);

CKINVDCx6p67_ASAP7_75t_R g1418 ( 
.A(n_1268),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1304),
.B(n_1312),
.Y(n_1419)
);

AO21x1_ASAP7_75t_L g1420 ( 
.A1(n_1278),
.A2(n_1282),
.B(n_1329),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1247),
.B(n_1312),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1330),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1324),
.A2(n_1294),
.B(n_1248),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1285),
.Y(n_1424)
);

INVx5_ASAP7_75t_L g1425 ( 
.A(n_1259),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1277),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1277),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1280),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1281),
.B(n_1283),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1322),
.A2(n_1287),
.B1(n_1313),
.B2(n_1278),
.Y(n_1430)
);

INVx6_ASAP7_75t_L g1431 ( 
.A(n_1218),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1204),
.Y(n_1432)
);

INVx6_ASAP7_75t_L g1433 ( 
.A(n_1308),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1308),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1322),
.A2(n_1227),
.B(n_1205),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_SL g1436 ( 
.A1(n_1313),
.A2(n_1289),
.B1(n_1216),
.B2(n_1327),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1286),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1294),
.A2(n_1244),
.B(n_1238),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1247),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1313),
.A2(n_1227),
.B1(n_1205),
.B2(n_1248),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_L g1441 ( 
.A(n_1247),
.B(n_1292),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1297),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1293),
.A2(n_1235),
.B1(n_1284),
.B2(n_1296),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1296),
.Y(n_1444)
);

INVx3_ASAP7_75t_SL g1445 ( 
.A(n_1284),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1235),
.A2(n_1279),
.B(n_1299),
.Y(n_1446)
);

INVx6_ASAP7_75t_L g1447 ( 
.A(n_1284),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1288),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1295),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1298),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1288),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1291),
.A2(n_1016),
.B1(n_1025),
.B2(n_1008),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1204),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1226),
.A2(n_1059),
.B(n_1273),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1335),
.A2(n_1016),
.B1(n_1025),
.B2(n_1008),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1335),
.A2(n_1016),
.B1(n_1156),
.B2(n_1195),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1242),
.B(n_1195),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1450),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1343),
.B(n_1348),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1442),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1454),
.A2(n_1423),
.B(n_1359),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1454),
.A2(n_1423),
.B(n_1359),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1429),
.B(n_1409),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1438),
.A2(n_1417),
.B(n_1371),
.Y(n_1464)
);

BUFx2_ASAP7_75t_SL g1465 ( 
.A(n_1439),
.Y(n_1465)
);

CKINVDCx11_ASAP7_75t_R g1466 ( 
.A(n_1432),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1449),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1457),
.B(n_1411),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1402),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1455),
.B(n_1390),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1444),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1457),
.B(n_1413),
.Y(n_1473)
);

OAI21xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1346),
.A2(n_1456),
.B(n_1360),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1340),
.B(n_1346),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1403),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1437),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1398),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1420),
.A2(n_1438),
.B(n_1412),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1399),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1440),
.A2(n_1384),
.B(n_1405),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1377),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1456),
.A2(n_1452),
.B(n_1360),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1352),
.B(n_1374),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1366),
.B(n_1428),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1412),
.A2(n_1446),
.B(n_1364),
.Y(n_1486)
);

AO31x2_ASAP7_75t_L g1487 ( 
.A1(n_1451),
.A2(n_1395),
.A3(n_1426),
.B(n_1427),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1391),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1344),
.B(n_1361),
.Y(n_1489)
);

OAI21xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1382),
.A2(n_1367),
.B(n_1344),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1357),
.B(n_1382),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1447),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1384),
.B(n_1366),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1380),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1447),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1341),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1396),
.B(n_1347),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1366),
.B(n_1430),
.Y(n_1498)
);

AO21x1_ASAP7_75t_SL g1499 ( 
.A1(n_1443),
.A2(n_1406),
.B(n_1405),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1440),
.A2(n_1406),
.B(n_1443),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1435),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1370),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1381),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1349),
.Y(n_1504)
);

INVxp33_ASAP7_75t_L g1505 ( 
.A(n_1414),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1345),
.A2(n_1358),
.B(n_1428),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1372),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1353),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1354),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1369),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1386),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1368),
.B(n_1339),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1448),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1373),
.B(n_1368),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1393),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1445),
.B(n_1375),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1381),
.Y(n_1517)
);

BUFx2_ASAP7_75t_R g1518 ( 
.A(n_1453),
.Y(n_1518)
);

AOI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1363),
.A2(n_1376),
.B1(n_1416),
.B2(n_1424),
.C(n_1404),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1381),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1444),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1441),
.B(n_1392),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1378),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1436),
.B(n_1379),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1421),
.B(n_1392),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1421),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1392),
.B(n_1410),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1407),
.B(n_1419),
.Y(n_1528)
);

INVx2_ASAP7_75t_SL g1529 ( 
.A(n_1401),
.Y(n_1529)
);

INVx4_ASAP7_75t_L g1530 ( 
.A(n_1401),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1342),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1401),
.Y(n_1532)
);

NAND2x1_ASAP7_75t_L g1533 ( 
.A(n_1342),
.B(n_1397),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1418),
.B(n_1397),
.Y(n_1534)
);

NAND2x1p5_ASAP7_75t_L g1535 ( 
.A(n_1389),
.B(n_1425),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1475),
.B(n_1425),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1481),
.B(n_1408),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1470),
.B(n_1408),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1487),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1460),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1481),
.B(n_1408),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1481),
.B(n_1408),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1464),
.B(n_1418),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1506),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_L g1545 ( 
.A(n_1533),
.B(n_1472),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1481),
.B(n_1422),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1494),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1491),
.A2(n_1383),
.B1(n_1439),
.B2(n_1350),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1464),
.B(n_1422),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1491),
.A2(n_1383),
.B1(n_1350),
.B2(n_1365),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1500),
.B(n_1415),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1469),
.B(n_1385),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1469),
.B(n_1400),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1500),
.B(n_1400),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1460),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1476),
.B(n_1389),
.Y(n_1556)
);

AOI211x1_ASAP7_75t_SL g1557 ( 
.A1(n_1483),
.A2(n_1383),
.B(n_1350),
.C(n_1365),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1476),
.B(n_1434),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1489),
.B(n_1362),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1501),
.B(n_1486),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1486),
.B(n_1362),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1478),
.B(n_1434),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1477),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1471),
.B(n_1394),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1506),
.B(n_1388),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1486),
.B(n_1463),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1502),
.B(n_1431),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1478),
.B(n_1431),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1531),
.B(n_1432),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1480),
.B(n_1431),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1486),
.B(n_1433),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1463),
.B(n_1499),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1564),
.A2(n_1483),
.B1(n_1459),
.B2(n_1519),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1566),
.B(n_1477),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1547),
.B(n_1488),
.Y(n_1575)
);

OAI211xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1550),
.A2(n_1507),
.B(n_1513),
.C(n_1484),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1537),
.B(n_1513),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1547),
.B(n_1482),
.Y(n_1578)
);

OAI211xp5_ASAP7_75t_L g1579 ( 
.A1(n_1548),
.A2(n_1474),
.B(n_1490),
.C(n_1524),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1564),
.A2(n_1550),
.B1(n_1548),
.B2(n_1465),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1537),
.B(n_1493),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1569),
.A2(n_1474),
.B1(n_1527),
.B2(n_1493),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1563),
.B(n_1480),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1561),
.B(n_1540),
.Y(n_1584)
);

OAI221xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1543),
.A2(n_1490),
.B1(n_1561),
.B2(n_1572),
.C(n_1514),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1561),
.B(n_1467),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1541),
.B(n_1498),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1541),
.B(n_1498),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1541),
.B(n_1468),
.Y(n_1589)
);

AOI211xp5_ASAP7_75t_L g1590 ( 
.A1(n_1543),
.A2(n_1505),
.B(n_1497),
.C(n_1507),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1538),
.B(n_1458),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1542),
.B(n_1468),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1542),
.B(n_1473),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1538),
.A2(n_1465),
.B1(n_1521),
.B2(n_1472),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1559),
.B(n_1458),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1558),
.A2(n_1516),
.B1(n_1534),
.B2(n_1530),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1557),
.A2(n_1522),
.B(n_1516),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1569),
.A2(n_1522),
.B1(n_1526),
.B2(n_1532),
.Y(n_1598)
);

OA21x2_ASAP7_75t_L g1599 ( 
.A1(n_1544),
.A2(n_1461),
.B(n_1462),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1558),
.A2(n_1521),
.B1(n_1472),
.B2(n_1524),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1546),
.B(n_1479),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1562),
.A2(n_1496),
.B1(n_1523),
.B2(n_1518),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1546),
.B(n_1551),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1567),
.B(n_1517),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1543),
.A2(n_1528),
.B1(n_1515),
.B2(n_1525),
.C(n_1492),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1572),
.A2(n_1509),
.B1(n_1511),
.B2(n_1508),
.Y(n_1606)
);

OAI31xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1572),
.A2(n_1522),
.A3(n_1525),
.B(n_1512),
.Y(n_1607)
);

AOI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1536),
.A2(n_1511),
.B1(n_1504),
.B2(n_1508),
.C(n_1510),
.Y(n_1608)
);

OAI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1557),
.A2(n_1520),
.B1(n_1529),
.B2(n_1517),
.C(n_1495),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1569),
.A2(n_1522),
.B1(n_1503),
.B2(n_1530),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_SL g1611 ( 
.A1(n_1536),
.A2(n_1485),
.B(n_1535),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1567),
.A2(n_1503),
.B1(n_1530),
.B2(n_1520),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1555),
.B(n_1510),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1545),
.B(n_1529),
.Y(n_1614)
);

NAND4xp25_ASAP7_75t_L g1615 ( 
.A(n_1552),
.B(n_1568),
.C(n_1570),
.D(n_1553),
.Y(n_1615)
);

NOR3xp33_ASAP7_75t_L g1616 ( 
.A(n_1568),
.B(n_1503),
.C(n_1530),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1599),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1584),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1603),
.B(n_1601),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1613),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1601),
.B(n_1544),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1613),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1599),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1583),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1574),
.B(n_1560),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1583),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1586),
.B(n_1560),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1586),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1581),
.B(n_1549),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1615),
.B(n_1560),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1577),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1589),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1599),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1599),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1581),
.B(n_1577),
.Y(n_1635)
);

NAND4xp25_ASAP7_75t_L g1636 ( 
.A(n_1573),
.B(n_1570),
.C(n_1552),
.D(n_1556),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1575),
.B(n_1571),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1575),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1587),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1615),
.B(n_1539),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1554),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1620),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1620),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1620),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1630),
.B(n_1591),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1630),
.B(n_1578),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1630),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1639),
.B(n_1607),
.Y(n_1648)
);

NOR2xp67_ASAP7_75t_L g1649 ( 
.A(n_1640),
.B(n_1611),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1622),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1622),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1622),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1624),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1634),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1634),
.Y(n_1655)
);

INVxp67_ASAP7_75t_SL g1656 ( 
.A(n_1640),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1633),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_1640),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1625),
.B(n_1592),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1638),
.B(n_1593),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1633),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1624),
.Y(n_1662)
);

OR2x6_ASAP7_75t_L g1663 ( 
.A(n_1617),
.B(n_1611),
.Y(n_1663)
);

NOR2x1p5_ASAP7_75t_L g1664 ( 
.A(n_1636),
.B(n_1595),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1636),
.B(n_1590),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1623),
.B(n_1573),
.C(n_1590),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1607),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1639),
.B(n_1614),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1634),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1588),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1624),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1638),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1631),
.B(n_1565),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1631),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1634),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1619),
.B(n_1629),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1625),
.B(n_1627),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1638),
.A2(n_1579),
.B1(n_1580),
.B2(n_1576),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1632),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1626),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1642),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1666),
.A2(n_1580),
.B1(n_1600),
.B2(n_1594),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1646),
.B(n_1627),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1642),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1643),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1643),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1644),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1672),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1668),
.Y(n_1689)
);

OAI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1666),
.A2(n_1665),
.B(n_1678),
.Y(n_1690)
);

OAI31xp33_ASAP7_75t_L g1691 ( 
.A1(n_1664),
.A2(n_1602),
.A3(n_1585),
.B(n_1600),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1644),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1648),
.B(n_1621),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1650),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1650),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1678),
.A2(n_1602),
.B(n_1594),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1663),
.Y(n_1697)
);

OAI31xp33_ASAP7_75t_L g1698 ( 
.A1(n_1664),
.A2(n_1596),
.A3(n_1605),
.B(n_1606),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1646),
.B(n_1627),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1651),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1656),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1648),
.B(n_1621),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1658),
.B(n_1637),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1647),
.B(n_1637),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1649),
.A2(n_1604),
.B(n_1608),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1621),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1651),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1652),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1645),
.B(n_1625),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1663),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1667),
.B(n_1619),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1645),
.B(n_1628),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1670),
.B(n_1641),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1668),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1660),
.B(n_1466),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1676),
.B(n_1635),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1670),
.B(n_1641),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1676),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1654),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1649),
.B(n_1635),
.Y(n_1720)
);

NAND2x1p5_ASAP7_75t_L g1721 ( 
.A(n_1668),
.B(n_1545),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1652),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1660),
.B(n_1641),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1701),
.B(n_1677),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1688),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1692),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1697),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1712),
.B(n_1677),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1719),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1689),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1714),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1692),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1719),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1718),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1720),
.B(n_1663),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1690),
.B(n_1668),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1688),
.Y(n_1737)
);

OR2x6_ASAP7_75t_L g1738 ( 
.A(n_1696),
.B(n_1663),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1715),
.A2(n_1663),
.B1(n_1679),
.B2(n_1674),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1694),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1711),
.B(n_1674),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1705),
.B(n_1453),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1691),
.A2(n_1582),
.B1(n_1616),
.B2(n_1673),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1682),
.B(n_1628),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1694),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1695),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1718),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1695),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1703),
.B(n_1351),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1698),
.B(n_1635),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1700),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1711),
.B(n_1618),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1697),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1693),
.B(n_1673),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1712),
.B(n_1659),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1683),
.B(n_1659),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1700),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1693),
.B(n_1673),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_L g1759 ( 
.A(n_1710),
.B(n_1653),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1727),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1753),
.B(n_1702),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1742),
.B(n_1749),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1741),
.B(n_1702),
.Y(n_1763)
);

OAI21xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1738),
.A2(n_1720),
.B(n_1706),
.Y(n_1764)
);

OAI32xp33_ASAP7_75t_L g1765 ( 
.A1(n_1736),
.A2(n_1721),
.A3(n_1704),
.B1(n_1706),
.B2(n_1699),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1730),
.B(n_1716),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1727),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1738),
.A2(n_1710),
.B1(n_1699),
.B2(n_1683),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1748),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1731),
.B(n_1716),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1750),
.B(n_1713),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1748),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1738),
.A2(n_1597),
.B1(n_1612),
.B2(n_1606),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1741),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1725),
.B(n_1717),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1759),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1759),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1739),
.A2(n_1721),
.B(n_1684),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1754),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1754),
.B(n_1721),
.Y(n_1780)
);

OAI32xp33_ASAP7_75t_L g1781 ( 
.A1(n_1744),
.A2(n_1709),
.A3(n_1633),
.B1(n_1661),
.B2(n_1657),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1748),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1726),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1758),
.B(n_1737),
.Y(n_1784)
);

AND2x4_ASAP7_75t_SL g1785 ( 
.A(n_1735),
.B(n_1673),
.Y(n_1785)
);

OAI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1738),
.A2(n_1709),
.B1(n_1707),
.B2(n_1686),
.C(n_1687),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_SL g1787 ( 
.A(n_1762),
.B(n_1738),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1760),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1761),
.B(n_1724),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1767),
.B(n_1737),
.Y(n_1790)
);

NOR2xp67_ASAP7_75t_L g1791 ( 
.A(n_1764),
.B(n_1728),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1760),
.B(n_1737),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1760),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1774),
.B(n_1743),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1774),
.B(n_1724),
.Y(n_1795)
);

NOR2x1_ASAP7_75t_L g1796 ( 
.A(n_1776),
.B(n_1726),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1784),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1784),
.B(n_1728),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1763),
.B(n_1758),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1784),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1766),
.B(n_1755),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1775),
.B(n_1755),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1769),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1784),
.B(n_1734),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1769),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1785),
.Y(n_1806)
);

NAND4xp75_ASAP7_75t_L g1807 ( 
.A(n_1791),
.B(n_1796),
.C(n_1764),
.D(n_1792),
.Y(n_1807)
);

AOI221x1_ASAP7_75t_L g1808 ( 
.A1(n_1788),
.A2(n_1776),
.B1(n_1777),
.B2(n_1782),
.C(n_1772),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1794),
.A2(n_1765),
.B1(n_1786),
.B2(n_1778),
.C(n_1768),
.Y(n_1809)
);

OAI211xp5_ASAP7_75t_L g1810 ( 
.A1(n_1790),
.A2(n_1765),
.B(n_1777),
.C(n_1781),
.Y(n_1810)
);

AOI221x1_ASAP7_75t_L g1811 ( 
.A1(n_1804),
.A2(n_1782),
.B1(n_1772),
.B2(n_1783),
.C(n_1770),
.Y(n_1811)
);

OAI321xp33_ASAP7_75t_L g1812 ( 
.A1(n_1798),
.A2(n_1773),
.A3(n_1779),
.B1(n_1780),
.B2(n_1771),
.C(n_1763),
.Y(n_1812)
);

AOI211xp5_ASAP7_75t_L g1813 ( 
.A1(n_1787),
.A2(n_1781),
.B(n_1773),
.C(n_1779),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1795),
.B(n_1783),
.C(n_1780),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1797),
.A2(n_1800),
.B1(n_1793),
.B2(n_1806),
.C(n_1789),
.Y(n_1815)
);

AOI211xp5_ASAP7_75t_L g1816 ( 
.A1(n_1806),
.A2(n_1793),
.B(n_1801),
.C(n_1802),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1802),
.A2(n_1805),
.B1(n_1803),
.B2(n_1799),
.C(n_1734),
.Y(n_1817)
);

O2A1O1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1799),
.A2(n_1745),
.B(n_1757),
.C(n_1740),
.Y(n_1818)
);

NOR4xp25_ASAP7_75t_L g1819 ( 
.A(n_1815),
.B(n_1734),
.C(n_1747),
.D(n_1745),
.Y(n_1819)
);

NOR3xp33_ASAP7_75t_L g1820 ( 
.A(n_1816),
.B(n_1747),
.C(n_1740),
.Y(n_1820)
);

OAI322xp33_ASAP7_75t_L g1821 ( 
.A1(n_1818),
.A2(n_1747),
.A3(n_1757),
.B1(n_1732),
.B2(n_1751),
.C1(n_1746),
.C2(n_1733),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1808),
.Y(n_1822)
);

NOR3xp33_ASAP7_75t_L g1823 ( 
.A(n_1809),
.B(n_1746),
.C(n_1732),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1807),
.A2(n_1785),
.B1(n_1735),
.B2(n_1751),
.Y(n_1824)
);

NOR2x1p5_ASAP7_75t_SL g1825 ( 
.A(n_1812),
.B(n_1733),
.Y(n_1825)
);

AOI211x1_ASAP7_75t_L g1826 ( 
.A1(n_1810),
.A2(n_1752),
.B(n_1708),
.C(n_1722),
.Y(n_1826)
);

NOR2x1p5_ASAP7_75t_SL g1827 ( 
.A(n_1811),
.B(n_1733),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1819),
.A2(n_1813),
.B(n_1814),
.C(n_1817),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1822),
.A2(n_1735),
.B(n_1756),
.Y(n_1829)
);

AOI32xp33_ASAP7_75t_L g1830 ( 
.A1(n_1823),
.A2(n_1735),
.A3(n_1729),
.B1(n_1756),
.B2(n_1623),
.Y(n_1830)
);

NAND4xp75_ASAP7_75t_L g1831 ( 
.A(n_1827),
.B(n_1825),
.C(n_1826),
.D(n_1824),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_L g1832 ( 
.A(n_1820),
.B(n_1729),
.C(n_1722),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1831),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1829),
.B(n_1681),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1832),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1828),
.A2(n_1708),
.B1(n_1685),
.B2(n_1387),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1830),
.A2(n_1387),
.B1(n_1723),
.B2(n_1680),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1832),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1834),
.Y(n_1839)
);

NAND5xp2_ASAP7_75t_L g1840 ( 
.A(n_1836),
.B(n_1821),
.C(n_1597),
.D(n_1610),
.E(n_1598),
.Y(n_1840)
);

NAND3x1_ASAP7_75t_L g1841 ( 
.A(n_1835),
.B(n_1661),
.C(n_1657),
.Y(n_1841)
);

XNOR2x1_ASAP7_75t_L g1842 ( 
.A(n_1833),
.B(n_1535),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1838),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1839),
.B(n_1837),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1843),
.Y(n_1845)
);

AND3x1_ASAP7_75t_L g1846 ( 
.A(n_1840),
.B(n_1661),
.C(n_1657),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1845),
.Y(n_1847)
);

OAI221xp5_ASAP7_75t_L g1848 ( 
.A1(n_1847),
.A2(n_1842),
.B1(n_1844),
.B2(n_1846),
.C(n_1841),
.Y(n_1848)
);

BUFx2_ASAP7_75t_L g1849 ( 
.A(n_1848),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1848),
.A2(n_1657),
.B1(n_1661),
.B2(n_1623),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1849),
.A2(n_1654),
.B(n_1675),
.C(n_1655),
.Y(n_1851)
);

OAI22x1_ASAP7_75t_L g1852 ( 
.A1(n_1850),
.A2(n_1654),
.B1(n_1675),
.B2(n_1655),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1852),
.A2(n_1655),
.B1(n_1675),
.B2(n_1669),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1851),
.Y(n_1854)
);

AOI21xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1854),
.A2(n_1535),
.B(n_1669),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1855),
.A2(n_1853),
.B(n_1669),
.Y(n_1856)
);

OAI221xp5_ASAP7_75t_R g1857 ( 
.A1(n_1856),
.A2(n_1617),
.B1(n_1671),
.B2(n_1662),
.C(n_1653),
.Y(n_1857)
);

AOI211xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1609),
.B(n_1680),
.C(n_1662),
.Y(n_1858)
);


endmodule