module real_jpeg_723_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_88, n_11, n_14, n_7, n_3, n_87, n_5, n_4, n_1, n_89, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_88;
input n_11;
input n_14;
input n_7;
input n_3;
input n_87;
input n_5;
input n_4;
input n_1;
input n_89;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_0),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_1),
.A2(n_17),
.B1(n_23),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_5),
.A2(n_55),
.B1(n_58),
.B2(n_69),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_5),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_87),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_8),
.B(n_10),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_20),
.B1(n_52),
.B2(n_53),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_11),
.A2(n_52),
.B1(n_71),
.B2(n_78),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_15),
.B(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_15),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_16),
.B(n_88),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_89),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_17),
.A2(n_23),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_17),
.A2(n_46),
.B(n_48),
.Y(n_45)
);

AOI221xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_54),
.B1(n_70),
.B2(n_79),
.C(n_84),
.Y(n_18)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_49),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_73),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_31),
.C(n_39),
.Y(n_38)
);

OAI211xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_34),
.B(n_37),
.C(n_45),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B(n_30),
.Y(n_27)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_38),
.B(n_42),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_29),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_31),
.A2(n_35),
.B(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_35),
.A2(n_38),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_74),
.C(n_77),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_65),
.B(n_68),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);


endmodule