module fake_aes_1357_n_694 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_694);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_694;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g80 ( .A(n_8), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_20), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_65), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_71), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_24), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_63), .Y(n_85) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_4), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_2), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_40), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_77), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_64), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_15), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_37), .Y(n_92) );
BUFx3_ASAP7_75t_L g93 ( .A(n_33), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_21), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_49), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_47), .Y(n_96) );
OR2x2_ASAP7_75t_L g97 ( .A(n_43), .B(n_17), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_5), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_27), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_21), .Y(n_100) );
BUFx10_ASAP7_75t_L g101 ( .A(n_79), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_30), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_51), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_42), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_78), .Y(n_105) );
INVxp33_ASAP7_75t_L g106 ( .A(n_15), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_44), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_53), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_34), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_18), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_12), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_55), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_35), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_38), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_23), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_3), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_25), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_17), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_41), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_11), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_1), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_7), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_76), .B(n_28), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_57), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_5), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_9), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_99), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_96), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_99), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_111), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_111), .Y(n_132) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_82), .A2(n_36), .B(n_74), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_89), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_103), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_101), .B(n_0), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_104), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_80), .Y(n_138) );
NOR2xp33_ASAP7_75t_R g139 ( .A(n_103), .B(n_32), .Y(n_139) );
OR2x6_ASAP7_75t_L g140 ( .A(n_86), .B(n_1), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_81), .B(n_2), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_122), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_80), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_124), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_109), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_108), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_101), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_100), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_81), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_101), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_101), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_97), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_87), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_88), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_126), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_87), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_119), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_106), .B(n_3), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_93), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_93), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_115), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_115), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_83), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_97), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_91), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_91), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_159), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_148), .B(n_94), .Y(n_172) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_141), .B(n_125), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_148), .B(n_94), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_159), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_148), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_141), .B(n_125), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_133), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_144), .B(n_118), .Y(n_183) );
AO22x2_ASAP7_75t_L g184 ( .A1(n_141), .A2(n_82), .B1(n_84), .B2(n_85), .Y(n_184) );
AND2x6_ASAP7_75t_L g185 ( .A(n_134), .B(n_84), .Y(n_185) );
NAND2xp33_ASAP7_75t_SL g186 ( .A(n_153), .B(n_110), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_133), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_137), .B(n_120), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_128), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_151), .B(n_117), .Y(n_190) );
OAI221xp5_ASAP7_75t_L g191 ( .A1(n_168), .A2(n_110), .B1(n_121), .B2(n_120), .C(n_118), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_164), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_133), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_151), .B(n_121), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_167), .B(n_105), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_133), .Y(n_197) );
INVxp67_ASAP7_75t_SL g198 ( .A(n_161), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_147), .B(n_116), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_166), .Y(n_201) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_128), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_166), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_162), .B(n_117), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
OAI22xp33_ASAP7_75t_L g208 ( .A1(n_140), .A2(n_98), .B1(n_116), .B2(n_114), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_162), .B(n_102), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_156), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_163), .B(n_102), .Y(n_212) );
BUFx4f_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_163), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_167), .B(n_105), .Y(n_215) );
AO22x2_ASAP7_75t_L g216 ( .A1(n_136), .A2(n_107), .B1(n_114), .B2(n_113), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_158), .B(n_98), .Y(n_217) );
BUFx4f_ASAP7_75t_L g218 ( .A(n_140), .Y(n_218) );
NAND3x1_ASAP7_75t_L g219 ( .A(n_140), .B(n_113), .C(n_112), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_168), .B(n_112), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_157), .B(n_107), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_169), .B(n_85), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_157), .B(n_92), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_170), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_160), .B(n_92), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_139), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_160), .A2(n_90), .B1(n_95), .B2(n_123), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_130), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_130), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_135), .Y(n_231) );
OAI21xp33_ASAP7_75t_SL g232 ( .A1(n_172), .A2(n_135), .B(n_154), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_213), .B(n_95), .Y(n_233) );
NOR2xp33_ASAP7_75t_R g234 ( .A(n_213), .B(n_145), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_189), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_213), .B(n_95), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_171), .Y(n_237) );
INVx5_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_175), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_175), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_176), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_213), .A2(n_145), .B(n_95), .C(n_149), .Y(n_244) );
NOR3xp33_ASAP7_75t_SL g245 ( .A(n_186), .B(n_146), .C(n_132), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_198), .B(n_131), .Y(n_246) );
AND2x6_ASAP7_75t_SL g247 ( .A(n_215), .B(n_142), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_220), .B(n_146), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_171), .Y(n_249) );
NOR3xp33_ASAP7_75t_SL g250 ( .A(n_191), .B(n_4), .C(n_6), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_218), .Y(n_251) );
INVx4_ASAP7_75t_L g252 ( .A(n_218), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_200), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_218), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_218), .Y(n_256) );
BUFx8_ASAP7_75t_SL g257 ( .A(n_189), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_172), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_174), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_184), .A2(n_95), .B1(n_7), .B2(n_8), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_174), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_210), .B(n_6), .Y(n_262) );
BUFx12f_ASAP7_75t_L g263 ( .A(n_230), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_200), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_231), .B(n_48), .Y(n_266) );
NOR2xp67_ASAP7_75t_L g267 ( .A(n_202), .B(n_9), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_200), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_205), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_230), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_173), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_212), .B(n_10), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_231), .B(n_196), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_190), .B(n_10), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_205), .Y(n_275) );
NOR3xp33_ASAP7_75t_SL g276 ( .A(n_208), .B(n_11), .C(n_12), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_230), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_183), .B(n_13), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_184), .A2(n_13), .B1(n_14), .B2(n_16), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_206), .B(n_14), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_207), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_173), .B(n_56), .Y(n_284) );
INVx5_ASAP7_75t_L g285 ( .A(n_185), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_206), .B(n_16), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_219), .Y(n_287) );
INVx5_ASAP7_75t_L g288 ( .A(n_185), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_207), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_201), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_201), .Y(n_291) );
NOR2xp33_ASAP7_75t_R g292 ( .A(n_229), .B(n_18), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_185), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_201), .Y(n_294) );
INVx4_ASAP7_75t_L g295 ( .A(n_173), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_184), .A2(n_19), .B1(n_20), .B2(n_22), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_240), .A2(n_187), .B(n_197), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g298 ( .A(n_295), .B(n_178), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_293), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_271), .A2(n_180), .B1(n_184), .B2(n_219), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_295), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_295), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_241), .Y(n_303) );
NOR2xp33_ASAP7_75t_SL g304 ( .A(n_293), .B(n_180), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_279), .A2(n_185), .B1(n_195), .B2(n_216), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_235), .B(n_195), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_258), .B(n_259), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_242), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_252), .B(n_229), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_238), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_243), .Y(n_311) );
BUFx12f_ASAP7_75t_L g312 ( .A(n_263), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_271), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_261), .B(n_214), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_241), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_254), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_277), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_263), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_249), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_264), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_252), .B(n_229), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_269), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_246), .B(n_183), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_275), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_249), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_283), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_252), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_273), .B(n_209), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_292), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_289), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_256), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_287), .A2(n_185), .B1(n_216), .B2(n_180), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_270), .B(n_223), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_280), .A2(n_185), .B1(n_216), .B2(n_211), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_238), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_238), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_246), .B(n_223), .Y(n_338) );
CKINVDCx12_ASAP7_75t_R g339 ( .A(n_257), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_238), .Y(n_340) );
BUFx10_ASAP7_75t_L g341 ( .A(n_251), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_238), .Y(n_342) );
BUFx12f_ASAP7_75t_L g343 ( .A(n_247), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_237), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_248), .B(n_229), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_246), .B(n_226), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_237), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_237), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g350 ( .A(n_301), .B(n_285), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_324), .A2(n_232), .B1(n_257), .B2(n_255), .Y(n_351) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_300), .A2(n_234), .B1(n_251), .B2(n_216), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_308), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_301), .B(n_255), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_311), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_301), .Y(n_357) );
NOR3xp33_ASAP7_75t_SL g358 ( .A(n_339), .B(n_224), .C(n_244), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_324), .A2(n_214), .B1(n_234), .B2(n_216), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_317), .B(n_285), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_338), .A2(n_250), .B1(n_296), .B2(n_260), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_318), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_303), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_302), .B(n_285), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_310), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_302), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_345), .A2(n_222), .B(n_204), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_306), .A2(n_267), .B1(n_227), .B2(n_188), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_338), .A2(n_188), .B1(n_245), .B2(n_217), .C(n_199), .Y(n_369) );
NAND2xp33_ASAP7_75t_R g370 ( .A(n_318), .B(n_276), .Y(n_370) );
INVx2_ASAP7_75t_SL g371 ( .A(n_302), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_305), .A2(n_244), .B1(n_227), .B2(n_272), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_303), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_306), .B(n_217), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_317), .Y(n_375) );
OR2x6_ASAP7_75t_L g376 ( .A(n_312), .B(n_233), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_333), .A2(n_262), .B1(n_274), .B2(n_286), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_334), .B(n_221), .Y(n_378) );
AOI21xp5_ASAP7_75t_SL g379 ( .A1(n_300), .A2(n_284), .B(n_266), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_315), .Y(n_380) );
INVx6_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_369), .A2(n_343), .B1(n_346), .B2(n_322), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_351), .A2(n_346), .B1(n_314), .B2(n_335), .C(n_329), .Y(n_383) );
OAI211xp5_ASAP7_75t_SL g384 ( .A1(n_362), .A2(n_228), .B(n_281), .C(n_335), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_361), .A2(n_343), .B1(n_322), .B2(n_330), .Y(n_385) );
CKINVDCx11_ASAP7_75t_R g386 ( .A(n_357), .Y(n_386) );
OAI211xp5_ASAP7_75t_L g387 ( .A1(n_368), .A2(n_307), .B(n_334), .C(n_233), .Y(n_387) );
OAI22xp33_ASAP7_75t_SL g388 ( .A1(n_361), .A2(n_330), .B1(n_304), .B2(n_302), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_353), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_353), .B(n_320), .Y(n_390) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_379), .A2(n_284), .B(n_297), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_352), .A2(n_320), .B1(n_323), .B2(n_325), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_370), .A2(n_304), .B1(n_343), .B2(n_312), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_359), .A2(n_323), .B1(n_325), .B2(n_331), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_378), .A2(n_327), .B1(n_331), .B2(n_332), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_375), .A2(n_312), .B1(n_329), .B2(n_311), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_354), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_377), .A2(n_321), .B(n_309), .Y(n_398) );
BUFx4f_ASAP7_75t_SL g399 ( .A(n_357), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_354), .Y(n_400) );
AO221x2_ASAP7_75t_L g401 ( .A1(n_356), .A2(n_327), .B1(n_316), .B2(n_339), .C(n_19), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_374), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_374), .B(n_316), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_349), .Y(n_404) );
OR2x2_ASAP7_75t_SL g405 ( .A(n_381), .B(n_315), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_356), .B(n_307), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_349), .A2(n_313), .B1(n_298), .B2(n_326), .Y(n_407) );
INVx4_ASAP7_75t_L g408 ( .A(n_357), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_367), .A2(n_358), .B1(n_372), .B2(n_379), .C(n_178), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_401), .A2(n_367), .B1(n_309), .B2(n_321), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_406), .B(n_199), .Y(n_411) );
AO21x2_ASAP7_75t_L g412 ( .A1(n_409), .A2(n_182), .B(n_194), .Y(n_412) );
AOI211xp5_ASAP7_75t_L g413 ( .A1(n_396), .A2(n_309), .B(n_321), .C(n_236), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_389), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_404), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_402), .Y(n_416) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_404), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_401), .A2(n_321), .B1(n_309), .B2(n_376), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_406), .B(n_209), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_389), .Y(n_420) );
OAI33xp33_ASAP7_75t_L g421 ( .A1(n_393), .A2(n_179), .A3(n_177), .B1(n_203), .B2(n_181), .B3(n_193), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_386), .Y(n_422) );
OAI221xp5_ASAP7_75t_SL g423 ( .A1(n_382), .A2(n_376), .B1(n_207), .B2(n_211), .C(n_221), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_399), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_397), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_383), .A2(n_381), .B1(n_376), .B2(n_366), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_403), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_392), .A2(n_381), .B1(n_376), .B2(n_380), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_388), .A2(n_366), .B(n_371), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_400), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g432 ( .A1(n_395), .A2(n_381), .B1(n_371), .B2(n_357), .Y(n_432) );
OAI211xp5_ASAP7_75t_L g433 ( .A1(n_385), .A2(n_236), .B(n_203), .C(n_193), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_400), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_405), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_390), .B(n_363), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_403), .B(n_181), .C(n_179), .D(n_177), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_405), .B(n_363), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_401), .B(n_357), .C(n_373), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_387), .B(n_192), .C(n_225), .D(n_355), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_401), .B(n_380), .Y(n_442) );
INVx4_ASAP7_75t_L g443 ( .A(n_408), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_408), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_428), .B(n_394), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_437), .B(n_408), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_414), .B(n_373), .Y(n_447) );
OAI211xp5_ASAP7_75t_SL g448 ( .A1(n_416), .A2(n_398), .B(n_192), .C(n_225), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_414), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_413), .B(n_384), .C(n_201), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_422), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_420), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_443), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_436), .B(n_388), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_427), .A2(n_355), .B1(n_391), .B2(n_407), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_417), .Y(n_456) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_443), .B(n_391), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_420), .B(n_391), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_413), .B(n_440), .C(n_410), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_425), .B(n_319), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_425), .A2(n_348), .A3(n_347), .B1(n_360), .B2(n_225), .B3(n_182), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_437), .B(n_315), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_442), .B(n_365), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_415), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_431), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_436), .B(n_355), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_431), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_434), .B(n_355), .Y(n_468) );
OAI21xp33_ASAP7_75t_L g469 ( .A1(n_440), .A2(n_201), .B(n_298), .Y(n_469) );
OAI31xp33_ASAP7_75t_SL g470 ( .A1(n_429), .A2(n_364), .A3(n_319), .B(n_326), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_434), .B(n_319), .Y(n_471) );
AOI21xp5_ASAP7_75t_SL g472 ( .A1(n_424), .A2(n_313), .B(n_350), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_443), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_442), .B(n_365), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_426), .Y(n_475) );
INVxp33_ASAP7_75t_L g476 ( .A(n_438), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_426), .B(n_326), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_423), .A2(n_298), .B1(n_328), .B2(n_365), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_415), .B(n_365), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_411), .B(n_201), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_424), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_444), .B(n_365), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_419), .B(n_347), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_439), .Y(n_484) );
AND2x4_ASAP7_75t_SL g485 ( .A(n_444), .B(n_364), .Y(n_485) );
NAND2xp33_ASAP7_75t_SL g486 ( .A(n_435), .B(n_364), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_418), .B(n_194), .C(n_182), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_412), .Y(n_488) );
INVxp33_ASAP7_75t_L g489 ( .A(n_438), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_439), .Y(n_490) );
OAI31xp33_ASAP7_75t_L g491 ( .A1(n_432), .A2(n_328), .A3(n_350), .B(n_348), .Y(n_491) );
AOI211xp5_ASAP7_75t_L g492 ( .A1(n_435), .A2(n_328), .B(n_187), .C(n_197), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_412), .B(n_26), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_481), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_449), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_458), .B(n_412), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_484), .B(n_422), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_452), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_464), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_458), .B(n_430), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_490), .B(n_441), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_453), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_465), .Y(n_503) );
NAND2xp33_ASAP7_75t_R g504 ( .A(n_453), .B(n_29), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_476), .A2(n_421), .B1(n_328), .B2(n_344), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_464), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_467), .B(n_433), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_475), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_463), .B(n_31), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_445), .B(n_197), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_463), .B(n_39), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_453), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_446), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_466), .B(n_194), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_481), .Y(n_515) );
NOR2x1_ASAP7_75t_L g516 ( .A(n_472), .B(n_457), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_446), .Y(n_517) );
NAND2xp33_ASAP7_75t_R g518 ( .A(n_493), .B(n_45), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_456), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_447), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_447), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_454), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_451), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_460), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_463), .B(n_46), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_460), .B(n_187), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_474), .B(n_50), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_477), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_462), .B(n_350), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_477), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_479), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_474), .B(n_52), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_462), .B(n_344), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_468), .B(n_344), .Y(n_534) );
AND4x1_ASAP7_75t_L g535 ( .A(n_470), .B(n_341), .C(n_58), .D(n_59), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_473), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_471), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_474), .B(n_54), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_473), .B(n_344), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_478), .A2(n_340), .B(n_336), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_476), .B(n_341), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_489), .B(n_341), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_488), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_488), .B(n_60), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_482), .B(n_61), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_479), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_482), .B(n_62), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_493), .B(n_66), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_493), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_455), .B(n_67), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_489), .B(n_68), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_459), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_499), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_513), .B(n_485), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_519), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_495), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_495), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_517), .B(n_485), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_536), .Y(n_559) );
OAI21xp33_ASAP7_75t_SL g560 ( .A1(n_516), .A2(n_491), .B(n_486), .Y(n_560) );
AOI21xp33_ASAP7_75t_L g561 ( .A1(n_552), .A2(n_480), .B(n_450), .Y(n_561) );
AOI22x1_ASAP7_75t_L g562 ( .A1(n_494), .A2(n_486), .B1(n_469), .B2(n_492), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_515), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_498), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_522), .B(n_483), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_498), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_523), .Y(n_567) );
AOI32xp33_ASAP7_75t_L g568 ( .A1(n_552), .A2(n_448), .A3(n_461), .B1(n_487), .B2(n_342), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_503), .Y(n_569) );
OAI21xp33_ASAP7_75t_SL g570 ( .A1(n_516), .A2(n_336), .B(n_340), .Y(n_570) );
AOI21xp33_ASAP7_75t_SL g571 ( .A1(n_504), .A2(n_69), .B(n_70), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_499), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_503), .Y(n_573) );
OAI21xp33_ASAP7_75t_L g574 ( .A1(n_522), .A2(n_290), .B(n_253), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_520), .B(n_72), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_512), .A2(n_502), .B(n_540), .Y(n_576) );
OR3x2_ASAP7_75t_L g577 ( .A(n_497), .B(n_73), .C(n_75), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_518), .A2(n_299), .B1(n_342), .B2(n_288), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_524), .B(n_239), .Y(n_579) );
OAI32xp33_ASAP7_75t_L g580 ( .A1(n_502), .A2(n_342), .A3(n_265), .B1(n_278), .B2(n_291), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_497), .B(n_239), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_520), .B(n_239), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_524), .B(n_239), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_508), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_541), .A2(n_299), .B1(n_310), .B2(n_337), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_542), .A2(n_299), .B1(n_310), .B2(n_337), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_512), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_521), .B(n_268), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_529), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_551), .B(n_268), .C(n_282), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_521), .B(n_268), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_537), .B(n_268), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_508), .Y(n_593) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_501), .A2(n_282), .B(n_294), .Y(n_594) );
AND3x2_ASAP7_75t_L g595 ( .A(n_548), .B(n_291), .C(n_299), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_546), .B(n_282), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_506), .Y(n_597) );
NAND2x1_ASAP7_75t_L g598 ( .A(n_502), .B(n_337), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_550), .A2(n_299), .B1(n_282), .B2(n_294), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_537), .B(n_294), .Y(n_600) );
OAI21xp5_ASAP7_75t_SL g601 ( .A1(n_535), .A2(n_310), .B(n_337), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_548), .A2(n_285), .B(n_288), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_506), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_528), .B(n_265), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_563), .B(n_507), .Y(n_605) );
NAND2xp33_ASAP7_75t_SL g606 ( .A(n_554), .B(n_549), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_555), .B(n_500), .Y(n_607) );
INVxp33_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
NAND2xp33_ASAP7_75t_SL g609 ( .A(n_558), .B(n_549), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_560), .A2(n_550), .B(n_505), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_555), .B(n_496), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_559), .B(n_531), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_603), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_565), .B(n_528), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_556), .B(n_530), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_567), .Y(n_616) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_603), .Y(n_617) );
XNOR2x2_ASAP7_75t_L g618 ( .A(n_576), .B(n_527), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_577), .A2(n_530), .B1(n_531), .B2(n_532), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_589), .B(n_509), .Y(n_620) );
NAND2x1_ASAP7_75t_L g621 ( .A(n_584), .B(n_593), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_570), .B(n_543), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_598), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_557), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_571), .A2(n_545), .B(n_547), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_578), .B(n_544), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_564), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_566), .B(n_510), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_587), .B(n_527), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_601), .A2(n_525), .B(n_538), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_569), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_573), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_561), .B(n_545), .C(n_547), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_553), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_572), .B(n_529), .Y(n_635) );
XOR2x2_ASAP7_75t_L g636 ( .A(n_595), .B(n_577), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_572), .B(n_544), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_581), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_597), .Y(n_639) );
AOI321xp33_ASAP7_75t_L g640 ( .A1(n_605), .A2(n_581), .A3(n_575), .B1(n_532), .B2(n_538), .C(n_525), .Y(n_640) );
OAI332xp33_ASAP7_75t_L g641 ( .A1(n_616), .A2(n_578), .A3(n_597), .B1(n_533), .B2(n_534), .B3(n_604), .C1(n_585), .C2(n_586), .Y(n_641) );
XNOR2xp5_ASAP7_75t_L g642 ( .A(n_636), .B(n_595), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_621), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g644 ( .A1(n_608), .A2(n_602), .B(n_599), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_624), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_627), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_607), .B(n_588), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_631), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_632), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_630), .A2(n_590), .B1(n_511), .B2(n_509), .Y(n_650) );
NAND4xp25_ASAP7_75t_L g651 ( .A(n_610), .B(n_568), .C(n_594), .D(n_511), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_608), .A2(n_605), .B1(n_614), .B2(n_609), .C(n_606), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_613), .Y(n_653) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_622), .B(n_539), .Y(n_654) );
OAI21xp33_ASAP7_75t_L g655 ( .A1(n_611), .A2(n_574), .B(n_596), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_613), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_615), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_617), .B(n_583), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_622), .Y(n_659) );
OA22x2_ASAP7_75t_L g660 ( .A1(n_619), .A2(n_591), .B1(n_582), .B2(n_579), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_657), .B(n_638), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_659), .A2(n_609), .B1(n_606), .B2(n_633), .C(n_612), .Y(n_662) );
AOI21xp33_ASAP7_75t_L g663 ( .A1(n_642), .A2(n_623), .B(n_628), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_656), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_652), .A2(n_636), .B1(n_625), .B2(n_626), .C(n_618), .Y(n_665) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_654), .B(n_623), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_660), .A2(n_629), .B1(n_626), .B2(n_620), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_641), .A2(n_635), .B1(n_634), .B2(n_639), .C(n_637), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_653), .B(n_639), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_651), .A2(n_623), .B1(n_539), .B2(n_533), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_644), .A2(n_580), .B(n_592), .C(n_600), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_651), .B(n_514), .C(n_526), .D(n_265), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_645), .Y(n_673) );
NAND5xp2_ASAP7_75t_L g674 ( .A(n_644), .B(n_285), .C(n_288), .D(n_299), .E(n_310), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_650), .A2(n_310), .B1(n_337), .B2(n_288), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_643), .B(n_278), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_646), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_648), .Y(n_678) );
AO221x1_ASAP7_75t_L g679 ( .A1(n_640), .A2(n_641), .B1(n_649), .B2(n_655), .C(n_658), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_647), .A2(n_659), .B1(n_652), .B2(n_641), .C(n_608), .Y(n_680) );
AOI221x1_ASAP7_75t_L g681 ( .A1(n_663), .A2(n_679), .B1(n_672), .B2(n_661), .C(n_676), .Y(n_681) );
INVx1_ASAP7_75t_SL g682 ( .A(n_664), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_665), .A2(n_680), .B1(n_662), .B2(n_670), .C(n_667), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_673), .Y(n_684) );
AOI22xp33_ASAP7_75t_R g685 ( .A1(n_678), .A2(n_677), .B1(n_666), .B2(n_675), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_682), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_684), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_683), .A2(n_668), .B1(n_676), .B2(n_669), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_686), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_687), .Y(n_690) );
BUFx3_ASAP7_75t_L g691 ( .A(n_690), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_689), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_692), .A2(n_688), .B1(n_681), .B2(n_685), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_693), .A2(n_691), .B1(n_681), .B2(n_671), .C(n_674), .Y(n_694) );
endmodule