module fake_ariane_1470_n_761 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_761);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_761;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_48),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_39),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_20),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_46),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_67),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_74),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_52),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_71),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_6),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_108),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_2),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_9),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_77),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_8),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_49),
.Y(n_174)
);

BUFx2_ASAP7_75t_SL g175 ( 
.A(n_55),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_51),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_94),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_92),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_90),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_112),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_86),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_30),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_63),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_78),
.B(n_50),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_1),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_85),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_13),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_122),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_27),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_82),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_8),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_64),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_87),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_45),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_98),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_32),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_88),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_0),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_0),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_167),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_1),
.Y(n_219)
);

OAI22x1_ASAP7_75t_SL g220 ( 
.A1(n_189),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_3),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_4),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_161),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_155),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_158),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_169),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_187),
.B(n_175),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_159),
.B(n_5),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_160),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_5),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_193),
.B(n_6),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_170),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_163),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_231),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_212),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_211),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_240),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_239),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_217),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_239),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_R g265 ( 
.A(n_216),
.B(n_185),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_239),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_216),
.B(n_174),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_239),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_228),
.Y(n_274)
);

NOR2x1p5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_165),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_234),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_234),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_226),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_R g279 ( 
.A(n_218),
.B(n_178),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_225),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_225),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_223),
.B(n_195),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_225),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_225),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_209),
.B(n_166),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_224),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_209),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_229),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_222),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_237),
.Y(n_294)
);

AOI221xp5_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_243),
.B1(n_238),
.B2(n_220),
.C(n_244),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_229),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_238),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_249),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_227),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_236),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_213),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_213),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_235),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_258),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_259),
.B(n_206),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_248),
.B(n_235),
.Y(n_315)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_267),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_229),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_229),
.Y(n_319)
);

OR2x2_ASAP7_75t_SL g320 ( 
.A(n_248),
.B(n_208),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_265),
.B(n_219),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_L g324 ( 
.A(n_268),
.B(n_221),
.C(n_243),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_257),
.B(n_230),
.Y(n_325)
);

NAND2x1p5_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_230),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_285),
.B(n_230),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_275),
.A2(n_232),
.B1(n_230),
.B2(n_201),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_257),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_232),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_265),
.B(n_232),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_251),
.Y(n_334)
);

NAND2x1_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_232),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_279),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_209),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_251),
.B(n_209),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_246),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_263),
.B(n_210),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_269),
.B(n_10),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_263),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_271),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_269),
.B(n_210),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_252),
.B(n_204),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_250),
.B(n_168),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_280),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_282),
.B(n_210),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_262),
.B(n_171),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_282),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_291),
.B(n_210),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_271),
.B(n_177),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_179),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_295),
.A2(n_194),
.B1(n_184),
.B2(n_190),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_317),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_297),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_300),
.B(n_253),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_309),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_316),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_301),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_307),
.B(n_181),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_330),
.B(n_192),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

OR2x6_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_247),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_315),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_11),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_330),
.B(n_196),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

BUFx4f_ASAP7_75t_L g374 ( 
.A(n_316),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_321),
.B(n_271),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_324),
.A2(n_215),
.B1(n_12),
.B2(n_13),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_313),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_293),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_339),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_293),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_326),
.B(n_11),
.Y(n_382)
);

BUFx12f_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_302),
.B(n_215),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_347),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_325),
.B(n_329),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_303),
.B(n_12),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_294),
.B(n_326),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_324),
.B(n_14),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_298),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_299),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_345),
.B(n_14),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_322),
.B(n_15),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_16),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_341),
.B(n_17),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_332),
.B(n_153),
.Y(n_400)
);

AND3x2_ASAP7_75t_SL g401 ( 
.A(n_314),
.B(n_18),
.C(n_19),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_305),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_306),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_344),
.A2(n_350),
.B1(n_353),
.B2(n_346),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_310),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_318),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_349),
.B(n_21),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_312),
.B(n_22),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_343),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_319),
.B(n_23),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_328),
.B(n_152),
.Y(n_414)
);

AND3x1_ASAP7_75t_L g415 ( 
.A(n_331),
.B(n_24),
.C(n_25),
.Y(n_415)
);

AND2x2_ASAP7_75t_SL g416 ( 
.A(n_343),
.B(n_26),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_338),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_343),
.B(n_28),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_355),
.B(n_29),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_374),
.B(n_354),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_354),
.Y(n_424)
);

NOR3xp33_ASAP7_75t_L g425 ( 
.A(n_359),
.B(n_337),
.C(n_351),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_361),
.B(n_351),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_417),
.A2(n_31),
.B(n_33),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_381),
.B(n_34),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_35),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_374),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_370),
.A2(n_151),
.B1(n_37),
.B2(n_38),
.Y(n_432)
);

OAI22x1_ASAP7_75t_L g433 ( 
.A1(n_357),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_358),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_370),
.B(n_42),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_422),
.A2(n_43),
.B(n_44),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_SL g438 ( 
.A(n_363),
.B(n_47),
.Y(n_438)
);

A2O1A1Ixp33_ASAP7_75t_L g439 ( 
.A1(n_387),
.A2(n_357),
.B(n_376),
.C(n_377),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_362),
.Y(n_440)
);

AOI21x1_ASAP7_75t_L g441 ( 
.A1(n_389),
.A2(n_53),
.B(n_54),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_356),
.B(n_56),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_380),
.B(n_416),
.Y(n_443)
);

A2O1A1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_376),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_60),
.Y(n_445)
);

AO21x1_ASAP7_75t_L g446 ( 
.A1(n_389),
.A2(n_61),
.B(n_62),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_369),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_368),
.A2(n_65),
.B(n_66),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_399),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_449)
);

CKINVDCx8_ASAP7_75t_R g450 ( 
.A(n_369),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_373),
.A2(n_72),
.B(n_73),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_399),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_453)
);

NOR3xp33_ASAP7_75t_L g454 ( 
.A(n_366),
.B(n_80),
.C(n_83),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_402),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_396),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_407),
.B(n_84),
.Y(n_458)
);

O2A1O1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_390),
.A2(n_89),
.B(n_91),
.C(n_93),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_SL g460 ( 
.A(n_397),
.B(n_95),
.C(n_96),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_360),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_403),
.A2(n_365),
.B1(n_379),
.B2(n_367),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_382),
.Y(n_463)
);

AND2x6_ASAP7_75t_L g464 ( 
.A(n_420),
.B(n_97),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_418),
.A2(n_419),
.B(n_394),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_358),
.B(n_99),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_394),
.A2(n_372),
.B(n_400),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_367),
.A2(n_379),
.B1(n_386),
.B2(n_413),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_404),
.B(n_100),
.Y(n_469)
);

O2A1O1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_393),
.A2(n_101),
.B(n_102),
.C(n_103),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_406),
.B(n_105),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_414),
.A2(n_106),
.B1(n_111),
.B2(n_113),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_385),
.B(n_114),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_375),
.A2(n_115),
.B(n_116),
.Y(n_475)
);

A2O1A1Ixp33_ASAP7_75t_L g476 ( 
.A1(n_421),
.A2(n_412),
.B(n_392),
.C(n_408),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_383),
.B(n_150),
.Y(n_477)
);

O2A1O1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_395),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_408),
.A2(n_120),
.B(n_121),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_431),
.Y(n_480)
);

BUFx2_ASAP7_75t_R g481 ( 
.A(n_450),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_456),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_467),
.A2(n_415),
.B(n_384),
.Y(n_484)
);

AOI22x1_ASAP7_75t_L g485 ( 
.A1(n_465),
.A2(n_395),
.B1(n_411),
.B2(n_398),
.Y(n_485)
);

AO21x2_ASAP7_75t_L g486 ( 
.A1(n_476),
.A2(n_415),
.B(n_401),
.Y(n_486)
);

OR2x6_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_398),
.Y(n_487)
);

BUFx12f_ASAP7_75t_L g488 ( 
.A(n_447),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_430),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_398),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_431),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_440),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_457),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

BUFx2_ASAP7_75t_SL g496 ( 
.A(n_451),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_411),
.Y(n_497)
);

BUFx4f_ASAP7_75t_SL g498 ( 
.A(n_474),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_426),
.B(n_411),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_437),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_461),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_441),
.A2(n_405),
.B(n_410),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_443),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_464),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_473),
.B(n_410),
.Y(n_505)
);

BUFx2_ASAP7_75t_SL g506 ( 
.A(n_464),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_435),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_439),
.B(n_410),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_429),
.B(n_410),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_479),
.A2(n_123),
.B(n_125),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_468),
.Y(n_512)
);

BUFx12f_ASAP7_75t_L g513 ( 
.A(n_477),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_455),
.B(n_126),
.Y(n_514)
);

INVx5_ASAP7_75t_SL g515 ( 
.A(n_432),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_445),
.Y(n_516)
);

AO21x2_ASAP7_75t_L g517 ( 
.A1(n_442),
.A2(n_127),
.B(n_128),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_434),
.B(n_129),
.Y(n_518)
);

AOI21x1_ASAP7_75t_L g519 ( 
.A1(n_462),
.A2(n_134),
.B(n_136),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_428),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_460),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_458),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_469),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_425),
.A2(n_142),
.B(n_143),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_449),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_523),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_493),
.B(n_495),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_524),
.A2(n_444),
.B(n_446),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_504),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_483),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_482),
.Y(n_531)
);

AO21x2_ASAP7_75t_L g532 ( 
.A1(n_502),
.A2(n_454),
.B(n_472),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_489),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_509),
.B(n_433),
.Y(n_534)
);

OA21x2_ASAP7_75t_L g535 ( 
.A1(n_484),
.A2(n_448),
.B(n_452),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_453),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g537 ( 
.A1(n_484),
.A2(n_427),
.B(n_436),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_515),
.A2(n_466),
.B1(n_423),
.B2(n_438),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_512),
.Y(n_539)
);

HB1xp67_ASAP7_75t_SL g540 ( 
.A(n_481),
.Y(n_540)
);

AO21x1_ASAP7_75t_L g541 ( 
.A1(n_508),
.A2(n_459),
.B(n_470),
.Y(n_541)
);

BUFx8_ASAP7_75t_L g542 ( 
.A(n_488),
.Y(n_542)
);

BUFx2_ASAP7_75t_SL g543 ( 
.A(n_504),
.Y(n_543)
);

INVx6_ASAP7_75t_L g544 ( 
.A(n_480),
.Y(n_544)
);

AO21x1_ASAP7_75t_L g545 ( 
.A1(n_525),
.A2(n_478),
.B(n_475),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_494),
.Y(n_546)
);

BUFx4f_ASAP7_75t_SL g547 ( 
.A(n_488),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_483),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_492),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

OA21x2_ASAP7_75t_L g551 ( 
.A1(n_502),
.A2(n_144),
.B(n_145),
.Y(n_551)
);

INVx6_ASAP7_75t_L g552 ( 
.A(n_480),
.Y(n_552)
);

AO21x1_ASAP7_75t_SL g553 ( 
.A1(n_510),
.A2(n_146),
.B(n_147),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_501),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_497),
.B(n_148),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_513),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_493),
.B(n_495),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_518),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_512),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_497),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_518),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_515),
.A2(n_487),
.B1(n_499),
.B2(n_521),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_485),
.A2(n_149),
.B(n_519),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_SL g564 ( 
.A1(n_515),
.A2(n_513),
.B1(n_498),
.B2(n_507),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_493),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_520),
.A2(n_516),
.B(n_521),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_495),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_511),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_526),
.B(n_503),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_529),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_531),
.B(n_497),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_530),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_496),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_539),
.Y(n_574)
);

OR2x6_ASAP7_75t_L g575 ( 
.A(n_543),
.B(n_487),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_543),
.B(n_487),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_539),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_560),
.B(n_487),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_529),
.B(n_560),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_564),
.B(n_515),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_559),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_542),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_534),
.A2(n_486),
.B1(n_506),
.B2(n_521),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_540),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_SL g585 ( 
.A1(n_534),
.A2(n_486),
.B1(n_505),
.B2(n_517),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_558),
.B(n_561),
.Y(n_586)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_563),
.A2(n_566),
.B(n_568),
.Y(n_587)
);

NAND2x1p5_ASAP7_75t_L g588 ( 
.A(n_529),
.B(n_480),
.Y(n_588)
);

BUFx4f_ASAP7_75t_L g589 ( 
.A(n_529),
.Y(n_589)
);

AND2x4_ASAP7_75t_SL g590 ( 
.A(n_529),
.B(n_491),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_530),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_559),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_R g593 ( 
.A(n_556),
.B(n_505),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_533),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_542),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_SL g596 ( 
.A(n_556),
.B(n_514),
.C(n_522),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_R g597 ( 
.A(n_555),
.B(n_505),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_546),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_536),
.A2(n_486),
.B1(n_562),
.B2(n_528),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_548),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_550),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_SL g602 ( 
.A1(n_528),
.A2(n_517),
.B1(n_520),
.B2(n_511),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_555),
.B(n_491),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_536),
.B(n_500),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_565),
.B(n_491),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_565),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_550),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_542),
.Y(n_608)
);

AND2x2_ASAP7_75t_SL g609 ( 
.A(n_538),
.B(n_551),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_SL g610 ( 
.A(n_547),
.B(n_500),
.C(n_490),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_527),
.B(n_557),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_SL g612 ( 
.A1(n_527),
.A2(n_520),
.B(n_490),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_554),
.B(n_500),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_594),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_574),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_598),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_586),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_574),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_580),
.A2(n_528),
.B1(n_541),
.B2(n_532),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_571),
.B(n_552),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_577),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_609),
.A2(n_541),
.B1(n_532),
.B2(n_517),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_604),
.B(n_567),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_577),
.Y(n_624)
);

AOI21xp33_ASAP7_75t_L g625 ( 
.A1(n_602),
.A2(n_532),
.B(n_551),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_569),
.B(n_554),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_600),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_599),
.B(n_567),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_581),
.Y(n_629)
);

OR2x2_ASAP7_75t_SL g630 ( 
.A(n_584),
.B(n_552),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_606),
.B(n_567),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_600),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_573),
.B(n_565),
.Y(n_633)
);

AOI221xp5_ASAP7_75t_L g634 ( 
.A1(n_596),
.A2(n_545),
.B1(n_568),
.B2(n_500),
.C(n_557),
.Y(n_634)
);

NAND2x1p5_ASAP7_75t_L g635 ( 
.A(n_589),
.B(n_551),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_585),
.B(n_570),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_570),
.B(n_557),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_601),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_611),
.B(n_576),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_613),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_603),
.B(n_544),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_612),
.A2(n_545),
.B(n_537),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_601),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_611),
.B(n_563),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_581),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_589),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_587),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_575),
.B(n_553),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_623),
.B(n_582),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_614),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_648),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_623),
.B(n_595),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_616),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_621),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_617),
.B(n_592),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_626),
.B(n_583),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_615),
.B(n_612),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_615),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_618),
.Y(n_659)
);

INVx5_ASAP7_75t_L g660 ( 
.A(n_648),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_620),
.B(n_605),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_605),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_618),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_624),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_624),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_627),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_620),
.B(n_590),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_628),
.B(n_553),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_640),
.B(n_591),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_633),
.B(n_572),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_636),
.B(n_576),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_631),
.B(n_607),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_632),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_668),
.A2(n_622),
.B(n_619),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_653),
.B(n_645),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_653),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_654),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_662),
.B(n_636),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_654),
.B(n_619),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_662),
.B(n_628),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_660),
.B(n_648),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_651),
.B(n_642),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_651),
.B(n_637),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_663),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_663),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_651),
.B(n_637),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_655),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_676),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_677),
.B(n_650),
.Y(n_689)
);

AOI32xp33_ASAP7_75t_L g690 ( 
.A1(n_679),
.A2(n_668),
.A3(n_622),
.B1(n_671),
.B2(n_673),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_687),
.B(n_672),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_675),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_684),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_679),
.B(n_666),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_674),
.B(n_634),
.C(n_657),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_685),
.B(n_670),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_681),
.Y(n_697)
);

OR4x1_ASAP7_75t_L g698 ( 
.A(n_688),
.B(n_664),
.C(n_665),
.D(n_682),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_695),
.A2(n_674),
.B(n_625),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_692),
.Y(n_700)
);

NAND2x1p5_ASAP7_75t_L g701 ( 
.A(n_697),
.B(n_660),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_697),
.B(n_681),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_698),
.Y(n_703)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_699),
.A2(n_690),
.B(n_694),
.C(n_656),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_700),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_699),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_702),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_701),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_706),
.B(n_608),
.Y(n_709)
);

CKINVDCx14_ASAP7_75t_R g710 ( 
.A(n_707),
.Y(n_710)
);

OAI221xp5_ASAP7_75t_L g711 ( 
.A1(n_704),
.A2(n_701),
.B1(n_691),
.B2(n_689),
.C(n_696),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_705),
.Y(n_712)
);

OAI211xp5_ASAP7_75t_L g713 ( 
.A1(n_710),
.A2(n_703),
.B(n_709),
.C(n_711),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_712),
.B(n_708),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_711),
.A2(n_693),
.B(n_652),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_714),
.Y(n_716)
);

AOI21xp33_ASAP7_75t_SL g717 ( 
.A1(n_713),
.A2(n_681),
.B(n_649),
.Y(n_717)
);

NAND3xp33_ASAP7_75t_L g718 ( 
.A(n_715),
.B(n_682),
.C(n_610),
.Y(n_718)
);

OAI21xp5_ASAP7_75t_L g719 ( 
.A1(n_713),
.A2(n_678),
.B(n_680),
.Y(n_719)
);

NOR2x1_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_646),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_718),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_719),
.Y(n_722)
);

NOR2x1_ASAP7_75t_L g723 ( 
.A(n_717),
.B(n_646),
.Y(n_723)
);

AO22x2_ASAP7_75t_L g724 ( 
.A1(n_716),
.A2(n_671),
.B1(n_639),
.B2(n_686),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_716),
.B(n_683),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_716),
.A2(n_660),
.B1(n_630),
.B2(n_661),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_720),
.B(n_660),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_R g728 ( 
.A1(n_722),
.A2(n_659),
.B1(n_658),
.B2(n_638),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_724),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_721),
.B(n_667),
.C(n_641),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_725),
.B(n_723),
.Y(n_731)
);

AOI211xp5_ASAP7_75t_L g732 ( 
.A1(n_726),
.A2(n_671),
.B(n_644),
.C(n_639),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_720),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_720),
.B(n_544),
.Y(n_734)
);

AOI221xp5_ASAP7_75t_SL g735 ( 
.A1(n_731),
.A2(n_647),
.B1(n_659),
.B2(n_658),
.C(n_643),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_733),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_729),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_734),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_727),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_730),
.A2(n_575),
.B(n_588),
.Y(n_740)
);

AOI221xp5_ASAP7_75t_L g741 ( 
.A1(n_732),
.A2(n_635),
.B1(n_644),
.B2(n_647),
.C(n_669),
.Y(n_741)
);

NAND4xp25_ASAP7_75t_L g742 ( 
.A(n_728),
.B(n_593),
.C(n_597),
.D(n_647),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_736),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_737),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_738),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_739),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_742),
.Y(n_747)
);

XOR2xp5_ASAP7_75t_L g748 ( 
.A(n_740),
.B(n_578),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_741),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_744),
.A2(n_735),
.B1(n_544),
.B2(n_552),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_746),
.Y(n_751)
);

AOI31xp33_ASAP7_75t_L g752 ( 
.A1(n_745),
.A2(n_635),
.A3(n_639),
.B(n_544),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_743),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_751),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_753),
.A2(n_747),
.B1(n_749),
.B2(n_748),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_754),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_755),
.B(n_750),
.Y(n_757)
);

AOI21xp33_ASAP7_75t_L g758 ( 
.A1(n_756),
.A2(n_752),
.B(n_644),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_758),
.A2(n_757),
.B1(n_552),
.B2(n_537),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_759),
.B(n_579),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_760),
.A2(n_535),
.B1(n_537),
.B2(n_629),
.Y(n_761)
);


endmodule