module fake_jpeg_10784_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_30),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_71),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_73),
.B1(n_62),
.B2(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_0),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_4),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_54),
.Y(n_87)
);

CKINVDCx6p67_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_62),
.B(n_60),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_92),
.B1(n_101),
.B2(n_17),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_65),
.B1(n_45),
.B2(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_52),
.B1(n_53),
.B2(n_61),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_97),
.B1(n_100),
.B2(n_105),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_52),
.A3(n_60),
.B1(n_59),
.B2(n_51),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_50),
.B1(n_49),
.B2(n_64),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_4),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_22),
.B1(n_42),
.B2(n_40),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_5),
.B(n_7),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_14),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_101),
.B1(n_102),
.B2(n_34),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_113),
.B(n_114),
.Y(n_126)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_116),
.B1(n_114),
.B2(n_107),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_18),
.C(n_21),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_115),
.C(n_38),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_25),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_104),
.C(n_106),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_33),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_118),
.B1(n_112),
.B2(n_110),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_118),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_108),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_123),
.B(n_124),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_129),
.C(n_121),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_125),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_116),
.B(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_122),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_122),
.Y(n_134)
);

INVxp33_ASAP7_75t_SL g137 ( 
.A(n_134),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_136),
.B(n_133),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_131),
.C(n_137),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_140),
.Y(n_141)
);


endmodule