module real_jpeg_4269_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_1),
.A2(n_91),
.B1(n_92),
.B2(n_95),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_1),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_1),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_2),
.A2(n_23),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_2),
.A2(n_44),
.B1(n_49),
.B2(n_52),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_2),
.A2(n_44),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_2),
.A2(n_44),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_2),
.A2(n_223),
.B(n_226),
.C(n_229),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_2),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_2),
.B(n_139),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_2),
.B(n_266),
.C(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_2),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_2),
.B(n_71),
.C(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_2),
.B(n_25),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_3),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_3),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_3),
.A2(n_71),
.B1(n_112),
.B2(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_4),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_4),
.A2(n_22),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_4),
.A2(n_22),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_4),
.A2(n_22),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_5),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_5),
.Y(n_111)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_7),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_8),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_8),
.Y(n_228)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_11),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_11),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_207),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_206),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_188),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_15),
.B(n_188),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_151),
.C(n_169),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_16),
.B(n_151),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_87),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_46),
.B1(n_47),
.B2(n_86),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_18),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_18),
.B(n_47),
.C(n_87),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_18),
.B(n_201),
.C(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_18),
.A2(n_86),
.B1(n_201),
.B2(n_305),
.Y(n_329)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_24),
.B1(n_40),
.B2(n_45),
.Y(n_18)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_19),
.A2(n_24),
.B1(n_40),
.B2(n_45),
.Y(n_187)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_23),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_24),
.A2(n_40),
.B(n_45),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_25)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_44),
.A2(n_49),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_46),
.A2(n_47),
.B1(n_172),
.B2(n_260),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_46),
.B(n_260),
.C(n_282),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_46),
.A2(n_47),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_47),
.B(n_187),
.C(n_315),
.Y(n_333)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_55),
.B1(n_69),
.B2(n_80),
.Y(n_47)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_48),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_48),
.A2(n_55),
.B1(n_69),
.B2(n_80),
.Y(n_201)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_55),
.B(n_69),
.Y(n_186)
);

NAND2x1_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_69),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_66),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_69),
.Y(n_275)
);

AOI22x1_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_73),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_85),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_119),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_88),
.A2(n_119),
.B1(n_120),
.B2(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_88),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_97),
.B1(n_106),
.B2(n_116),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_90),
.A2(n_175),
.B(n_178),
.Y(n_174)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_95),
.Y(n_250)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_96),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_97),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_97),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_98),
.A2(n_180),
.B1(n_232),
.B2(n_237),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_98),
.A2(n_176),
.B1(n_180),
.B2(n_232),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_105),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_113),
.Y(n_267)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_115),
.Y(n_233)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_119),
.A2(n_120),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_119),
.A2(n_120),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_120),
.B(n_231),
.C(n_274),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_120),
.B(n_297),
.C(n_299),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_128),
.B1(n_144),
.B2(n_145),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_139),
.Y(n_173)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_128),
.B(n_144),
.Y(n_316)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_129),
.A2(n_139),
.B1(n_154),
.B2(n_199),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_133),
.B1(n_136),
.B2(n_138),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AO22x1_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_154),
.B(n_161),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_146),
.B(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_163),
.B2(n_168),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_163),
.Y(n_195)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_160),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_162),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_163),
.A2(n_168),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_164),
.B(n_180),
.Y(n_290)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_184),
.C(n_187),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_215),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_172),
.A2(n_260),
.B1(n_261),
.B2(n_268),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_172),
.A2(n_174),
.B1(n_260),
.B2(n_332),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_174),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_184),
.A2(n_187),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_187),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_187),
.A2(n_216),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_204),
.B2(n_205),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_196),
.B1(n_197),
.B2(n_203),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_201),
.B(n_202),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_201),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_201),
.A2(n_301),
.B1(n_302),
.B2(n_305),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_201),
.Y(n_305)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_240),
.B(n_344),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_210),
.B(n_212),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_218),
.C(n_220),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_213),
.A2(n_214),
.B1(n_218),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_218),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_220),
.B(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_221),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_222),
.A2(n_230),
.B1(n_231),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_222),
.Y(n_323)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_230),
.A2(n_231),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_255),
.Y(n_256)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_325),
.B(n_341),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_309),
.B(n_324),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_294),
.B(n_308),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_279),
.B(n_293),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_270),
.B(n_278),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_257),
.B(n_269),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_254),
.B(n_256),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_253),
.A2(n_258),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_259),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_258),
.B(n_303),
.C(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_277),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_277),
.Y(n_278)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_281),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_292),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_290),
.B2(n_291),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_291),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_290),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_307),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_307),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_299),
.B1(n_300),
.B2(n_306),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_311),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_320),
.C(n_321),
.Y(n_334)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2x1_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_335),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_334),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_334),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_328),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_333),
.C(n_337),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_335),
.A2(n_342),
.B(n_343),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_336),
.B(n_338),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);


endmodule