module fake_jpeg_3146_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_54),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_53),
.Y(n_56)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_41),
.C(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_47),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_43),
.B1(n_46),
.B2(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_53),
.A2(n_42),
.B1(n_45),
.B2(n_35),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_52),
.B1(n_36),
.B2(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_49),
.B1(n_53),
.B2(n_52),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_59),
.B1(n_40),
.B2(n_4),
.Y(n_86)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_1),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_72),
.B1(n_59),
.B2(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_43),
.B(n_46),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_60),
.A3(n_40),
.B1(n_2),
.B2(n_4),
.Y(n_80)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_89),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_68),
.B(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_2),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_75),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_29),
.B(n_28),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_70),
.B(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_100),
.B1(n_101),
.B2(n_11),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_95),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_66),
.B(n_89),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_102),
.B(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_1),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_6),
.C(n_8),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_6),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_19),
.C(n_7),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_82),
.C(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_103),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_82),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_108),
.C(n_113),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_77),
.B(n_10),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_9),
.B(n_10),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_114),
.B1(n_101),
.B2(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_9),
.C(n_11),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_116),
.B(n_117),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_113),
.A3(n_108),
.B1(n_114),
.B2(n_15),
.C1(n_12),
.C2(n_17),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_107),
.C(n_110),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_122),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_122),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_125),
.B(n_115),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_119),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C(n_13),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_16),
.Y(n_130)
);


endmodule