module fake_jpeg_743_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_52),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_49),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_69),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_66),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_43),
.B1(n_45),
.B2(n_51),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_45),
.B1(n_47),
.B2(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_81),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_82),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_57),
.B(n_51),
.C(n_40),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_39),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_42),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_41),
.B1(n_67),
.B2(n_47),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_72),
.B1(n_78),
.B2(n_44),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_41),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_47),
.B1(n_44),
.B2(n_15),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_108),
.B1(n_98),
.B2(n_7),
.Y(n_121)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_105),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_1),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_109),
.Y(n_126)
);

NOR4xp25_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_18),
.C(n_35),
.D(n_34),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_6),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_36),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_122),
.B1(n_127),
.B2(n_108),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_10),
.C(n_11),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_21),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_126),
.B(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_104),
.B1(n_114),
.B2(n_22),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_16),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_116),
.B(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_133),
.C(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_137),
.Y(n_139)
);

AOI321xp33_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_118),
.A3(n_120),
.B1(n_119),
.B2(n_124),
.C(n_32),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_118),
.B(n_136),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_139),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_29),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_24),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_25),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_144),
.Y(n_145)
);


endmodule