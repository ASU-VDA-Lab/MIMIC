module fake_jpeg_14421_n_453 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_453);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_453;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_4),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_16),
.B(n_15),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_47),
.B(n_52),
.Y(n_143)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_49),
.A2(n_22),
.B1(n_26),
.B2(n_20),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_67),
.Y(n_99)
);

AND2x6_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_0),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_55),
.B(n_39),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_10),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_88),
.Y(n_111)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_21),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_73),
.A2(n_34),
.B1(n_17),
.B2(n_32),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_79),
.Y(n_110)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_10),
.B(n_1),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_80),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_27),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_39),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_91),
.Y(n_116)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g145 ( 
.A(n_90),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_105),
.B(n_114),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_52),
.A2(n_42),
.B1(n_28),
.B2(n_23),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_115),
.A2(n_29),
.B1(n_25),
.B2(n_18),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_138),
.Y(n_154)
);

CKINVDCx12_ASAP7_75t_R g118 ( 
.A(n_57),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_51),
.B(n_35),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_119),
.B(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_35),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_33),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_123),
.B(n_125),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_73),
.B1(n_115),
.B2(n_143),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_33),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_30),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_134),
.B(n_136),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_50),
.B(n_30),
.Y(n_136)
);

CKINVDCx12_ASAP7_75t_R g137 ( 
.A(n_83),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_54),
.B(n_34),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_17),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_64),
.B(n_22),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_89),
.B1(n_91),
.B2(n_46),
.Y(n_177)
);

BUFx16f_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_147),
.A2(n_31),
.B(n_8),
.C(n_9),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_77),
.Y(n_149)
);

NAND2x1_ASAP7_75t_L g205 ( 
.A(n_149),
.B(n_101),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_141),
.A2(n_32),
.B1(n_69),
.B2(n_24),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_150),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_151),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_80),
.B1(n_25),
.B2(n_29),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_SL g215 ( 
.A(n_153),
.B(n_182),
.Y(n_215)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_155),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_92),
.A2(n_87),
.B1(n_90),
.B2(n_63),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_177),
.B1(n_104),
.B2(n_127),
.Y(n_213)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_158),
.Y(n_246)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_159),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_24),
.B1(n_26),
.B2(n_23),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_162),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_68),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_186),
.B1(n_199),
.B2(n_200),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_95),
.B(n_93),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_168),
.B(n_192),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

BUFx2_ASAP7_75t_SL g203 ( 
.A(n_171),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_98),
.A2(n_24),
.B1(n_23),
.B2(n_29),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_110),
.B(n_42),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_178),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_100),
.B(n_86),
.C(n_81),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_193),
.C(n_131),
.Y(n_229)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_124),
.A2(n_25),
.B(n_18),
.C(n_6),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_184),
.Y(n_223)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

BUFx24_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_116),
.A2(n_74),
.B1(n_66),
.B2(n_61),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_130),
.B(n_3),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_189),
.Y(n_220)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_194),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_120),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_113),
.B(n_78),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_60),
.C(n_31),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_94),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_120),
.A2(n_31),
.B1(n_6),
.B2(n_7),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_8),
.B1(n_9),
.B2(n_160),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_113),
.B(n_5),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_146),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_142),
.A2(n_31),
.B1(n_8),
.B2(n_9),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_106),
.A2(n_31),
.B1(n_8),
.B2(n_9),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_222),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_106),
.B1(n_142),
.B2(n_132),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_206),
.A2(n_208),
.B1(n_213),
.B2(n_226),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_108),
.B1(n_132),
.B2(n_126),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_216),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_153),
.A2(n_126),
.B1(n_104),
.B2(n_108),
.Y(n_208)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_163),
.A3(n_179),
.B1(n_174),
.B2(n_157),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_212),
.A2(n_164),
.B(n_161),
.C(n_189),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_163),
.A2(n_128),
.B1(n_97),
.B2(n_122),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_101),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_193),
.C(n_152),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_221),
.B(n_238),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_154),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_180),
.A2(n_128),
.B1(n_97),
.B2(n_122),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_229),
.B(n_187),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_151),
.B1(n_172),
.B2(n_190),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_182),
.A2(n_152),
.B(n_165),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_191),
.B(n_169),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_148),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_178),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_245),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_184),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_155),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_149),
.B(n_198),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_247),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_197),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_249),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_183),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_210),
.Y(n_250)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_251),
.B(n_273),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_245),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_253),
.B(n_254),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_181),
.Y(n_254)
);

INVx4_ASAP7_75t_SL g255 ( 
.A(n_209),
.Y(n_255)
);

INVx11_ASAP7_75t_L g317 ( 
.A(n_255),
.Y(n_317)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_257),
.Y(n_295)
);

BUFx12_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_258),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_259),
.A2(n_263),
.B(n_282),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_274),
.C(n_280),
.Y(n_308)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_170),
.B(n_173),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_264),
.A2(n_271),
.B1(n_281),
.B2(n_209),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_223),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_266),
.B(n_268),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_158),
.Y(n_268)
);

OR2x6_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_233),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_225),
.A2(n_208),
.B1(n_206),
.B2(n_226),
.Y(n_271)
);

INVx6_ASAP7_75t_SL g272 ( 
.A(n_236),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_272),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_159),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_211),
.B(n_229),
.C(n_218),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_161),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_223),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_201),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_224),
.B(n_171),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_287),
.B(n_237),
.Y(n_296)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_211),
.B(n_204),
.C(n_205),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_225),
.A2(n_185),
.B1(n_194),
.B2(n_211),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_231),
.A2(n_232),
.B(n_244),
.Y(n_282)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_204),
.B(n_216),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_285),
.C(n_251),
.Y(n_315)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_236),
.Y(n_284)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_215),
.B(n_201),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_246),
.B(n_214),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_237),
.B(n_241),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_250),
.A2(n_231),
.B1(n_256),
.B2(n_244),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_288),
.A2(n_303),
.B1(n_310),
.B2(n_264),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_291),
.Y(n_345)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_215),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_296),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_267),
.A2(n_233),
.B1(n_217),
.B2(n_228),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_294),
.A2(n_297),
.B(n_269),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_SL g297 ( 
.A(n_277),
.B(n_207),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_256),
.A2(n_233),
.B1(n_230),
.B2(n_241),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_299),
.A2(n_304),
.B1(n_306),
.B2(n_318),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_203),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_275),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_301),
.A2(n_277),
.B(n_287),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_240),
.B1(n_217),
.B2(n_228),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_271),
.A2(n_259),
.B1(n_261),
.B2(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_260),
.A2(n_253),
.B1(n_276),
.B2(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_265),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_282),
.A2(n_260),
.B1(n_265),
.B2(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_262),
.Y(n_321)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_321),
.Y(n_341)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_323),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_280),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_324),
.B(n_325),
.C(n_331),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_292),
.B(n_248),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_327),
.B(n_352),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_281),
.Y(n_330)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_330),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_283),
.C(n_249),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_283),
.C(n_286),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_350),
.C(n_319),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_317),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_333),
.B(n_340),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_291),
.B1(n_313),
.B2(n_302),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_247),
.Y(n_336)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_348),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_268),
.Y(n_338)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

AO22x1_ASAP7_75t_L g376 ( 
.A1(n_339),
.A2(n_317),
.B1(n_298),
.B2(n_323),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_300),
.A2(n_278),
.B(n_252),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_296),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_343),
.B(n_302),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_306),
.A2(n_291),
.B1(n_318),
.B2(n_299),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_346),
.A2(n_349),
.B1(n_303),
.B2(n_301),
.Y(n_360)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_312),
.Y(n_347)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_347),
.Y(n_365)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_295),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_272),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_255),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_289),
.B(n_255),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_309),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_290),
.B(n_284),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_311),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_353),
.B(n_358),
.Y(n_380)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_345),
.A2(n_316),
.B1(n_301),
.B2(n_293),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_359),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_322),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_361),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_342),
.A2(n_301),
.B1(n_294),
.B2(n_319),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_332),
.B(n_331),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_376),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_320),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_374),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_305),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_368),
.Y(n_392)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_371),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_336),
.B(n_314),
.Y(n_372)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_328),
.C(n_326),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_301),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_346),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_330),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_397),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_367),
.B(n_328),
.C(n_342),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_383),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_371),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_373),
.C(n_366),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_326),
.C(n_338),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_374),
.B(n_339),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_389),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_345),
.C(n_340),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_391),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_362),
.B(n_330),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_337),
.C(n_351),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_SL g403 ( 
.A(n_396),
.B(n_395),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_341),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_380),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_389),
.Y(n_418)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_393),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_400),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_390),
.A2(n_369),
.B(n_356),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_381),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_402),
.B(n_409),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_395),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_388),
.A2(n_361),
.B1(n_378),
.B2(n_386),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_406),
.A2(n_412),
.B1(n_396),
.B2(n_365),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_392),
.A2(n_370),
.B1(n_354),
.B2(n_364),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_407),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_397),
.A2(n_364),
.B1(n_356),
.B2(n_369),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_394),
.A2(n_377),
.B(n_376),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_413),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_379),
.A2(n_377),
.B1(n_376),
.B2(n_365),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_382),
.A2(n_341),
.B(n_348),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_416),
.B(n_404),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_398),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_419),
.Y(n_430)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_418),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_384),
.C(n_385),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_408),
.B(n_387),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_408),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_422),
.A2(n_400),
.B1(n_412),
.B2(n_406),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_401),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_425),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_335),
.C(n_347),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_428),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_425),
.C(n_411),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_434),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_422),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_414),
.C(n_344),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_335),
.B1(n_344),
.B2(n_314),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_435),
.B(n_436),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_298),
.Y(n_436)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_416),
.C(n_418),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_441),
.B(n_442),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_430),
.B(n_426),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_437),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_445),
.B(n_446),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_441),
.A2(n_431),
.B(n_432),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_443),
.A2(n_433),
.B(n_434),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_447),
.B(n_438),
.Y(n_449)
);

AOI32xp33_ASAP7_75t_L g451 ( 
.A1(n_449),
.A2(n_450),
.A3(n_439),
.B1(n_420),
.B2(n_258),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_448),
.B(n_444),
.C(n_440),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_284),
.C(n_258),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_258),
.Y(n_453)
);


endmodule