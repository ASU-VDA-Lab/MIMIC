module fake_jpeg_13468_n_300 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_247;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_273;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx9p33_ASAP7_75t_R g42 ( 
.A(n_41),
.Y(n_42)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_43),
.B(n_14),
.Y(n_71)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_59),
.Y(n_70)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_1),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx2_ASAP7_75t_SL g83 ( 
.A(n_62),
.Y(n_83)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_63),
.Y(n_107)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_19),
.B(n_1),
.CON(n_67),
.SN(n_67)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_3),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_78),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_35),
.B1(n_33),
.B2(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_73),
.A2(n_77),
.B1(n_80),
.B2(n_84),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_40),
.B1(n_39),
.B2(n_25),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_75),
.A2(n_79),
.B1(n_7),
.B2(n_8),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_35),
.B1(n_33),
.B2(n_32),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_40),
.B1(n_27),
.B2(n_25),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_32),
.B1(n_22),
.B2(n_27),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_22),
.B1(n_27),
.B2(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_101),
.Y(n_128)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_38),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_106),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_17),
.B1(n_36),
.B2(n_19),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_37),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_37),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_5),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_42),
.A2(n_20),
.B1(n_17),
.B2(n_28),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_80),
.B1(n_82),
.B2(n_74),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_36),
.B1(n_17),
.B2(n_20),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_112),
.A2(n_133),
.B1(n_110),
.B2(n_104),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_145),
.B1(n_111),
.B2(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_120),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_3),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_128),
.B(n_136),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_70),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_3),
.C(n_5),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_127),
.C(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_89),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_135),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_7),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_69),
.B1(n_74),
.B2(n_88),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

AOI32xp33_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_73),
.A3(n_77),
.B1(n_89),
.B2(n_84),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_144),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_75),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_15),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_9),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_102),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_15),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_141),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_83),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_16),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_76),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_144),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_85),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_69),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_139),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_147),
.A2(n_151),
.B1(n_160),
.B2(n_157),
.Y(n_195)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_154),
.B1(n_137),
.B2(n_162),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_104),
.B1(n_102),
.B2(n_105),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_167),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_134),
.B1(n_127),
.B2(n_133),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_170),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_117),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_119),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_134),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_113),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_163),
.C(n_153),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_115),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_121),
.A2(n_114),
.B(n_142),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_153),
.B(n_155),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_124),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_123),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_159),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_179),
.A2(n_146),
.B(n_137),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_160),
.A2(n_129),
.B1(n_131),
.B2(n_118),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_208),
.B1(n_186),
.B2(n_204),
.Y(n_213)
);

AO22x1_ASAP7_75t_SL g182 ( 
.A1(n_179),
.A2(n_146),
.B1(n_131),
.B2(n_139),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_188),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_187),
.B(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_202),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_191),
.B(n_193),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_158),
.C(n_148),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_201),
.C(n_192),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_151),
.A2(n_147),
.B1(n_154),
.B2(n_172),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_176),
.B1(n_173),
.B2(n_171),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_171),
.A2(n_156),
.B(n_152),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_204),
.B(n_209),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_177),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_149),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_205),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_208),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_230),
.C(n_191),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_229),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_228),
.B(n_217),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_209),
.B(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_180),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_207),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_233),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_226),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_182),
.B1(n_193),
.B2(n_181),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_238),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_219),
.B1(n_222),
.B2(n_227),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_221),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_239),
.A2(n_251),
.B(n_252),
.Y(n_265)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_215),
.C(n_212),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_182),
.B1(n_201),
.B2(n_200),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_210),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_218),
.C(n_232),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_250),
.C(n_228),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_224),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_216),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_249),
.B(n_252),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_222),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_248),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_214),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_231),
.B(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_221),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_256),
.C(n_257),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_244),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_212),
.C(n_211),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g258 ( 
.A(n_235),
.B(n_211),
.C(n_220),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_243),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_242),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_250),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_210),
.B(n_220),
.C(n_235),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_238),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_239),
.B(n_248),
.Y(n_267)
);

BUFx12f_ASAP7_75t_SL g266 ( 
.A(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_273),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_268),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_272),
.Y(n_283)
);

NOR4xp25_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_234),
.C(n_236),
.D(n_242),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_275),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_257),
.C(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_280),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_261),
.B1(n_264),
.B2(n_237),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_262),
.B1(n_237),
.B2(n_263),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_237),
.B1(n_242),
.B2(n_255),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_278),
.A2(n_234),
.B(n_270),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_287),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_254),
.Y(n_285)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_285),
.B(n_286),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_247),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_255),
.C(n_247),
.Y(n_288)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_288),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_289),
.A2(n_282),
.B1(n_279),
.B2(n_277),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_288),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_290),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_295),
.B(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_296),
.B(n_290),
.Y(n_297)
);

OAI21xp33_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_292),
.B(n_251),
.Y(n_298)
);

OAI211xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_258),
.B(n_280),
.C(n_240),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_287),
.Y(n_300)
);


endmodule