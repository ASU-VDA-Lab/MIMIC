module real_jpeg_31076_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_626, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_626;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_602;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_0),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_0),
.Y(n_271)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_0),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_1),
.B(n_181),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_1),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_2),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_2),
.B(n_152),
.Y(n_258)
);

NAND2x1_ASAP7_75t_L g277 ( 
.A(n_2),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_2),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_2),
.B(n_359),
.Y(n_358)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_2),
.B(n_160),
.C(n_465),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_2),
.B(n_470),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_2),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_2),
.B(n_465),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_SL g548 ( 
.A(n_2),
.B(n_160),
.C(n_465),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_3),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_4),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_5),
.Y(n_126)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_5),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_5),
.Y(n_467)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_5),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_6),
.B(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_6),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_6),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g337 ( 
.A(n_6),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_6),
.B(n_427),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_6),
.B(n_220),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_6),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_6),
.B(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_7),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_7),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_7),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_7),
.B(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_7),
.B(n_499),
.Y(n_498)
);

BUFx2_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_8),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_8),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_8),
.B(n_100),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_8),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_8),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_8),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_8),
.B(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_9),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_9),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_10),
.Y(n_342)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_11),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_12),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_12),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_13),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_13),
.B(n_220),
.Y(n_219)
);

AOI22x1_ASAP7_75t_L g343 ( 
.A1(n_13),
.A2(n_14),
.B1(n_344),
.B2(n_347),
.Y(n_343)
);

NAND2x1_ASAP7_75t_L g267 ( 
.A(n_14),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_14),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_14),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_14),
.B(n_424),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_14),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_14),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_14),
.B(n_526),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_15),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_16),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_16),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_16),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_16),
.B(n_124),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g150 ( 
.A(n_16),
.B(n_107),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_16),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_17),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_17),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_17),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_SL g332 ( 
.A(n_17),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_17),
.B(n_385),
.Y(n_384)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_182),
.A3(n_603),
.B1(n_616),
.B2(n_617),
.C(n_622),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_179),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI332xp33_ASAP7_75t_L g622 ( 
.A1(n_21),
.A2(n_179),
.A3(n_603),
.B1(n_618),
.B2(n_619),
.B3(n_623),
.C1(n_624),
.C2(n_626),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_111),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_86),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_23),
.B(n_86),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_52),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_24),
.B(n_52),
.C(n_86),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.C(n_47),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_26),
.A2(n_27),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_26),
.B(n_123),
.C(n_127),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_26),
.A2(n_27),
.B1(n_306),
.B2(n_419),
.Y(n_418)
);

CKINVDCx11_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_27),
.B(n_306),
.C(n_309),
.Y(n_305)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_29),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_29),
.Y(n_520)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_30),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_30),
.A2(n_174),
.B1(n_609),
.B2(n_610),
.Y(n_608)
);

NAND2x1_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_36),
.Y(n_163)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_36),
.Y(n_361)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_37),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_38),
.A2(n_59),
.B1(n_68),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_38),
.A2(n_59),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_38),
.A2(n_59),
.B1(n_315),
.B2(n_320),
.Y(n_314)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2x1_ASAP7_75t_R g103 ( 
.A(n_43),
.B(n_104),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_43),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_43),
.B(n_228),
.Y(n_236)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_50),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_51),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_51),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_74),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_54),
.B(n_74),
.C(n_613),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_58),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.C(n_68),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_59),
.B(n_315),
.C(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_62),
.B(n_123),
.C(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_63),
.B(n_131),
.Y(n_208)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_67),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_67),
.Y(n_434)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_69),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_68),
.A2(n_69),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_69),
.B(n_80),
.C(n_84),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_70),
.B(n_267),
.C(n_269),
.Y(n_266)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_71),
.Y(n_454)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_72),
.Y(n_359)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_73),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_73),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_84),
.B2(n_85),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

XOR2x2_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_75),
.B(n_142),
.C(n_144),
.Y(n_175)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_79),
.B(n_214),
.C(n_218),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_79),
.A2(n_80),
.B1(n_149),
.B2(n_150),
.Y(n_610)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_80),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_83),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.C(n_108),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2x1_ASAP7_75t_L g177 ( 
.A(n_88),
.B(n_178),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_91),
.B(n_109),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.C(n_103),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_92),
.A2(n_93),
.B1(n_99),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_94),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_94),
.B(n_398),
.Y(n_397)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_99),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_99),
.B(n_160),
.C(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_100),
.Y(n_308)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2x1_ASAP7_75t_L g166 ( 
.A(n_103),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_111),
.B(n_621),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_169),
.C(n_177),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_112),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_113),
.A2(n_170),
.B(n_177),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_146),
.C(n_165),
.Y(n_113)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_129),
.C(n_136),
.Y(n_114)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_115),
.Y(n_287)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_123),
.B1(n_127),
.B2(n_128),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_118),
.Y(n_127)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_120),
.Y(n_268)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_123),
.B(n_269),
.Y(n_382)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_128),
.B(n_208),
.Y(n_207)
);

XOR2x2_ASAP7_75t_L g461 ( 
.A(n_128),
.B(n_269),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_129),
.A2(n_130),
.B1(n_136),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_134),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_136),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_137)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_138),
.A2(n_144),
.B1(n_257),
.B2(n_258),
.Y(n_355)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_140),
.Y(n_429)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_141),
.Y(n_312)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_144),
.B(n_252),
.C(n_256),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_144),
.A2(n_252),
.B(n_256),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_146),
.A2(n_147),
.B1(n_166),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_155),
.B(n_164),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_151),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_149),
.B(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_149),
.A2(n_150),
.B1(n_227),
.B2(n_236),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_150),
.A2(n_227),
.B(n_230),
.C(n_235),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_162),
.Y(n_155)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_156),
.A2(n_210),
.B1(n_357),
.B2(n_358),
.Y(n_407)
);

OR2x2_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_157),
.Y(n_471)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_158),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_162),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_160),
.A2(n_231),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

XNOR2x2_ASAP7_75t_L g484 ( 
.A(n_160),
.B(n_485),
.Y(n_484)
);

INVx8_ASAP7_75t_L g399 ( 
.A(n_161),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_168),
.A2(n_245),
.B(n_248),
.Y(n_244)
);

OAI211xp5_ASAP7_75t_L g248 ( 
.A1(n_168),
.A2(n_231),
.B(n_247),
.C(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_177),
.B1(n_189),
.B2(n_190),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.C(n_176),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_180),
.B(n_619),
.Y(n_618)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_182),
.Y(n_616)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_290),
.B(n_599),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_237),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_186),
.A2(n_601),
.B(n_602),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_194),
.Y(n_186)
);

NOR2xp67_ASAP7_75t_L g602 ( 
.A(n_187),
.B(n_194),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_191),
.B(n_192),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.C(n_203),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_201),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_223),
.C(n_226),
.Y(n_204)
);

XOR2x1_ASAP7_75t_SL g288 ( 
.A(n_205),
.B(n_289),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.C(n_212),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_207),
.B(n_213),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_209),
.B(n_573),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_210),
.B(n_357),
.C(n_360),
.Y(n_356)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_222),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_223),
.B(n_226),
.Y(n_289)
);

INVx5_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_247),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_231),
.B(n_301),
.Y(n_300)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_234),
.Y(n_323)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_234),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_L g601 ( 
.A(n_238),
.B(n_240),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_283),
.C(n_288),
.Y(n_240)
);

INVxp33_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_242),
.B(n_284),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_263),
.C(n_280),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_243),
.B(n_570),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.C(n_260),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_244),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_L g420 ( 
.A(n_246),
.B(n_301),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_250),
.B(n_261),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_257),
.B(n_259),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_252),
.B(n_256),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_264),
.B(n_281),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.C(n_277),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_266),
.B(n_368),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_270),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_271),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_273),
.A2(n_274),
.B1(n_277),
.B2(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_277),
.Y(n_369)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_279),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g580 ( 
.A(n_288),
.B(n_581),
.Y(n_580)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_590),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_440),
.C(n_565),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_412),
.Y(n_293)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_294),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_374),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_295),
.B(n_374),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_350),
.B2(n_373),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_296),
.B(n_584),
.C(n_585),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_325),
.C(n_329),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_298),
.B(n_376),
.Y(n_375)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_313),
.B(n_324),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_305),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_300),
.B(n_305),
.Y(n_437)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_302),
.B(n_510),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_302),
.B(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_306),
.Y(n_419)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_SL g417 ( 
.A(n_309),
.B(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_312),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_313),
.B(n_437),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_321),
.Y(n_313)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_315),
.Y(n_320)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx4f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_329),
.Y(n_376)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_343),
.B2(n_349),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_337),
.Y(n_331)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_332),
.Y(n_365)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_343),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_365),
.C(n_366),
.Y(n_364)
);

INVx3_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_345),
.B(n_480),
.Y(n_479)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_397),
.B(n_400),
.Y(n_396)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_370),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_351),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_363),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g575 ( 
.A(n_352),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_356),
.C(n_362),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_353),
.B(n_356),
.Y(n_411)
);

XNOR2x1_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_360),
.Y(n_406)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

XNOR2x1_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_364),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_367),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_370),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.C(n_408),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_375),
.B(n_439),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_409),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_396),
.C(n_404),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_415),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.C(n_389),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_381),
.A2(n_382),
.B1(n_550),
.B2(n_551),
.Y(n_549)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_383),
.A2(n_384),
.B1(n_390),
.B2(n_391),
.Y(n_551)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_388),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_405),
.Y(n_415)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_438),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_413),
.B(n_438),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.C(n_435),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_414),
.B(n_558),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_416),
.A2(n_436),
.B1(n_559),
.B2(n_560),
.Y(n_558)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_416),
.Y(n_560)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_420),
.C(n_421),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_417),
.B(n_542),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_420),
.A2(n_421),
.B1(n_543),
.B2(n_544),
.Y(n_542)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_420),
.Y(n_544)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_421),
.Y(n_543)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_426),
.C(n_430),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_422),
.A2(n_423),
.B1(n_430),
.B2(n_431),
.Y(n_449)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_449),
.Y(n_448)
);

INVx3_ASAP7_75t_SL g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_436),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_555),
.B(n_564),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_443),
.A2(n_538),
.B(n_554),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_486),
.B(n_537),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_472),
.C(n_473),
.Y(n_444)
);

AOI21xp33_ASAP7_75t_SL g537 ( 
.A1(n_445),
.A2(n_472),
.B(n_473),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_459),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_447),
.Y(n_446)
);

NAND2xp33_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_460),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_450),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_448),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_450),
.B(n_459),
.C(n_553),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_455),
.C(n_456),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_451),
.A2(n_452),
.B1(n_455),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_455),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_475),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_457),
.B(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_461),
.B(n_468),
.C(n_548),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_R g563 ( 
.A(n_461),
.B(n_468),
.C(n_548),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_464),
.B1(n_468),
.B2(n_469),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.C(n_484),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_474),
.B(n_501),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_477),
.A2(n_478),
.B1(n_484),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_479),
.A2(n_481),
.B1(n_482),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_479),
.Y(n_491)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_484),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_503),
.B(n_536),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_500),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_488),
.B(n_500),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_492),
.C(n_498),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_489),
.A2(n_490),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_493),
.B(n_498),
.Y(n_532)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_530),
.B(n_535),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_515),
.B(n_529),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_509),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_521),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_521),
.Y(n_529)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_524),
.B1(n_525),
.B2(n_528),
.Y(n_521)
);

CKINVDCx14_ASAP7_75t_R g528 ( 
.A(n_522),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_528),
.Y(n_534)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_531),
.B(n_534),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_534),
.Y(n_535)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_532),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_552),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_552),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_540),
.A2(n_541),
.B1(n_545),
.B2(n_546),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_540),
.B(n_562),
.C(n_563),
.Y(n_561)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_549),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_549),
.Y(n_562)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_557),
.B(n_561),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_557),
.B(n_561),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_565),
.A2(n_591),
.B(n_595),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_566),
.A2(n_579),
.B1(n_582),
.B2(n_586),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

NOR2xp67_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_580),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_567),
.B(n_580),
.Y(n_598)
);

OAI22x1_ASAP7_75t_L g567 ( 
.A1(n_568),
.A2(n_571),
.B1(n_574),
.B2(n_578),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_569),
.B(n_572),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_574),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_572),
.Y(n_578)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_574),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_576),
.C(n_577),
.Y(n_574)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_583),
.B(n_587),
.Y(n_597)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_589),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_592),
.A2(n_593),
.B(n_594),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_596),
.A2(n_597),
.B(n_598),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_603),
.B(n_618),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_603),
.Y(n_623)
);

AO21x1_ASAP7_75t_L g603 ( 
.A1(n_604),
.A2(n_614),
.B(n_615),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_614),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_612),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_606),
.A2(n_607),
.B1(n_608),
.B2(n_611),
.Y(n_605)
);

CKINVDCx11_ASAP7_75t_R g606 ( 
.A(n_607),
.Y(n_606)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_608),
.Y(n_611)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);


endmodule