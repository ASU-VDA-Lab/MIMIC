module fake_ibex_484_n_1615 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_9, n_293, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_239, n_94, n_134, n_88, n_142, n_226, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_105, n_187, n_1, n_154, n_182, n_196, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_143, n_106, n_8, n_224, n_183, n_67, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_57, n_301, n_296, n_120, n_168, n_155, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_211, n_218, n_132, n_277, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_55, n_291, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_119, n_72, n_195, n_212, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1615);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_9;
input n_293;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_211;
input n_218;
input n_132;
input n_277;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_55;
input n_291;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_119;
input n_72;
input n_195;
input n_212;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1615;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1614;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1558;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_422;
wire n_1609;
wire n_324;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1610;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_1591;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_1577;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_1568;
wire n_325;
wire n_1477;
wire n_1184;
wire n_1364;
wire n_1540;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_1115;
wire n_998;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_650;
wire n_409;
wire n_1575;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_633;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_1607;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_1604;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1415;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_416;
wire n_1472;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_87),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_47),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_107),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_81),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_56),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_271),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_281),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_136),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_25),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_149),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_161),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_236),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_214),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_230),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_217),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_309),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_300),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_78),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_10),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_248),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_249),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_196),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_84),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_264),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_176),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_258),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_160),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_246),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_89),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_134),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_18),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_103),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_239),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_60),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_251),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_245),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_99),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_267),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_220),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_146),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_86),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_6),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_55),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_155),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_223),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_8),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_170),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_14),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_168),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_180),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_216),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_193),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_234),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_273),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_247),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_122),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_206),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_201),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_12),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_106),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_227),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_280),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_229),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_265),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_294),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_148),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_138),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_182),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_296),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_211),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_76),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_241),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_144),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_169),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_108),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_290),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_179),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_183),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_224),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_63),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_215),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_151),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_304),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_291),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_175),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_293),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_226),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_261),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_242),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_213),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_9),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_112),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_145),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_270),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_126),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_98),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_63),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_67),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_235),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_56),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_174),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_96),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_87),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_43),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_228),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_233),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_34),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_11),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_252),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_181),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_6),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_61),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_282),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_27),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_250),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_255),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_28),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_210),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_292),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_65),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_272),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_307),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_269),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_238),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_263),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_189),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_59),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_266),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_101),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_256),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_163),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_133),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_287),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_244),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_221),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_297),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_208),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_310),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_302),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_7),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_72),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_16),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_89),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_132),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_11),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_232),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_284),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_31),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_166),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_113),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_64),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_283),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_42),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_204),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_259),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_81),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_57),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_231),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_14),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_157),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_167),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_79),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_171),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_152),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_159),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_121),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_212),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_184),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_219),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_37),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_253),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_202),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_82),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_301),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_94),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_195),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_30),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_240),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_118),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_276),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_22),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_222),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_218),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_42),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_62),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_21),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_286),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_44),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_83),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_298),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_299),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_140),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_116),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_205),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_274),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_279),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_243),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_203),
.Y(n_513)
);

CKINVDCx14_ASAP7_75t_R g514 ( 
.A(n_295),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_268),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_177),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_285),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_190),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_275),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_254),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_225),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_40),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_117),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_8),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_72),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_93),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_100),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_129),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_142),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_262),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_260),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_303),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_55),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_288),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_154),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_153),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_58),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_200),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_209),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_191),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_257),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_412),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_432),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_313),
.B(n_0),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_327),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_328),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_352),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_331),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_463),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_423),
.B(n_0),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_392),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_369),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_539),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g554 ( 
.A(n_356),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_350),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_439),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_372),
.Y(n_557)
);

NOR2xp67_ASAP7_75t_L g558 ( 
.A(n_352),
.B(n_1),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_345),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_477),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_446),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_516),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_395),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_315),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_373),
.B(n_1),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_379),
.B(n_2),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_395),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_442),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_315),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_442),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_312),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_456),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_364),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_505),
.B(n_2),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_456),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_530),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_316),
.Y(n_577)
);

NOR2xp67_ASAP7_75t_L g578 ( 
.A(n_526),
.B(n_3),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_397),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_347),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_332),
.Y(n_581)
);

INVxp33_ASAP7_75t_SL g582 ( 
.A(n_343),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_386),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_435),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_415),
.B(n_3),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_397),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_311),
.B(n_4),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_435),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_499),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_427),
.B(n_4),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_317),
.B(n_5),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_319),
.B(n_5),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_455),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_483),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_458),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_314),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_483),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_460),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_323),
.Y(n_599)
);

INVxp33_ASAP7_75t_SL g600 ( 
.A(n_349),
.Y(n_600)
);

INVxp33_ASAP7_75t_SL g601 ( 
.A(n_358),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_468),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_362),
.Y(n_603)
);

NOR2xp67_ASAP7_75t_L g604 ( 
.A(n_471),
.B(n_7),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_472),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_485),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_362),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_492),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_361),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_514),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_501),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_499),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_514),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_323),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_314),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_314),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_467),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_363),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_374),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_406),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_364),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_467),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_323),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_573),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_580),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_545),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_573),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_596),
.B(n_419),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_559),
.A2(n_452),
.B(n_380),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_583),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_618),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_593),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_548),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_621),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_595),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_621),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_560),
.B(n_554),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_602),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_605),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_555),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_556),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_561),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_606),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_608),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_559),
.A2(n_452),
.B(n_380),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_611),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_563),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_596),
.B(n_461),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_567),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_568),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_570),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_547),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_547),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_562),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_572),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_575),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_596),
.B(n_615),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_585),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_599),
.B(n_357),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_564),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_547),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_579),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_616),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_586),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_617),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_622),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_546),
.B(n_419),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_594),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_587),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_591),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_598),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_544),
.B(n_419),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_592),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_565),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_551),
.B(n_553),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_557),
.B(n_434),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_571),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_552),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_597),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_566),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_574),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_558),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_564),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_550),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_603),
.B(n_461),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_582),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_578),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_542),
.B(n_357),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_577),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_590),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_569),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_604),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_581),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_607),
.B(n_497),
.Y(n_694)
);

OA21x2_ASAP7_75t_L g695 ( 
.A1(n_609),
.A2(n_507),
.B(n_497),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_619),
.B(n_419),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_600),
.A2(n_511),
.B(n_507),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_610),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_582),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_613),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_601),
.B(n_511),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_601),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_543),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_569),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_543),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_620),
.B(n_576),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_549),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_614),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_614),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_623),
.B(n_512),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_549),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_623),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_584),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_584),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_588),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_588),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_589),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_589),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_612),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_612),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_564),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_573),
.B(n_512),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_573),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_596),
.B(n_517),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_596),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_545),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_596),
.B(n_517),
.Y(n_727)
);

CKINVDCx16_ASAP7_75t_R g728 ( 
.A(n_552),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_573),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_545),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_618),
.Y(n_731)
);

BUFx8_ASAP7_75t_L g732 ( 
.A(n_585),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_596),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_545),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_580),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_573),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_573),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_573),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_545),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_596),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_573),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_545),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_580),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_596),
.B(n_540),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_571),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_573),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_580),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_564),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_580),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_571),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_573),
.Y(n_751)
);

NOR2x1_ASAP7_75t_L g752 ( 
.A(n_596),
.B(n_324),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_573),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_596),
.B(n_540),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_580),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_545),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_580),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_596),
.B(n_336),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_573),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_596),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_545),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_596),
.B(n_338),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_545),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_573),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_628),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_689),
.Y(n_766)
);

INVx6_ASAP7_75t_L g767 ( 
.A(n_678),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_629),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_741),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_741),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_657),
.B(n_333),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_631),
.B(n_339),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_645),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_703),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_697),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_689),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_628),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_684),
.B(n_318),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_653),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_741),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_710),
.B(n_413),
.C(n_411),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_731),
.Y(n_782)
);

AND2x6_ASAP7_75t_L g783 ( 
.A(n_659),
.B(n_443),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_686),
.A2(n_418),
.B1(n_422),
.B2(n_417),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_667),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_657),
.B(n_337),
.Y(n_786)
);

INVx8_ASAP7_75t_L g787 ( 
.A(n_678),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_L g788 ( 
.A1(n_699),
.A2(n_429),
.B1(n_444),
.B2(n_426),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_745),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_746),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_667),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_725),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_725),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_746),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_675),
.A2(n_466),
.B1(n_474),
.B2(n_457),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_745),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_684),
.A2(n_357),
.B1(n_355),
.B2(n_342),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_705),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_750),
.B(n_488),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_674),
.B(n_467),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_671),
.B(n_320),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_733),
.Y(n_802)
);

INVx5_ASAP7_75t_L g803 ( 
.A(n_759),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_733),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_740),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_678),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_702),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_740),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_677),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_750),
.Y(n_810)
);

AND2x6_ASAP7_75t_L g811 ( 
.A(n_752),
.B(n_443),
.Y(n_811)
);

INVx4_ASAP7_75t_SL g812 ( 
.A(n_672),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_663),
.B(n_321),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_760),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_760),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_732),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_663),
.B(n_329),
.Y(n_817)
);

AND2x2_ASAP7_75t_SL g818 ( 
.A(n_728),
.B(n_365),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_665),
.B(n_330),
.Y(n_819)
);

INVxp33_ASAP7_75t_L g820 ( 
.A(n_713),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_661),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_665),
.B(n_334),
.Y(n_822)
);

BUFx4f_ASAP7_75t_L g823 ( 
.A(n_675),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_764),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_732),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_688),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_764),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_680),
.B(n_335),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_666),
.B(n_340),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_701),
.B(n_658),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_674),
.B(n_341),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_698),
.B(n_453),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_637),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_701),
.B(n_322),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_685),
.B(n_325),
.Y(n_835)
);

OR2x2_ASAP7_75t_L g836 ( 
.A(n_693),
.B(n_346),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_674),
.B(n_344),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_708),
.B(n_366),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_685),
.B(n_326),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_681),
.B(n_669),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_678),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_764),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_672),
.A2(n_676),
.B1(n_710),
.B2(n_625),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_653),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_661),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_653),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_706),
.B(n_490),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_624),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_698),
.B(n_496),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_634),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_652),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_627),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_672),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_SL g854 ( 
.A(n_626),
.B(n_500),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_636),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_647),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_696),
.B(n_503),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_649),
.Y(n_858)
);

AND2x6_ASAP7_75t_L g859 ( 
.A(n_681),
.B(n_453),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_681),
.B(n_348),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_696),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_707),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_723),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_662),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_650),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_651),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_695),
.Y(n_867)
);

NAND3x1_ASAP7_75t_L g868 ( 
.A(n_714),
.B(n_378),
.C(n_370),
.Y(n_868)
);

AO22x1_ASAP7_75t_L g869 ( 
.A1(n_758),
.A2(n_387),
.B1(n_399),
.B2(n_382),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_711),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_695),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_729),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_694),
.B(n_368),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_736),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_630),
.B(n_504),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_737),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_655),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_738),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_751),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_669),
.B(n_351),
.Y(n_880)
);

BUFx8_ASAP7_75t_SL g881 ( 
.A(n_704),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_753),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_656),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_633),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_694),
.B(n_394),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_700),
.B(n_522),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_669),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_722),
.Y(n_888)
);

AND2x4_ASAP7_75t_SL g889 ( 
.A(n_709),
.B(n_720),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_722),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_632),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_635),
.B(n_353),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_638),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_639),
.B(n_354),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_690),
.B(n_692),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_640),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_643),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_644),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_763),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_646),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_670),
.B(n_410),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_641),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_735),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_670),
.A2(n_405),
.B1(n_414),
.B2(n_408),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_648),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_743),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_747),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_749),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_648),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_755),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_757),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_670),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_724),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_724),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_673),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_727),
.Y(n_916)
);

INVxp33_ASAP7_75t_L g917 ( 
.A(n_713),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_673),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_673),
.B(n_421),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_682),
.B(n_524),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_727),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_642),
.Y(n_922)
);

AND2x6_ASAP7_75t_L g923 ( 
.A(n_758),
.B(n_493),
.Y(n_923)
);

NAND3x1_ASAP7_75t_L g924 ( 
.A(n_715),
.B(n_424),
.C(n_416),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_676),
.B(n_525),
.Y(n_925)
);

OR2x6_ASAP7_75t_L g926 ( 
.A(n_720),
.B(n_431),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_654),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_687),
.B(n_527),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_762),
.B(n_359),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_720),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_762),
.B(n_360),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_726),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_744),
.B(n_371),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_744),
.B(n_375),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_754),
.B(n_376),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_754),
.B(n_377),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_730),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_717),
.B(n_381),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_664),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_668),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_679),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_L g942 ( 
.A(n_734),
.B(n_537),
.C(n_533),
.Y(n_942)
);

AND2x6_ASAP7_75t_L g943 ( 
.A(n_719),
.B(n_493),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_712),
.B(n_9),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_739),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_742),
.B(n_383),
.Y(n_946)
);

INVxp67_ASAP7_75t_SL g947 ( 
.A(n_660),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_756),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_761),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_716),
.B(n_384),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_718),
.Y(n_951)
);

BUFx10_ASAP7_75t_L g952 ( 
.A(n_683),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_691),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_748),
.Y(n_954)
);

BUFx4f_ASAP7_75t_L g955 ( 
.A(n_704),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_721),
.B(n_541),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_721),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_684),
.B(n_385),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_657),
.B(n_438),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_741),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_689),
.Y(n_961)
);

CKINVDCx8_ASAP7_75t_R g962 ( 
.A(n_728),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_741),
.Y(n_963)
);

AND2x6_ASAP7_75t_L g964 ( 
.A(n_659),
.B(n_450),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_628),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_631),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_684),
.B(n_388),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_741),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_703),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_628),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_628),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_741),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_684),
.B(n_389),
.Y(n_973)
);

AND2x6_ASAP7_75t_L g974 ( 
.A(n_659),
.B(n_538),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_684),
.B(n_390),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_657),
.B(n_459),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_629),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_689),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_741),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_628),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_663),
.B(n_393),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_741),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_888),
.B(n_396),
.Y(n_983)
);

AND2x6_ASAP7_75t_L g984 ( 
.A(n_775),
.B(n_469),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_905),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_830),
.A2(n_888),
.B(n_914),
.C(n_913),
.Y(n_986)
);

AOI21x1_ASAP7_75t_L g987 ( 
.A1(n_768),
.A2(n_536),
.B(n_478),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_905),
.B(n_398),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_SL g989 ( 
.A1(n_776),
.A2(n_401),
.B1(n_402),
.B2(n_400),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_789),
.B(n_535),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_905),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_978),
.B(n_403),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_809),
.B(n_404),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_810),
.B(n_10),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_909),
.A2(n_470),
.B1(n_484),
.B2(n_479),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_909),
.Y(n_996)
);

AND2x6_ASAP7_75t_SL g997 ( 
.A(n_881),
.B(n_486),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_890),
.B(n_407),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_823),
.A2(n_495),
.B1(n_506),
.B2(n_494),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_796),
.A2(n_518),
.B1(n_529),
.B2(n_515),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_768),
.A2(n_532),
.B(n_420),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_961),
.B(n_12),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_L g1003 ( 
.A(n_775),
.B(n_105),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_823),
.B(n_409),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_890),
.B(n_425),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_890),
.B(n_428),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_766),
.B(n_534),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_914),
.A2(n_367),
.B(n_487),
.C(n_391),
.Y(n_1008)
);

AND2x6_ASAP7_75t_SL g1009 ( 
.A(n_954),
.B(n_13),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_787),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_921),
.A2(n_345),
.B1(n_433),
.B2(n_430),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_952),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_834),
.B(n_436),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_787),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_858),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_816),
.B(n_367),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_833),
.B(n_437),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_835),
.B(n_440),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_891),
.A2(n_531),
.B1(n_445),
.B2(n_447),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_853),
.B(n_441),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_853),
.B(n_812),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_839),
.B(n_448),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_893),
.A2(n_451),
.B1(n_454),
.B2(n_449),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_820),
.B(n_462),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_812),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_917),
.B(n_464),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_799),
.A2(n_465),
.B1(n_475),
.B2(n_473),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_858),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_773),
.A2(n_480),
.B(n_476),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_883),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_778),
.B(n_481),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_873),
.B(n_482),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_847),
.B(n_491),
.Y(n_1033)
);

BUFx5_ASAP7_75t_L g1034 ( 
.A(n_977),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_885),
.B(n_498),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_958),
.B(n_502),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_882),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_967),
.B(n_508),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_972),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_883),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_973),
.B(n_509),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_SL g1042 ( 
.A1(n_901),
.A2(n_510),
.B(n_519),
.C(n_513),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_916),
.A2(n_521),
.B(n_520),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_877),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_782),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_966),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_SL g1047 ( 
.A1(n_818),
.A2(n_528),
.B1(n_523),
.B2(n_391),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_975),
.B(n_345),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_962),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_964),
.A2(n_345),
.B1(n_391),
.B2(n_367),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_SL g1051 ( 
.A(n_952),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_877),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_900),
.B(n_903),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_897),
.B(n_345),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_898),
.A2(n_367),
.B(n_487),
.C(n_391),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_806),
.B(n_13),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_906),
.A2(n_489),
.B1(n_487),
.B2(n_17),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_907),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_883),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_840),
.A2(n_489),
.B(n_487),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_767),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_882),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_807),
.B(n_15),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_972),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_841),
.B(n_15),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_908),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_921),
.A2(n_345),
.B1(n_489),
.B2(n_18),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_849),
.B(n_345),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_856),
.A2(n_489),
.B(n_110),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_886),
.B(n_16),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_849),
.B(n_17),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_910),
.B(n_19),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_911),
.B(n_19),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_912),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_875),
.B(n_20),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_921),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_767),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_843),
.B(n_23),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_SL g1079 ( 
.A1(n_854),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_869),
.B(n_26),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_869),
.B(n_27),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_865),
.B(n_28),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_785),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_886),
.B(n_29),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_866),
.B(n_29),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_867),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1086)
);

O2A1O1Ixp5_ASAP7_75t_L g1087 ( 
.A1(n_867),
.A2(n_871),
.B(n_931),
.C(n_800),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_783),
.B(n_33),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_918),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_959),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_981),
.B(n_35),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_791),
.Y(n_1092)
);

NAND2x1_ASAP7_75t_L g1093 ( 
.A(n_779),
.B(n_109),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_783),
.B(n_36),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_826),
.B(n_36),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_971),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_871),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_813),
.B(n_38),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_959),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1099)
);

OR2x6_ASAP7_75t_L g1100 ( 
.A(n_825),
.B(n_41),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_971),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_783),
.B(n_43),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_864),
.B(n_44),
.Y(n_1103)
);

AND3x1_ASAP7_75t_L g1104 ( 
.A(n_957),
.B(n_45),
.C(n_46),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_976),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_783),
.B(n_797),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_772),
.B(n_48),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_887),
.Y(n_1108)
);

O2A1O1Ixp5_ASAP7_75t_L g1109 ( 
.A1(n_831),
.A2(n_114),
.B(n_115),
.C(n_111),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_980),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_L g1111 ( 
.A(n_832),
.B(n_119),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_925),
.B(n_48),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_915),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_980),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_976),
.B(n_49),
.Y(n_1115)
);

AND2x6_ASAP7_75t_SL g1116 ( 
.A(n_772),
.B(n_49),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_817),
.B(n_50),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_915),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_902),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_SL g1120 ( 
.A(n_884),
.B(n_50),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_L g1121 ( 
.A(n_781),
.B(n_51),
.C(n_52),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_972),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_819),
.B(n_822),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_857),
.B(n_51),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_771),
.B(n_52),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_771),
.B(n_53),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_786),
.B(n_53),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_930),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_930),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_765),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_777),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_964),
.A2(n_58),
.B1(n_54),
.B2(n_57),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_964),
.A2(n_61),
.B1(n_54),
.B2(n_59),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_922),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_965),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_784),
.B(n_788),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_964),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_855),
.Y(n_1138)
);

O2A1O1Ixp5_ASAP7_75t_L g1139 ( 
.A1(n_837),
.A2(n_207),
.B(n_308),
.C(n_306),
.Y(n_1139)
);

NOR3xp33_ASAP7_75t_SL g1140 ( 
.A(n_948),
.B(n_66),
.C(n_67),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_786),
.B(n_937),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_929),
.B(n_919),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_828),
.B(n_895),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_857),
.B(n_66),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_895),
.B(n_68),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_836),
.B(n_68),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_892),
.B(n_69),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_974),
.B(n_69),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_974),
.B(n_70),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_970),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_974),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_920),
.B(n_71),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_974),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_945),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_896),
.Y(n_1155)
);

OAI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_949),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_940),
.B(n_77),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_923),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_861),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_930),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_851),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_795),
.B(n_80),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_940),
.B(n_82),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_932),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_899),
.B(n_83),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_801),
.B(n_84),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_894),
.B(n_832),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1015),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1014),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1014),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1039),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1134),
.B(n_798),
.C(n_774),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1010),
.B(n_927),
.Y(n_1173)
);

INVxp67_ASAP7_75t_SL g1174 ( 
.A(n_1014),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1164),
.B(n_957),
.Y(n_1175)
);

NOR3xp33_ASAP7_75t_SL g1176 ( 
.A(n_1049),
.B(n_870),
.C(n_862),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1012),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1058),
.Y(n_1178)
);

AO22x1_ASAP7_75t_L g1179 ( 
.A1(n_984),
.A2(n_832),
.B1(n_945),
.B2(n_943),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1025),
.B(n_945),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_986),
.B(n_928),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1028),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1066),
.B(n_838),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1025),
.B(n_852),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1039),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1037),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1046),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_1119),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1044),
.B(n_838),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_989),
.B(n_1045),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1052),
.B(n_904),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1016),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1155),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1016),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1141),
.A2(n_969),
.B1(n_956),
.B2(n_951),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_994),
.B(n_953),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1039),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1083),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1143),
.B(n_939),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1136),
.B(n_947),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1107),
.B(n_926),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1092),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1130),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1146),
.B(n_941),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1154),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1100),
.B(n_993),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1016),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1131),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1112),
.B(n_934),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1100),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_1100),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1135),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1154),
.B(n_852),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1056),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1033),
.B(n_889),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1047),
.A2(n_926),
.B1(n_944),
.B2(n_950),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1150),
.Y(n_1217)
);

BUFx4f_ASAP7_75t_L g1218 ( 
.A(n_1056),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_SL g1219 ( 
.A(n_1051),
.B(n_955),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_985),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1065),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1065),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1051),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1027),
.B(n_1120),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1021),
.B(n_1002),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_997),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1162),
.A2(n_924),
.B1(n_868),
.B2(n_955),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1017),
.B(n_946),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1116),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1053),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1070),
.A2(n_938),
.B1(n_942),
.B2(n_943),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1072),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1101),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_992),
.B(n_874),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1075),
.B(n_832),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1073),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1082),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1064),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1085),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1064),
.Y(n_1240)
);

NOR2x1_ASAP7_75t_L g1241 ( 
.A(n_1121),
.B(n_860),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1161),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1063),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1125),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1037),
.B(n_829),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1024),
.B(n_935),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1126),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1009),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1026),
.B(n_792),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_984),
.Y(n_1250)
);

NOR3xp33_ASAP7_75t_SL g1251 ( 
.A(n_1156),
.B(n_1071),
.C(n_1090),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1007),
.B(n_1095),
.Y(n_1252)
);

AND3x1_ASAP7_75t_SL g1253 ( 
.A(n_1104),
.B(n_845),
.C(n_821),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1165),
.B(n_880),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1062),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1127),
.B(n_811),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1101),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1159),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_991),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1145),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1064),
.Y(n_1261)
);

INVxp67_ASAP7_75t_SL g1262 ( 
.A(n_1034),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1000),
.B(n_811),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1096),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1122),
.Y(n_1265)
);

AOI211xp5_ASAP7_75t_L g1266 ( 
.A1(n_1084),
.A2(n_936),
.B(n_933),
.C(n_802),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1062),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1103),
.B(n_793),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1078),
.A2(n_943),
.B1(n_923),
.B2(n_811),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1054),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1128),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1157),
.B(n_804),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1142),
.A2(n_808),
.B(n_814),
.C(n_805),
.Y(n_1273)
);

AND2x6_ASAP7_75t_L g1274 ( 
.A(n_996),
.B(n_815),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1110),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_1124),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1122),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1163),
.B(n_876),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1144),
.B(n_1115),
.Y(n_1279)
);

NOR3xp33_ASAP7_75t_SL g1280 ( 
.A(n_1152),
.B(n_943),
.C(n_859),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1122),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1114),
.Y(n_1282)
);

INVx6_ASAP7_75t_L g1283 ( 
.A(n_984),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_R g1284 ( 
.A(n_1111),
.B(n_859),
.Y(n_1284)
);

NOR2xp67_ASAP7_75t_L g1285 ( 
.A(n_1132),
.B(n_803),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1132),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1019),
.B(n_803),
.Y(n_1287)
);

NOR3xp33_ASAP7_75t_SL g1288 ( 
.A(n_999),
.B(n_859),
.C(n_85),
.Y(n_1288)
);

NOR3xp33_ASAP7_75t_SL g1289 ( 
.A(n_990),
.B(n_859),
.C(n_85),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1133),
.Y(n_1290)
);

NOR3xp33_ASAP7_75t_SL g1291 ( 
.A(n_1020),
.B(n_86),
.C(n_88),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1140),
.Y(n_1292)
);

BUFx8_ASAP7_75t_L g1293 ( 
.A(n_1129),
.Y(n_1293)
);

INVx6_ASAP7_75t_L g1294 ( 
.A(n_984),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1048),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1034),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1034),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1133),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1106),
.B(n_923),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1286),
.B(n_983),
.Y(n_1300)
);

CKINVDCx11_ASAP7_75t_R g1301 ( 
.A(n_1226),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1178),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1242),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1168),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1198),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1296),
.A2(n_1069),
.B(n_1003),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1218),
.B(n_1148),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1290),
.A2(n_1081),
.B1(n_1080),
.B2(n_1099),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1298),
.B(n_1013),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1209),
.A2(n_1167),
.B(n_1123),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1181),
.A2(n_1003),
.B(n_1060),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1230),
.B(n_1018),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1235),
.A2(n_1166),
.B(n_1087),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1193),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1299),
.A2(n_987),
.B(n_1001),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1202),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1188),
.B(n_1201),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1218),
.A2(n_1151),
.B1(n_1153),
.B2(n_1137),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1262),
.A2(n_1068),
.B(n_1091),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1199),
.B(n_1022),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1296),
.A2(n_1093),
.B(n_1109),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1297),
.A2(n_1139),
.B(n_1040),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1297),
.A2(n_1008),
.B(n_1055),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1295),
.A2(n_1059),
.B(n_1030),
.Y(n_1324)
);

AOI21xp33_ASAP7_75t_L g1325 ( 
.A1(n_1200),
.A2(n_1042),
.B(n_1088),
.Y(n_1325)
);

AOI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1227),
.A2(n_1285),
.B1(n_1216),
.B2(n_1292),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1279),
.A2(n_1050),
.B(n_1029),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1222),
.B(n_1187),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1203),
.Y(n_1329)
);

OAI22x1_ASAP7_75t_L g1330 ( 
.A1(n_1211),
.A2(n_1149),
.B1(n_1160),
.B2(n_1147),
.Y(n_1330)
);

NAND3xp33_ASAP7_75t_SL g1331 ( 
.A(n_1248),
.B(n_1079),
.C(n_1105),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1241),
.A2(n_1089),
.B(n_1074),
.Y(n_1332)
);

INVx3_ASAP7_75t_SL g1333 ( 
.A(n_1177),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1211),
.B(n_1138),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1211),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1206),
.B(n_1043),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1259),
.A2(n_770),
.B(n_769),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1208),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1295),
.A2(n_1117),
.B(n_1098),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1283),
.A2(n_1158),
.B1(n_995),
.B2(n_1097),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_SL g1341 ( 
.A1(n_1192),
.A2(n_1102),
.B(n_1094),
.Y(n_1341)
);

NAND2x1p5_ASAP7_75t_L g1342 ( 
.A(n_1192),
.B(n_1061),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_L g1343 ( 
.A1(n_1179),
.A2(n_1006),
.B(n_1057),
.C(n_1031),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1228),
.B(n_1251),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1212),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1220),
.A2(n_794),
.B(n_780),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1293),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1273),
.A2(n_1067),
.B(n_1086),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1294),
.A2(n_1214),
.B1(n_1221),
.B2(n_1250),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1294),
.A2(n_1076),
.B1(n_1035),
.B2(n_1032),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1232),
.A2(n_1038),
.B(n_1036),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1236),
.A2(n_842),
.B(n_827),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1287),
.A2(n_963),
.B(n_960),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1183),
.B(n_1189),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1182),
.B(n_1041),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1237),
.A2(n_1005),
.B(n_998),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1171),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1186),
.A2(n_979),
.B(n_968),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1204),
.A2(n_1113),
.B(n_1108),
.Y(n_1359)
);

AO21x1_ASAP7_75t_L g1360 ( 
.A1(n_1224),
.A2(n_790),
.B(n_988),
.Y(n_1360)
);

NAND2xp33_ASAP7_75t_L g1361 ( 
.A(n_1284),
.B(n_1034),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1217),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1239),
.A2(n_850),
.B(n_848),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1179),
.A2(n_982),
.B(n_1118),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1186),
.A2(n_1034),
.B(n_779),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1255),
.A2(n_846),
.B(n_844),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1170),
.B(n_1180),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1255),
.A2(n_876),
.B(n_863),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1194),
.B(n_1023),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1293),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1246),
.B(n_1077),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1260),
.A2(n_879),
.B(n_878),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1258),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1245),
.A2(n_1011),
.B(n_1004),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_L g1375 ( 
.A(n_1267),
.B(n_790),
.Y(n_1375)
);

AO31x2_ASAP7_75t_L g1376 ( 
.A1(n_1244),
.A2(n_872),
.A3(n_824),
.B(n_91),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1196),
.B(n_872),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1282),
.Y(n_1378)
);

BUFx8_ASAP7_75t_SL g1379 ( 
.A(n_1370),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1352),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1326),
.A2(n_1210),
.B1(n_1288),
.B2(n_1243),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1306),
.A2(n_1256),
.B(n_1269),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1301),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1344),
.B(n_1195),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1333),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1322),
.A2(n_1272),
.B(n_1270),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1321),
.A2(n_1257),
.B(n_1233),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1347),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1302),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1367),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1354),
.B(n_1175),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1314),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1357),
.B(n_1171),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1313),
.A2(n_1280),
.B(n_1247),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1352),
.Y(n_1395)
);

NOR2x1_ASAP7_75t_L g1396 ( 
.A(n_1361),
.B(n_1205),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1304),
.Y(n_1397)
);

BUFx2_ASAP7_75t_SL g1398 ( 
.A(n_1375),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1320),
.A2(n_1276),
.B(n_1190),
.C(n_1252),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1314),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1331),
.A2(n_1263),
.B(n_1215),
.C(n_1266),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1305),
.B(n_1264),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1316),
.B(n_1275),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1364),
.A2(n_1191),
.B(n_1249),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1357),
.B(n_1171),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1303),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1326),
.A2(n_1289),
.B1(n_1291),
.B2(n_1231),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1336),
.B(n_1229),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1311),
.A2(n_1268),
.B(n_1278),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1378),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1353),
.A2(n_1169),
.B(n_1185),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1335),
.Y(n_1412)
);

AOI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1309),
.A2(n_1234),
.B1(n_1225),
.B2(n_1219),
.C(n_1172),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1357),
.B(n_1185),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1341),
.A2(n_1169),
.B(n_1185),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1373),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1328),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1332),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1329),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1376),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1376),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1389),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_SL g1423 ( 
.A(n_1388),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1384),
.A2(n_1318),
.B1(n_1300),
.B2(n_1356),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1407),
.A2(n_1308),
.B1(n_1349),
.B2(n_1312),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1417),
.B(n_1338),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1389),
.Y(n_1427)
);

CKINVDCx16_ASAP7_75t_R g1428 ( 
.A(n_1385),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1381),
.A2(n_1408),
.B1(n_1391),
.B2(n_1413),
.Y(n_1429)
);

CKINVDCx16_ASAP7_75t_R g1430 ( 
.A(n_1383),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1380),
.A2(n_1315),
.B(n_1360),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1400),
.A2(n_1398),
.B1(n_1308),
.B2(n_1392),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1406),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1398),
.A2(n_1340),
.B1(n_1369),
.B2(n_1355),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1401),
.B(n_1371),
.Y(n_1435)
);

BUFx8_ASAP7_75t_L g1436 ( 
.A(n_1379),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1380),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1388),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1395),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1402),
.B(n_1317),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1412),
.Y(n_1441)
);

BUFx12f_ASAP7_75t_L g1442 ( 
.A(n_1390),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1396),
.B(n_1415),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1395),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1390),
.B(n_1334),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1399),
.A2(n_1343),
.B(n_1339),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1406),
.A2(n_1207),
.B1(n_1225),
.B2(n_1367),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1419),
.B(n_1345),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1397),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1410),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1429),
.A2(n_1396),
.B1(n_1419),
.B2(n_1416),
.Y(n_1451)
);

BUFx12f_ASAP7_75t_L g1452 ( 
.A(n_1436),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1426),
.B(n_1410),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1422),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1435),
.A2(n_1425),
.B1(n_1424),
.B2(n_1429),
.Y(n_1455)
);

OAI211xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1424),
.A2(n_1176),
.B(n_1416),
.C(n_1351),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1435),
.A2(n_1351),
.B(n_1325),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1425),
.A2(n_1397),
.B1(n_1377),
.B2(n_1342),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1434),
.A2(n_1327),
.B1(n_1350),
.B2(n_1330),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1448),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1439),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1431),
.A2(n_1415),
.B(n_1420),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1442),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1443),
.B(n_1420),
.Y(n_1464)
);

AOI222xp33_ASAP7_75t_L g1465 ( 
.A1(n_1432),
.A2(n_1403),
.B1(n_1402),
.B2(n_1362),
.C1(n_1356),
.C2(n_1348),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1438),
.B(n_1223),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1440),
.A2(n_1403),
.B1(n_1348),
.B2(n_1394),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1438),
.A2(n_1394),
.B1(n_1307),
.B2(n_1310),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1442),
.A2(n_1421),
.B1(n_1409),
.B2(n_1394),
.Y(n_1469)
);

OAI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1447),
.A2(n_1254),
.B1(n_1271),
.B2(n_1421),
.C(n_1174),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1428),
.A2(n_1173),
.B1(n_1180),
.B2(n_1254),
.Y(n_1471)
);

NAND2x1_ASAP7_75t_L g1472 ( 
.A(n_1443),
.B(n_1393),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1436),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1446),
.A2(n_1411),
.B(n_1404),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1427),
.A2(n_1409),
.B1(n_1278),
.B2(n_1315),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1475),
.B(n_1461),
.Y(n_1476)
);

NOR2x1_ASAP7_75t_L g1477 ( 
.A(n_1463),
.B(n_1443),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1475),
.B(n_1439),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1454),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1461),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1460),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1464),
.B(n_1437),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1472),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1464),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1474),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1467),
.B(n_1437),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1467),
.B(n_1444),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1453),
.B(n_1433),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1469),
.B(n_1444),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1463),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1474),
.B(n_1450),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1474),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1462),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1457),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1468),
.B(n_1449),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1458),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1494),
.B(n_1455),
.C(n_1465),
.Y(n_1497)
);

OAI332xp33_ASAP7_75t_L g1498 ( 
.A1(n_1494),
.A2(n_1430),
.A3(n_1441),
.B1(n_1471),
.B2(n_1451),
.B3(n_1455),
.C1(n_1470),
.C2(n_1466),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1481),
.B(n_1468),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1484),
.B(n_1482),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1494),
.A2(n_1456),
.B1(n_1459),
.B2(n_1445),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_R g1502 ( 
.A(n_1490),
.B(n_1473),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_L g1503 ( 
.A(n_1496),
.B(n_1409),
.C(n_1449),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1479),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_L g1505 ( 
.A(n_1477),
.B(n_1423),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1479),
.Y(n_1506)
);

OAI33xp33_ASAP7_75t_L g1507 ( 
.A1(n_1488),
.A2(n_1480),
.A3(n_1493),
.B1(n_1492),
.B2(n_1485),
.B3(n_1452),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1496),
.A2(n_1445),
.B1(n_1409),
.B2(n_1334),
.Y(n_1508)
);

OR2x6_ASAP7_75t_L g1509 ( 
.A(n_1477),
.B(n_1483),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1499),
.B(n_1488),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1504),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1500),
.B(n_1484),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1497),
.A2(n_1476),
.B1(n_1487),
.B2(n_1486),
.Y(n_1513)
);

NOR2x1_ASAP7_75t_L g1514 ( 
.A(n_1505),
.B(n_1509),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1502),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1506),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1509),
.Y(n_1517)
);

NOR2x1_ASAP7_75t_L g1518 ( 
.A(n_1509),
.B(n_1483),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1498),
.B(n_1480),
.Y(n_1519)
);

NAND2x1_ASAP7_75t_L g1520 ( 
.A(n_1503),
.B(n_1483),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1508),
.B(n_1484),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1501),
.B(n_1484),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1507),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1504),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1504),
.Y(n_1525)
);

AOI211xp5_ASAP7_75t_L g1526 ( 
.A1(n_1515),
.A2(n_1476),
.B(n_1489),
.C(n_1483),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1510),
.Y(n_1527)
);

AOI32xp33_ASAP7_75t_L g1528 ( 
.A1(n_1514),
.A2(n_1489),
.A3(n_1487),
.B1(n_1486),
.B2(n_1478),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1511),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1522),
.B(n_1491),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1523),
.A2(n_1492),
.B(n_1485),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1513),
.B(n_1491),
.Y(n_1532)
);

NOR3xp33_ASAP7_75t_L g1533 ( 
.A(n_1526),
.B(n_1519),
.C(n_1520),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1527),
.Y(n_1534)
);

NAND2xp33_ASAP7_75t_SL g1535 ( 
.A(n_1532),
.B(n_1513),
.Y(n_1535)
);

OAI211xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1528),
.A2(n_1519),
.B(n_1517),
.C(n_1518),
.Y(n_1536)
);

NAND2x1_ASAP7_75t_L g1537 ( 
.A(n_1533),
.B(n_1531),
.Y(n_1537)
);

AOI31xp33_ASAP7_75t_L g1538 ( 
.A1(n_1535),
.A2(n_1532),
.A3(n_1521),
.B(n_1530),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1538),
.B(n_1536),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1537),
.A2(n_1534),
.B1(n_1531),
.B2(n_1529),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1538),
.B(n_1529),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1537),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1541),
.B(n_1512),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1542),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1540),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1539),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1542),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1541),
.B(n_1511),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1548),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1547),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1547),
.B(n_1516),
.Y(n_1551)
);

OAI21xp33_ASAP7_75t_L g1552 ( 
.A1(n_1545),
.A2(n_1525),
.B(n_1524),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1543),
.B(n_1544),
.Y(n_1553)
);

NOR2x1_ASAP7_75t_L g1554 ( 
.A(n_1546),
.B(n_1184),
.Y(n_1554)
);

O2A1O1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1550),
.A2(n_1184),
.B(n_1213),
.C(n_1363),
.Y(n_1555)
);

O2A1O1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1549),
.A2(n_1213),
.B(n_1372),
.C(n_1375),
.Y(n_1556)
);

NAND3xp33_ASAP7_75t_L g1557 ( 
.A(n_1554),
.B(n_1267),
.C(n_1372),
.Y(n_1557)
);

OAI221xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1551),
.A2(n_1495),
.B1(n_1253),
.B2(n_1319),
.C(n_1359),
.Y(n_1558)
);

O2A1O1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1552),
.A2(n_93),
.B(n_90),
.C(n_92),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1550),
.Y(n_1560)
);

OA22x2_ASAP7_75t_L g1561 ( 
.A1(n_1550),
.A2(n_1482),
.B1(n_1393),
.B2(n_1414),
.Y(n_1561)
);

OAI221xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1553),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.C(n_98),
.Y(n_1562)
);

AOI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1550),
.A2(n_1482),
.B1(n_1324),
.B2(n_1418),
.C(n_1405),
.Y(n_1563)
);

AOI21xp33_ASAP7_75t_L g1564 ( 
.A1(n_1550),
.A2(n_97),
.B(n_99),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1550),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1560),
.A2(n_1374),
.B(n_102),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1565),
.A2(n_1482),
.B1(n_1274),
.B2(n_1414),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1561),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_R g1569 ( 
.A(n_1562),
.B(n_102),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1559),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1557),
.A2(n_1558),
.B1(n_1555),
.B2(n_1556),
.Y(n_1571)
);

BUFx12f_ASAP7_75t_L g1572 ( 
.A(n_1564),
.Y(n_1572)
);

NOR3xp33_ASAP7_75t_L g1573 ( 
.A(n_1563),
.B(n_103),
.C(n_104),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1560),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1565),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1560),
.A2(n_104),
.B(n_1414),
.C(n_1405),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_SL g1577 ( 
.A(n_1569),
.B(n_120),
.C(n_123),
.Y(n_1577)
);

NOR2x1_ASAP7_75t_L g1578 ( 
.A(n_1575),
.B(n_1323),
.Y(n_1578)
);

NOR3xp33_ASAP7_75t_L g1579 ( 
.A(n_1570),
.B(n_1368),
.C(n_1405),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1574),
.Y(n_1580)
);

AO22x2_ASAP7_75t_L g1581 ( 
.A1(n_1572),
.A2(n_1418),
.B1(n_1274),
.B2(n_1323),
.Y(n_1581)
);

NAND3xp33_ASAP7_75t_L g1582 ( 
.A(n_1574),
.B(n_1238),
.C(n_1197),
.Y(n_1582)
);

NOR2x1_ASAP7_75t_L g1583 ( 
.A(n_1568),
.B(n_872),
.Y(n_1583)
);

NOR3xp33_ASAP7_75t_L g1584 ( 
.A(n_1576),
.B(n_1365),
.C(n_1358),
.Y(n_1584)
);

NAND4xp75_ASAP7_75t_L g1585 ( 
.A(n_1566),
.B(n_124),
.C(n_125),
.D(n_127),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1573),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1571),
.A2(n_1382),
.B1(n_1386),
.B2(n_1238),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1567),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1580),
.B(n_1382),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_L g1590 ( 
.A(n_1577),
.B(n_1366),
.C(n_128),
.Y(n_1590)
);

XNOR2xp5_ASAP7_75t_L g1591 ( 
.A(n_1585),
.B(n_130),
.Y(n_1591)
);

OR3x2_ASAP7_75t_L g1592 ( 
.A(n_1586),
.B(n_131),
.C(n_135),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1583),
.A2(n_1261),
.B(n_1240),
.Y(n_1593)
);

XNOR2xp5_ASAP7_75t_L g1594 ( 
.A(n_1588),
.B(n_137),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1578),
.A2(n_1587),
.B1(n_1584),
.B2(n_1582),
.Y(n_1595)
);

OAI211xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1579),
.A2(n_139),
.B(n_141),
.C(n_143),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_SL g1597 ( 
.A(n_1581),
.B(n_147),
.C(n_150),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1590),
.B(n_156),
.Y(n_1598)
);

XNOR2x1_ASAP7_75t_SL g1599 ( 
.A(n_1594),
.B(n_158),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1591),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1595),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1589),
.Y(n_1602)
);

AOI211xp5_ASAP7_75t_L g1603 ( 
.A1(n_1596),
.A2(n_1277),
.B(n_1261),
.C(n_1265),
.Y(n_1603)
);

AOI211xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1601),
.A2(n_1597),
.B(n_1592),
.C(n_1593),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1600),
.A2(n_1281),
.B1(n_1261),
.B2(n_1265),
.Y(n_1605)
);

OA22x2_ASAP7_75t_L g1606 ( 
.A1(n_1602),
.A2(n_1387),
.B1(n_1411),
.B2(n_1346),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1604),
.A2(n_1598),
.B(n_1599),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1605),
.A2(n_1603),
.B(n_1337),
.Y(n_1608)
);

NOR2x1p5_ASAP7_75t_L g1609 ( 
.A(n_1607),
.B(n_1606),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1608),
.Y(n_1610)
);

OAI31xp33_ASAP7_75t_L g1611 ( 
.A1(n_1609),
.A2(n_162),
.A3(n_164),
.B(n_165),
.Y(n_1611)
);

OAI22x1_ASAP7_75t_L g1612 ( 
.A1(n_1611),
.A2(n_1610),
.B1(n_172),
.B2(n_173),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1612),
.A2(n_178),
.B1(n_185),
.B2(n_186),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1613),
.A2(n_187),
.B1(n_188),
.B2(n_192),
.C(n_194),
.Y(n_1614)
);

AOI211xp5_ASAP7_75t_L g1615 ( 
.A1(n_1614),
.A2(n_197),
.B(n_198),
.C(n_199),
.Y(n_1615)
);


endmodule