module fake_jpeg_31841_n_545 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_545);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_545;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_56),
.Y(n_170)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_18),
.A2(n_36),
.B1(n_39),
.B2(n_42),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_60),
.A2(n_16),
.B1(n_23),
.B2(n_27),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_108),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_64),
.Y(n_161)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_66),
.Y(n_169)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_18),
.B(n_14),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_104),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_82),
.Y(n_173)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_94),
.Y(n_124)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g176 ( 
.A(n_95),
.Y(n_176)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_97),
.Y(n_136)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_103),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g145 ( 
.A(n_105),
.B(n_107),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_106),
.A2(n_27),
.B1(n_49),
.B2(n_22),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_109),
.B(n_118),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_36),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_81),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_121),
.B(n_125),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_56),
.B(n_39),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_42),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_126),
.B(n_130),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_29),
.B(n_30),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_128),
.A2(n_49),
.A3(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_61),
.A2(n_26),
.B1(n_47),
.B2(n_37),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_129),
.A2(n_132),
.B1(n_140),
.B2(n_160),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_63),
.A2(n_37),
.B1(n_47),
.B2(n_43),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_52),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_139),
.B(n_155),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_98),
.B(n_52),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_101),
.B(n_21),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_72),
.B(n_21),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_165),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_91),
.A2(n_27),
.B1(n_47),
.B2(n_43),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_102),
.B(n_23),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_16),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_172),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_44),
.B1(n_14),
.B2(n_13),
.Y(n_220)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_111),
.A2(n_75),
.B1(n_66),
.B2(n_92),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_178),
.A2(n_192),
.B1(n_204),
.B2(n_206),
.Y(n_237)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_117),
.Y(n_181)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_22),
.C(n_104),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_183),
.B(n_188),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_32),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_203),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

INVx11_ASAP7_75t_L g274 ( 
.A(n_186),
.Y(n_274)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_22),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_106),
.C(n_89),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_189),
.B(n_201),
.Y(n_247)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_119),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_191),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_68),
.B1(n_78),
.B2(n_74),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_195),
.A2(n_211),
.B(n_213),
.Y(n_268)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_145),
.A2(n_31),
.A3(n_45),
.B1(n_33),
.B2(n_64),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_118),
.B(n_45),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_160),
.A2(n_84),
.B1(n_73),
.B2(n_69),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_47),
.B1(n_43),
.B2(n_37),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_122),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_209),
.B(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_43),
.B1(n_37),
.B2(n_45),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_176),
.A2(n_33),
.B1(n_25),
.B2(n_38),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_110),
.A2(n_33),
.B1(n_25),
.B2(n_38),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_215),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_233)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_216),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_120),
.A2(n_25),
.B1(n_38),
.B2(n_13),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_218),
.A2(n_131),
.B1(n_147),
.B2(n_154),
.Y(n_253)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g264 ( 
.A1(n_220),
.A2(n_223),
.B1(n_147),
.B2(n_131),
.Y(n_264)
);

BUFx4f_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_224),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_130),
.A2(n_136),
.B1(n_124),
.B2(n_153),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_152),
.B(n_0),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_115),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_143),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_120),
.B(n_14),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_232),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_140),
.A2(n_44),
.B1(n_13),
.B2(n_12),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_230),
.A2(n_231),
.B1(n_10),
.B2(n_1),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_141),
.A2(n_11),
.B1(n_10),
.B2(n_44),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_119),
.B1(n_123),
.B2(n_135),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_235),
.A2(n_255),
.B(n_264),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_194),
.A2(n_124),
.B1(n_136),
.B2(n_135),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_238),
.A2(n_223),
.B(n_204),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_146),
.C(n_11),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_220),
.Y(n_283)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_195),
.A2(n_170),
.B(n_137),
.C(n_112),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_251),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_180),
.A2(n_141),
.B1(n_169),
.B2(n_161),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_252),
.A2(n_263),
.B1(n_197),
.B2(n_188),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_253),
.A2(n_221),
.B1(n_191),
.B2(n_168),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_179),
.A2(n_137),
.B1(n_113),
.B2(n_116),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_169),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_269),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_180),
.A2(n_163),
.B1(n_162),
.B2(n_150),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_168),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_271),
.A2(n_185),
.B1(n_198),
.B2(n_216),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_205),
.A2(n_10),
.B(n_138),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_SL g286 ( 
.A(n_273),
.B(n_275),
.C(n_221),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g275 ( 
.A1(n_184),
.A2(n_113),
.B(n_168),
.C(n_114),
.D(n_44),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_277),
.A2(n_286),
.B(n_272),
.Y(n_330)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_282),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_247),
.A2(n_203),
.B(n_183),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_281),
.A2(n_286),
.B(n_289),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_251),
.B(n_264),
.C(n_201),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_285),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g287 ( 
.A1(n_234),
.A2(n_228),
.A3(n_217),
.B1(n_214),
.B2(n_210),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_290),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_288),
.A2(n_289),
.B1(n_296),
.B2(n_237),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_265),
.A2(n_230),
.B1(n_188),
.B2(n_189),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_296),
.B1(n_238),
.B2(n_233),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_222),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_293),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_234),
.B(n_207),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_244),
.B(n_262),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_298),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_190),
.C(n_187),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_264),
.C(n_252),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_265),
.A2(n_202),
.B1(n_181),
.B2(n_196),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_297),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_237),
.A2(n_182),
.B1(n_212),
.B2(n_232),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_302),
.Y(n_322)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_301),
.Y(n_327)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_250),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_226),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_225),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_304),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_261),
.B(n_227),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_199),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_305),
.B(n_248),
.Y(n_335)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_246),
.Y(n_334)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_307),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_276),
.Y(n_309)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_310),
.A2(n_323),
.B1(n_328),
.B2(n_331),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_275),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_311),
.B(n_312),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_263),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_303),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_329),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_333),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_308),
.A2(n_271),
.B1(n_264),
.B2(n_242),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_304),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g357 ( 
.A1(n_330),
.A2(n_291),
.B(n_295),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_308),
.A2(n_242),
.B1(n_246),
.B2(n_245),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_305),
.A2(n_272),
.B1(n_267),
.B2(n_261),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_332),
.A2(n_300),
.B1(n_297),
.B2(n_284),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_278),
.B(n_267),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_334),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_296),
.Y(n_340)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_354),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_282),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g380 ( 
.A1(n_342),
.A2(n_349),
.B(n_343),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_287),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_344),
.B(n_312),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_325),
.A2(n_288),
.B1(n_282),
.B2(n_292),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_345),
.A2(n_312),
.B1(n_328),
.B2(n_311),
.Y(n_378)
);

OAI21xp33_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_293),
.B(n_302),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g387 ( 
.A1(n_346),
.A2(n_336),
.B(n_334),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_313),
.A2(n_277),
.B(n_283),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_347),
.A2(n_357),
.B(n_335),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_R g349 ( 
.A(n_330),
.B(n_281),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_318),
.A2(n_288),
.B1(n_291),
.B2(n_298),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_351),
.A2(n_322),
.B1(n_325),
.B2(n_321),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_278),
.Y(n_352)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_353),
.Y(n_371)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_337),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_331),
.A2(n_299),
.B1(n_291),
.B2(n_279),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_358),
.A2(n_359),
.B1(n_360),
.B2(n_362),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_310),
.A2(n_295),
.B1(n_306),
.B2(n_301),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_317),
.B(n_307),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_364),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_323),
.A2(n_306),
.B1(n_301),
.B2(n_245),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_276),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_327),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_329),
.Y(n_375)
);

BUFx8_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_369),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_347),
.A2(n_315),
.B(n_321),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_361),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_367),
.B(n_314),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_374),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_380),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_333),
.C(n_311),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_385),
.C(n_386),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_377),
.A2(n_392),
.B(n_342),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_378),
.B(n_397),
.Y(n_418)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_381),
.A2(n_383),
.B1(n_359),
.B2(n_350),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_348),
.B(n_333),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_387),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_355),
.A2(n_322),
.B1(n_336),
.B2(n_326),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_365),
.C(n_345),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_326),
.C(n_327),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_355),
.A2(n_338),
.B1(n_320),
.B2(n_309),
.Y(n_388)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_388),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_338),
.B1(n_324),
.B2(n_320),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_363),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_309),
.B(n_320),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_324),
.C(n_241),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_382),
.C(n_385),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_248),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_339),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_343),
.B(n_324),
.Y(n_396)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_352),
.B(n_256),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_399),
.A2(n_407),
.B1(n_415),
.B2(n_421),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_401),
.A2(n_405),
.B(n_413),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_396),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_414),
.Y(n_430)
);

AO22x1_ASAP7_75t_L g405 ( 
.A1(n_380),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_405)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_408),
.Y(n_432)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_410),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_349),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_425),
.C(n_193),
.Y(n_444)
);

BUFx12_ASAP7_75t_L g414 ( 
.A(n_380),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_370),
.A2(n_362),
.B1(n_364),
.B2(n_354),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_378),
.Y(n_429)
);

NAND2x1_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_395),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_417),
.B(n_394),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_256),
.Y(n_419)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_370),
.A2(n_356),
.B1(n_353),
.B2(n_258),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_368),
.Y(n_422)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_422),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_383),
.A2(n_356),
.B1(n_258),
.B2(n_254),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_423),
.A2(n_371),
.B1(n_274),
.B2(n_266),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_285),
.Y(n_424)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_424),
.Y(n_440)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_393),
.Y(n_426)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_426),
.Y(n_445)
);

XNOR2x1_ASAP7_75t_SL g428 ( 
.A(n_417),
.B(n_373),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_428),
.B(n_429),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_384),
.B1(n_390),
.B2(n_387),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_433),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_401),
.A2(n_384),
.B(n_392),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_393),
.Y(n_434)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_443),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_389),
.Y(n_436)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_372),
.B1(n_389),
.B2(n_371),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_450),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_409),
.B(n_372),
.Y(n_442)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_391),
.Y(n_443)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_424),
.C(n_423),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_446),
.A2(n_405),
.B1(n_410),
.B2(n_422),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_239),
.C(n_243),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_407),
.C(n_416),
.Y(n_459)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_420),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_449),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_418),
.A2(n_369),
.B1(n_266),
.B2(n_274),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_448),
.Y(n_451)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_452),
.A2(n_441),
.B1(n_431),
.B2(n_449),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_404),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_467),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_461),
.C(n_468),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_438),
.A2(n_398),
.B1(n_405),
.B2(n_400),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_428),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_412),
.C(n_400),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_434),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_462),
.B(n_442),
.Y(n_476)
);

FAx1_ASAP7_75t_SL g464 ( 
.A(n_439),
.B(n_414),
.CI(n_399),
.CON(n_464),
.SN(n_464)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_465),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_414),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_415),
.C(n_421),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_454),
.A2(n_438),
.B1(n_470),
.B2(n_466),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_474),
.A2(n_460),
.B1(n_468),
.B2(n_457),
.Y(n_492)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_476),
.Y(n_489)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_455),
.Y(n_477)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_477),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_456),
.C(n_461),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_483),
.C(n_484),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_240),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_463),
.A2(n_433),
.B(n_430),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_480),
.A2(n_475),
.B(n_479),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_481),
.A2(n_369),
.B1(n_239),
.B2(n_186),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_437),
.Y(n_482)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_429),
.C(n_439),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_440),
.C(n_437),
.Y(n_484)
);

AOI21x1_ASAP7_75t_L g485 ( 
.A1(n_464),
.A2(n_445),
.B(n_440),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_485),
.A2(n_369),
.B(n_243),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_452),
.A2(n_445),
.B1(n_450),
.B2(n_427),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_219),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_446),
.C(n_406),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_240),
.C(n_114),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_478),
.B(n_464),
.Y(n_491)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_491),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_492),
.B(n_493),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_457),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_494),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_495),
.B(n_496),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_497),
.B(n_498),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_488),
.B(n_177),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_500),
.B(n_501),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_471),
.B(n_44),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_502),
.A2(n_504),
.B(n_480),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_475),
.A2(n_0),
.B(n_1),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_505),
.B(n_507),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_489),
.A2(n_474),
.B1(n_484),
.B2(n_485),
.Y(n_507)
);

OAI21xp33_ASAP7_75t_L g510 ( 
.A1(n_503),
.A2(n_482),
.B(n_481),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_496),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_471),
.C(n_488),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_518),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_492),
.A2(n_472),
.B1(n_473),
.B2(n_483),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_495),
.Y(n_525)
);

OA21x2_ASAP7_75t_SL g515 ( 
.A1(n_502),
.A2(n_1),
.B(n_2),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_515),
.A2(n_504),
.B(n_4),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_490),
.A2(n_1),
.B(n_2),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_516),
.A2(n_497),
.B(n_4),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_494),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_508),
.A2(n_499),
.B(n_500),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_528),
.B(n_513),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_522),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_527),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_526),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_506),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_511),
.B(n_3),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_3),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_530),
.B(n_525),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_524),
.A2(n_517),
.B(n_512),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_533),
.B(n_529),
.C(n_532),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_524),
.A2(n_507),
.B(n_509),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_534),
.A2(n_510),
.B(n_518),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_R g535 ( 
.A(n_531),
.B(n_521),
.Y(n_535)
);

O2A1O1Ixp33_ASAP7_75t_SL g539 ( 
.A1(n_535),
.A2(n_536),
.B(n_537),
.C(n_5),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_5),
.C(n_6),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_539),
.Y(n_541)
);

NOR5xp2_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_540),
.C(n_6),
.D(n_7),
.E(n_9),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_542),
.A2(n_5),
.B(n_7),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_7),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_7),
.Y(n_545)
);


endmodule