module fake_jpeg_30318_n_371 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_371);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_371;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_7),
.B(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_55),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_65),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_30),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_27),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_27),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_78),
.Y(n_112)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_32),
.B1(n_25),
.B2(n_29),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_32),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_67),
.Y(n_85)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_85),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_92),
.B(n_94),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_57),
.B(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_35),
.B1(n_34),
.B2(n_48),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_76),
.B1(n_67),
.B2(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_59),
.B(n_40),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_29),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

BUFx4f_ASAP7_75t_SL g137 ( 
.A(n_115),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_46),
.B(n_51),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_121),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_127),
.Y(n_157)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_80),
.A2(n_32),
.B1(n_47),
.B2(n_44),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_35),
.B1(n_77),
.B2(n_60),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_140),
.B1(n_95),
.B2(n_82),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_96),
.A2(n_38),
.B1(n_44),
.B2(n_47),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_72),
.B1(n_56),
.B2(n_54),
.Y(n_168)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

HAxp5_ASAP7_75t_SL g138 ( 
.A(n_81),
.B(n_68),
.CON(n_138),
.SN(n_138)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_63),
.Y(n_169)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_35),
.B1(n_55),
.B2(n_75),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_144),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_78),
.C(n_74),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_65),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_149),
.Y(n_166)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_114),
.B1(n_55),
.B2(n_95),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_168),
.A2(n_123),
.B1(n_104),
.B2(n_98),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_62),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_141),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_136),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_82),
.B1(n_144),
.B2(n_134),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_120),
.B(n_145),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_185),
.B(n_137),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_153),
.B1(n_170),
.B2(n_154),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_178),
.B(n_192),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_188),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_181),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_132),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_118),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_120),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_186),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_124),
.B(n_128),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_127),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_130),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_123),
.B(n_139),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_137),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_126),
.B(n_143),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_155),
.C(n_152),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_173),
.B1(n_167),
.B2(n_162),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_194),
.B1(n_188),
.B2(n_185),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_151),
.C(n_152),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_192),
.C(n_161),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_183),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_182),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_179),
.A2(n_168),
.B1(n_104),
.B2(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_213),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_170),
.B1(n_160),
.B2(n_142),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_205),
.B1(n_215),
.B2(n_158),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_167),
.B1(n_154),
.B2(n_153),
.Y(n_206)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_185),
.B(n_175),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_174),
.B(n_151),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_164),
.B1(n_158),
.B2(n_64),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_184),
.B(n_192),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_199),
.B(n_137),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_178),
.C(n_180),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_195),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_193),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_222),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_224),
.A2(n_150),
.B(n_23),
.Y(n_257)
);

INVx13_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_200),
.C(n_208),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_191),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_228),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_216),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_209),
.B(n_210),
.Y(n_230)
);

NOR4xp25_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_209),
.C(n_197),
.D(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_191),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_203),
.B1(n_197),
.B2(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_237),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_176),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_256),
.B1(n_231),
.B2(n_229),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_197),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_242),
.B(n_255),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_217),
.C(n_232),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_253),
.B(n_254),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_222),
.A2(n_211),
.B(n_207),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_199),
.B(n_205),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_167),
.B1(n_161),
.B2(n_150),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_257),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_233),
.B1(n_221),
.B2(n_220),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_181),
.B1(n_225),
.B2(n_148),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_275),
.C(n_256),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_220),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_244),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_227),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_266),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_223),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_271),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_225),
.B1(n_122),
.B2(n_103),
.Y(n_291)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_274),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_223),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_273),
.B(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_229),
.C(n_236),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_240),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_279),
.B1(n_252),
.B2(n_255),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_246),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_252),
.C(n_257),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_281),
.A2(n_280),
.B(n_297),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_289),
.Y(n_314)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

AND3x1_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_248),
.C(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_290),
.C(n_294),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_223),
.B1(n_181),
.B2(n_28),
.Y(n_288)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_164),
.C(n_23),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_265),
.A2(n_41),
.B(n_51),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_298),
.B(n_300),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_41),
.C(n_125),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_273),
.A2(n_159),
.B(n_103),
.C(n_149),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_113),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_38),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_50),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_262),
.B1(n_275),
.B2(n_269),
.Y(n_300)
);

AO221x1_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_278),
.B1(n_159),
.B2(n_13),
.C(n_19),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_303),
.Y(n_324)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_308),
.A2(n_310),
.B1(n_37),
.B2(n_25),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_278),
.B(n_17),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_40),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_113),
.C(n_116),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_286),
.C(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_321),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_318),
.B(n_320),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_298),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_323),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_285),
.C(n_295),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_28),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_307),
.A2(n_295),
.B(n_50),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_322),
.B(n_326),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_316),
.A2(n_295),
.B1(n_37),
.B2(n_34),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_114),
.C(n_79),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_313),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_306),
.B1(n_312),
.B2(n_309),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_330),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_301),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_320),
.A2(n_312),
.B1(n_316),
.B2(n_302),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_331),
.A2(n_326),
.B1(n_16),
.B2(n_3),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_315),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_339),
.Y(n_349)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

AOI221xp5_ASAP7_75t_L g338 ( 
.A1(n_322),
.A2(n_48),
.B1(n_42),
.B2(n_3),
.C(n_4),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_338),
.A2(n_1),
.B(n_2),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_42),
.C(n_106),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_16),
.C(n_2),
.Y(n_340)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_340),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_338),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_341),
.B(n_350),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_335),
.B(n_325),
.Y(n_343)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_343),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_344),
.B(n_337),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_SL g346 ( 
.A(n_336),
.B(n_106),
.Y(n_346)
);

OAI33xp33_ASAP7_75t_L g354 ( 
.A1(n_346),
.A2(n_115),
.A3(n_49),
.B1(n_6),
.B2(n_7),
.B3(n_8),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_348),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_87),
.C(n_71),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_352),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_342),
.A2(n_336),
.B1(n_340),
.B2(n_6),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_71),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_357),
.Y(n_360)
);

AOI21x1_ASAP7_75t_SL g358 ( 
.A1(n_354),
.A2(n_347),
.B(n_9),
.Y(n_358)
);

OAI21x1_ASAP7_75t_L g365 ( 
.A1(n_358),
.A2(n_361),
.B(n_5),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_355),
.B(n_345),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_356),
.A2(n_350),
.B(n_346),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_362),
.B(n_351),
.C(n_10),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_365),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_359),
.A2(n_5),
.B(n_10),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_360),
.C(n_12),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_L g368 ( 
.A1(n_367),
.A2(n_115),
.A3(n_71),
.B1(n_12),
.B2(n_11),
.C1(n_49),
.C2(n_83),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_368),
.B(n_366),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_369),
.B(n_83),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_370),
.A2(n_49),
.B(n_359),
.Y(n_371)
);


endmodule