module fake_jpeg_22662_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_46),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_17),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_20),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_68),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_72),
.B(n_76),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_77),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_83),
.B1(n_56),
.B2(n_54),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_79),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_36),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_45),
.B1(n_43),
.B2(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_32),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_86),
.B(n_93),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_30),
.B1(n_43),
.B2(n_37),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_37),
.B1(n_38),
.B2(n_43),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_20),
.B(n_35),
.C(n_39),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_20),
.B(n_35),
.C(n_49),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_20),
.Y(n_90)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_39),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_96),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_97),
.B(n_111),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_37),
.B1(n_38),
.B2(n_20),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_115),
.B1(n_123),
.B2(n_42),
.Y(n_129)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_110),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_109),
.A2(n_118),
.B(n_67),
.Y(n_151)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_36),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_116),
.Y(n_130)
);

OAI22x1_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_35),
.B1(n_27),
.B2(n_40),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_36),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_36),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_125),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_42),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_49),
.B1(n_42),
.B2(n_18),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_44),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_44),
.C(n_41),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_67),
.C(n_90),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_115),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_131),
.B(n_147),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_146),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_134),
.B1(n_74),
.B2(n_102),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_69),
.B(n_80),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_89),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_52),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_29),
.B(n_23),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_34),
.B(n_31),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_126),
.B1(n_113),
.B2(n_103),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_44),
.C(n_41),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_141),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_91),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_70),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_74),
.Y(n_166)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_40),
.A3(n_41),
.B1(n_44),
.B2(n_49),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_122),
.B1(n_107),
.B2(n_66),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_152),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_52),
.B(n_27),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_100),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_108),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_168),
.B1(n_169),
.B2(n_174),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_152),
.A2(n_104),
.B1(n_102),
.B2(n_121),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_186),
.B1(n_151),
.B2(n_132),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_123),
.A3(n_31),
.B1(n_23),
.B2(n_29),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g187 ( 
.A(n_159),
.B(n_176),
.C(n_179),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_162),
.B(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_185),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_99),
.B1(n_77),
.B2(n_95),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_129),
.B1(n_149),
.B2(n_135),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_177),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_175),
.C(n_136),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_122),
.B1(n_88),
.B2(n_108),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_120),
.C(n_41),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_182),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_130),
.A2(n_122),
.B1(n_88),
.B2(n_64),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_183),
.B1(n_148),
.B2(n_146),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_181),
.A2(n_147),
.B1(n_131),
.B2(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_176),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_127),
.A2(n_19),
.B1(n_34),
.B2(n_28),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_188),
.B(n_194),
.Y(n_227)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_68),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_143),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_127),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_205),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_210),
.C(n_217),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_158),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_156),
.B(n_143),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_212),
.B1(n_167),
.B2(n_163),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_161),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_207),
.Y(n_224)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_209),
.Y(n_238)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_136),
.C(n_146),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_155),
.A2(n_22),
.B1(n_33),
.B2(n_28),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_215),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_11),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_19),
.B(n_168),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_160),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_0),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_157),
.B(n_92),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_0),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_218),
.A2(n_26),
.B(n_33),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_11),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_159),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_229),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_175),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_234),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_164),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_241),
.Y(n_258)
);

NOR3xp33_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_187),
.C(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_201),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_0),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_25),
.C(n_22),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_187),
.C(n_216),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_9),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_9),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_204),
.C(n_208),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_1),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_202),
.A2(n_25),
.B1(n_1),
.B2(n_3),
.Y(n_245)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_246),
.B(n_236),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_189),
.C(n_192),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_189),
.C(n_193),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_219),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_263),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_244),
.B1(n_237),
.B2(n_232),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_190),
.B(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_231),
.B1(n_227),
.B2(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_191),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_197),
.C(n_198),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_1),
.Y(n_264)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_229),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_273),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_230),
.B1(n_222),
.B2(n_220),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_274),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_243),
.B1(n_224),
.B2(n_233),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_240),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_276),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_226),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_283),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_247),
.C(n_263),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_2),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_249),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_293),
.C(n_296),
.Y(n_304)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_270),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_248),
.C(n_255),
.Y(n_293)
);

NOR3xp33_ASAP7_75t_SL g294 ( 
.A(n_269),
.B(n_246),
.C(n_252),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_277),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_279),
.C(n_255),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_257),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_251),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_6),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_282),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_300),
.A2(n_310),
.B(n_12),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_309),
.B(n_285),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_278),
.CI(n_250),
.CON(n_302),
.SN(n_302)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_302),
.B(n_306),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_267),
.B1(n_3),
.B2(n_5),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_2),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_2),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_12),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_6),
.C(n_7),
.Y(n_309)
);

XOR2x2_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_6),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_10),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_288),
.B1(n_294),
.B2(n_286),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_316),
.B1(n_311),
.B2(n_306),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_317),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_287),
.B(n_297),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_308),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_302),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_300),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_326),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_327),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_325),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_329),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_330),
.A2(n_321),
.B(n_320),
.C(n_15),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_12),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_13),
.B(n_15),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_15),
.Y(n_338)
);


endmodule