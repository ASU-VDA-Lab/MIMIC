module fake_ariane_980_n_2336 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2336);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2336;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_279;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2271;
wire n_2116;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_348;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1860;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_2315;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_363;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_149),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_47),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_78),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_66),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_15),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_9),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_43),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_42),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_2),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_41),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_3),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_92),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_23),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_102),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_218),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_104),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_126),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_223),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_192),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_188),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_221),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_133),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_205),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_174),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_18),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_110),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_198),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_164),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_75),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_108),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_119),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_56),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_75),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_69),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_78),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_200),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_37),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_166),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_79),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_1),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_224),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_22),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_130),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_180),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_225),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_202),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_148),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_51),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_131),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_41),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_162),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_38),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_155),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_64),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_173),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_147),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_90),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_39),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_216),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_99),
.Y(n_303)
);

BUFx8_ASAP7_75t_SL g304 ( 
.A(n_220),
.Y(n_304)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_168),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_63),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_146),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_123),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_177),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_101),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_124),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_106),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_19),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_232),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_57),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_237),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_158),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_27),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_190),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_186),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_211),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_175),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_36),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_182),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_42),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_195),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_46),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_184),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_206),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_54),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_65),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_152),
.Y(n_332)
);

INVx4_ASAP7_75t_R g333 ( 
.A(n_39),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_66),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_47),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_57),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_68),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_153),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_145),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_122),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_31),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_235),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_65),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_125),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_29),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_76),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_217),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_19),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_4),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_128),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_127),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_25),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_187),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_132),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_37),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_112),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_86),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_170),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_105),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_22),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_71),
.Y(n_361)
);

BUFx5_ASAP7_75t_L g362 ( 
.A(n_52),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_199),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_63),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_114),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_144),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_5),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_59),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_24),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_227),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_87),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_94),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_234),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_87),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_214),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_49),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_171),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_64),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_15),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_156),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_137),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_88),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_91),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_7),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_142),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_53),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_143),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_80),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_116),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_139),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_154),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_13),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_113),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_157),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_98),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_229),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_29),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_5),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_44),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_4),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_135),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_172),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_136),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_95),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_151),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_140),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_207),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_53),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_107),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_191),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_58),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_71),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_35),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_61),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_11),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_17),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_176),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_161),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_50),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_212),
.Y(n_420)
);

CKINVDCx11_ASAP7_75t_R g421 ( 
.A(n_213),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_165),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_76),
.Y(n_423)
);

BUFx5_ASAP7_75t_L g424 ( 
.A(n_40),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_68),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_7),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_129),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_83),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_45),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_100),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_81),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_69),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_51),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_9),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_150),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_49),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_20),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_28),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_2),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_230),
.Y(n_440)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_77),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_67),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_120),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_16),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_81),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_35),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_109),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_181),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_61),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_97),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_89),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_167),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_74),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_219),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_60),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_34),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_118),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_23),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_208),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_215),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_1),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_50),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_70),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_179),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_45),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_345),
.B(n_0),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_304),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_362),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_441),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_421),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_251),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_283),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_465),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_362),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_287),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_320),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_362),
.Y(n_479)
);

INVxp33_ASAP7_75t_SL g480 ( 
.A(n_240),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_362),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_351),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_447),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_274),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_362),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_362),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_362),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_313),
.B(n_0),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_362),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_386),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_424),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_284),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_290),
.Y(n_494)
);

BUFx2_ASAP7_75t_SL g495 ( 
.A(n_282),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_424),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_240),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_295),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_424),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_424),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_424),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_415),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_465),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_6),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_266),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_247),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_297),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_266),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_266),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_323),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_266),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_266),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_318),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_247),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_331),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_431),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_318),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_334),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_425),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_335),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_405),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_282),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_461),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_336),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_291),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_239),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_291),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_301),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_442),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_337),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_391),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_243),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_298),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_341),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_244),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_282),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_348),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_298),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_349),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_456),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_352),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_302),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_248),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_245),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_301),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_302),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_248),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_339),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_321),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_289),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_390),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_249),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_313),
.B(n_6),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_390),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_396),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_249),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_357),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_396),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_250),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_252),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_270),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_367),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_270),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_273),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_255),
.B(n_8),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_340),
.B(n_8),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_275),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_301),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_278),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_368),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_292),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_293),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_369),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_306),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_289),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_325),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_371),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_376),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_289),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_327),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_404),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_330),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_350),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_378),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_379),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_384),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_404),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_398),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_350),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_343),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_586),
.B(n_358),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_552),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_552),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_552),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_514),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_552),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_514),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_514),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_514),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_534),
.B(n_393),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_470),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_586),
.B(n_305),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_471),
.B(n_406),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_552),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_468),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_586),
.B(n_350),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_476),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_468),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_468),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_551),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_476),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_551),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_534),
.B(n_584),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_551),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_584),
.B(n_253),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_479),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_479),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_481),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_481),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_485),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_485),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_486),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_586),
.B(n_321),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_486),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_475),
.B(n_505),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_487),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_487),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_471),
.B(n_420),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_489),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_489),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_491),
.B(n_267),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_491),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_492),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_492),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_472),
.Y(n_639)
);

OA21x2_ASAP7_75t_L g640 ( 
.A1(n_496),
.A2(n_277),
.B(n_272),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_471),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_590),
.B(n_406),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_496),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_499),
.B(n_285),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_590),
.B(n_420),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_499),
.B(n_288),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_500),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_500),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_501),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_501),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_495),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_503),
.B(n_296),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_503),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_590),
.B(n_409),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_504),
.A2(n_309),
.B(n_307),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_504),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_507),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_507),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_510),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_528),
.B(n_409),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_569),
.B(n_305),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_510),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_511),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_511),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_513),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_528),
.A2(n_319),
.B(n_310),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_513),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_562),
.B(n_420),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_530),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_530),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_562),
.B(n_346),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_536),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_536),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_541),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_541),
.B(n_324),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_497),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_545),
.B(n_326),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_484),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_545),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_549),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_549),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_554),
.A2(n_359),
.B(n_344),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_554),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_557),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_557),
.B(n_370),
.Y(n_685)
);

XNOR2xp5_ASAP7_75t_L g686 ( 
.A(n_490),
.B(n_275),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_558),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_558),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_561),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_561),
.B(n_529),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_480),
.B(n_526),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_515),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_651),
.B(n_523),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_610),
.B(n_495),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_614),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_648),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_624),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_668),
.A2(n_568),
.B1(n_466),
.B2(n_556),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_605),
.B(n_523),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_SL g700 ( 
.A1(n_686),
.A2(n_518),
.B1(n_532),
.B2(n_502),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_627),
.B(n_339),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_678),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_614),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_661),
.A2(n_668),
.B1(n_594),
.B2(n_606),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_651),
.B(n_493),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_624),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_605),
.B(n_525),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_610),
.B(n_535),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_605),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_691),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_691),
.B(n_494),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_614),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_676),
.B(n_525),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_624),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_678),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_618),
.Y(n_716)
);

AND2x6_ASAP7_75t_L g717 ( 
.A(n_668),
.B(n_321),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_627),
.B(n_339),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_625),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_606),
.B(n_498),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_612),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_612),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_648),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_661),
.B(n_539),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_639),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_639),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_625),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_610),
.B(n_509),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_639),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_594),
.B(n_512),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_625),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_660),
.A2(n_466),
.B1(n_488),
.B2(n_506),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_629),
.B(n_517),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_612),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_648),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_618),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_613),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_627),
.B(n_339),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_634),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_648),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_641),
.B(n_539),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_611),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_613),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_632),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_613),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_616),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_648),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_629),
.B(n_520),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_618),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_611),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_618),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_616),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_641),
.B(n_522),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_616),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_660),
.A2(n_506),
.B1(n_516),
.B2(n_508),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_616),
.Y(n_756)
);

BUFx6f_ASAP7_75t_SL g757 ( 
.A(n_607),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_634),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_676),
.B(n_546),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_632),
.B(n_527),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_641),
.B(n_533),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_615),
.Y(n_762)
);

INVx5_ASAP7_75t_L g763 ( 
.A(n_627),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_660),
.A2(n_555),
.B1(n_559),
.B2(n_550),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_627),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_617),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_686),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_SL g768 ( 
.A(n_632),
.B(n_467),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_616),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_645),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_629),
.B(n_537),
.Y(n_771)
);

INVx8_ASAP7_75t_L g772 ( 
.A(n_627),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_645),
.B(n_540),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_634),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_609),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_609),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_686),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_609),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_645),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_618),
.Y(n_780)
);

INVx5_ASAP7_75t_L g781 ( 
.A(n_627),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_607),
.A2(n_542),
.B1(n_560),
.B2(n_544),
.Y(n_782)
);

BUFx6f_ASAP7_75t_SL g783 ( 
.A(n_607),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_627),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_607),
.B(n_565),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_643),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_609),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_SL g788 ( 
.A1(n_690),
.A2(n_548),
.B1(n_571),
.B2(n_531),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_607),
.B(n_573),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_642),
.B(n_576),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_609),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_643),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_671),
.B(n_692),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_690),
.A2(n_241),
.B1(n_355),
.B2(n_315),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_618),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_643),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_647),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_654),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_647),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_647),
.Y(n_800)
);

BUFx10_ASAP7_75t_L g801 ( 
.A(n_642),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_649),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_649),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_627),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_649),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_642),
.B(n_580),
.Y(n_806)
);

BUFx4f_ASAP7_75t_L g807 ( 
.A(n_627),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_601),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_642),
.B(n_581),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_604),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_601),
.Y(n_811)
);

BUFx10_ASAP7_75t_L g812 ( 
.A(n_642),
.Y(n_812)
);

BUFx6f_ASAP7_75t_SL g813 ( 
.A(n_654),
.Y(n_813)
);

BUFx10_ASAP7_75t_L g814 ( 
.A(n_654),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_601),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_671),
.B(n_538),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_654),
.B(n_587),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_671),
.B(n_547),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_604),
.B(n_564),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_598),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_601),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_641),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_641),
.B(n_588),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_617),
.B(n_654),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_692),
.B(n_563),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_SL g826 ( 
.A(n_660),
.B(n_553),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_598),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_619),
.B(n_566),
.Y(n_828)
);

BUFx10_ASAP7_75t_L g829 ( 
.A(n_660),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_601),
.Y(n_830)
);

AND2x6_ASAP7_75t_L g831 ( 
.A(n_618),
.B(n_321),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_602),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_653),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_653),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_635),
.B(n_589),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_653),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_653),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_653),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_602),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_603),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_628),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_628),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_615),
.B(n_591),
.C(n_570),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_635),
.B(n_473),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_620),
.B(n_593),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_603),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_644),
.B(n_478),
.Y(n_847)
);

OAI22xp33_ASAP7_75t_L g848 ( 
.A1(n_675),
.A2(n_280),
.B1(n_281),
.B2(n_276),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_640),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_628),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_644),
.A2(n_437),
.B1(n_444),
.B2(n_436),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_646),
.B(n_242),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_628),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_628),
.Y(n_854)
);

NAND2xp33_ASAP7_75t_L g855 ( 
.A(n_628),
.B(n_339),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_619),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_695),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_704),
.B(n_620),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_810),
.B(n_621),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_710),
.B(n_694),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_856),
.B(n_621),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_856),
.B(n_622),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_820),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_L g864 ( 
.A(n_724),
.B(n_688),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_708),
.B(n_622),
.Y(n_865)
);

NOR2xp67_ASAP7_75t_L g866 ( 
.A(n_707),
.B(n_688),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_708),
.B(n_623),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_708),
.B(n_623),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_766),
.B(n_626),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_744),
.B(n_626),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_726),
.B(n_578),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_720),
.B(n_630),
.Y(n_872)
);

INVx8_ASAP7_75t_L g873 ( 
.A(n_772),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_696),
.B(n_723),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_827),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_827),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_832),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_744),
.B(n_630),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_760),
.B(n_633),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_773),
.B(n_633),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_725),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_715),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_725),
.B(n_582),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_759),
.B(n_474),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_699),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_770),
.B(n_779),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_698),
.A2(n_640),
.B1(n_592),
.B2(n_669),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_709),
.B(n_469),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_816),
.B(n_477),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_770),
.B(n_669),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_702),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_696),
.B(n_723),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_SL g893 ( 
.A(n_699),
.B(n_482),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_832),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_779),
.B(n_638),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_839),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_730),
.B(n_638),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_703),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_772),
.B(n_628),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_839),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_840),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_713),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_712),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_840),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_733),
.B(n_650),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_712),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_721),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_713),
.B(n_688),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_721),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_717),
.B(n_656),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_717),
.B(n_741),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_722),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_782),
.B(n_652),
.C(n_646),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_696),
.B(n_656),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_717),
.B(n_688),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_717),
.B(n_688),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_846),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_793),
.B(n_672),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_711),
.B(n_361),
.C(n_360),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_723),
.B(n_735),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_717),
.A2(n_652),
.B1(n_402),
.B2(n_672),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_793),
.B(n_845),
.Y(n_922)
);

NOR3xp33_ASAP7_75t_L g923 ( 
.A(n_729),
.B(n_374),
.C(n_364),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_753),
.B(n_673),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_798),
.A2(n_674),
.B1(n_679),
.B2(n_673),
.Y(n_925)
);

AOI221xp5_ASAP7_75t_L g926 ( 
.A1(n_794),
.A2(n_281),
.B1(n_280),
.B2(n_276),
.C(n_408),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_814),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_735),
.B(n_628),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_722),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_846),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_835),
.A2(n_392),
.B(n_397),
.C(n_388),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_742),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_735),
.B(n_631),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_748),
.B(n_631),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_761),
.B(n_674),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_734),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_734),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_771),
.B(n_631),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_728),
.B(n_631),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_737),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_742),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_825),
.B(n_816),
.Y(n_942)
);

NAND2xp33_ASAP7_75t_L g943 ( 
.A(n_772),
.B(n_631),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_825),
.B(n_679),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_818),
.B(n_681),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_818),
.B(n_681),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_SL g947 ( 
.A(n_826),
.B(n_483),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_750),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_819),
.B(n_543),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_750),
.B(n_684),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_762),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_798),
.A2(n_687),
.B1(n_684),
.B2(n_242),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_762),
.B(n_687),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_808),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_828),
.B(n_670),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_819),
.B(n_567),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_808),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_844),
.B(n_631),
.Y(n_958)
);

AND2x6_ASAP7_75t_L g959 ( 
.A(n_740),
.B(n_670),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_759),
.B(n_729),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_828),
.B(n_670),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_847),
.B(n_631),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_811),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_740),
.B(n_631),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_768),
.B(n_567),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_740),
.B(n_636),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_823),
.A2(n_637),
.B(n_636),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_811),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_R g969 ( 
.A(n_772),
.B(n_408),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_815),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_747),
.B(n_829),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_747),
.B(n_680),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_747),
.B(n_829),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_777),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_716),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_789),
.B(n_680),
.Y(n_976)
);

NAND2xp33_ASAP7_75t_L g977 ( 
.A(n_833),
.B(n_636),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_829),
.B(n_636),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_790),
.B(n_680),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_824),
.B(n_572),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_806),
.B(n_689),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_737),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_809),
.B(n_689),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_785),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_732),
.B(n_689),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_693),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_815),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_767),
.B(n_685),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_814),
.B(n_636),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_746),
.B(n_675),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_700),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_821),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_743),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_746),
.B(n_677),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_821),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_743),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_705),
.B(n_636),
.Y(n_997)
);

AND2x6_ASAP7_75t_L g998 ( 
.A(n_833),
.B(n_636),
.Y(n_998)
);

AND2x6_ASAP7_75t_SL g999 ( 
.A(n_767),
.B(n_399),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_814),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_745),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_807),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_824),
.A2(n_640),
.B1(n_683),
.B2(n_677),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_788),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_752),
.B(n_685),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_848),
.A2(n_411),
.B(n_423),
.C(n_400),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_824),
.B(n_817),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_851),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_745),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_792),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_752),
.B(n_636),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_754),
.B(n_637),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_754),
.B(n_637),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_852),
.B(n_637),
.Y(n_1014)
);

AND2x2_ASAP7_75t_SL g1015 ( 
.A(n_701),
.B(n_640),
.Y(n_1015)
);

NAND3x1_ASAP7_75t_L g1016 ( 
.A(n_764),
.B(n_428),
.C(n_426),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_765),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_813),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_843),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_756),
.B(n_637),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_792),
.Y(n_1021)
);

AO221x1_ASAP7_75t_L g1022 ( 
.A1(n_697),
.A2(n_453),
.B1(n_438),
.B2(n_455),
.C(n_458),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_756),
.B(n_637),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_769),
.B(n_637),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_860),
.B(n_755),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_863),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_860),
.A2(n_783),
.B1(n_757),
.B2(n_824),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_874),
.A2(n_836),
.B(n_834),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_873),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_1008),
.B(n_757),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_942),
.B(n_757),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_879),
.B(n_801),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_875),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_988),
.B(n_783),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_869),
.A2(n_967),
.B(n_935),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_922),
.A2(n_834),
.B(n_837),
.C(n_836),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_873),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_965),
.Y(n_1038)
);

INVxp33_ASAP7_75t_SL g1039 ( 
.A(n_882),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_858),
.A2(n_706),
.B(n_697),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_891),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_857),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_887),
.A2(n_783),
.B1(n_714),
.B2(n_719),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_879),
.B(n_801),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_880),
.B(n_801),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_SL g1046 ( 
.A1(n_947),
.A2(n_432),
.B1(n_813),
.B2(n_412),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_880),
.B(n_812),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_859),
.B(n_812),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_861),
.B(n_812),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_862),
.B(n_945),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_924),
.A2(n_838),
.B(n_837),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_946),
.B(n_706),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_874),
.A2(n_838),
.B(n_841),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_918),
.B(n_714),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_1017),
.B(n_716),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_892),
.A2(n_842),
.B(n_841),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_918),
.B(n_719),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_881),
.B(n_830),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_866),
.A2(n_813),
.B1(n_830),
.B2(n_731),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_1006),
.A2(n_775),
.B(n_776),
.C(n_769),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_892),
.A2(n_731),
.B(n_727),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_920),
.A2(n_739),
.B(n_727),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_873),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1019),
.B(n_850),
.Y(n_1064)
);

INVx11_ASAP7_75t_L g1065 ( 
.A(n_959),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_898),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_1017),
.B(n_716),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_920),
.A2(n_758),
.B(n_739),
.Y(n_1068)
);

NOR2xp67_ASAP7_75t_L g1069 ( 
.A(n_871),
.B(n_775),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_928),
.A2(n_842),
.B(n_850),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_913),
.A2(n_774),
.B(n_786),
.C(n_758),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_928),
.A2(n_853),
.B(n_850),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_898),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_986),
.B(n_853),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_925),
.A2(n_822),
.B1(n_849),
.B2(n_853),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_933),
.A2(n_854),
.B(n_822),
.Y(n_1076)
);

OR2x2_ASAP7_75t_SL g1077 ( 
.A(n_884),
.B(n_462),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_872),
.A2(n_786),
.B(n_799),
.C(n_774),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_918),
.B(n_799),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_956),
.B(n_800),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_885),
.B(n_854),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_889),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_960),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_933),
.A2(n_854),
.B(n_822),
.Y(n_1084)
);

BUFx4f_ASAP7_75t_L g1085 ( 
.A(n_1007),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_1017),
.B(n_716),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_902),
.B(n_897),
.Y(n_1087)
);

NOR3xp33_ASAP7_75t_L g1088 ( 
.A(n_926),
.B(n_883),
.C(n_923),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_964),
.A2(n_849),
.B(n_803),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_964),
.A2(n_803),
.B(n_800),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_903),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_890),
.B(n_776),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_858),
.A2(n_797),
.B(n_802),
.C(n_796),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_890),
.B(n_778),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_903),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_890),
.B(n_778),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_966),
.A2(n_791),
.B(n_787),
.Y(n_1097)
);

OAI321xp33_ASAP7_75t_L g1098 ( 
.A1(n_949),
.A2(n_577),
.A3(n_572),
.B1(n_574),
.B2(n_575),
.C(n_579),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_893),
.B(n_574),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_886),
.A2(n_878),
.B(n_895),
.C(n_870),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_955),
.B(n_787),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_975),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_974),
.B(n_791),
.Y(n_1103)
);

NAND2x1p5_ASAP7_75t_L g1104 ( 
.A(n_1002),
.B(n_765),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_961),
.B(n_865),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_966),
.A2(n_736),
.B(n_716),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_972),
.A2(n_749),
.B(n_736),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_876),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_867),
.B(n_796),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_975),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_868),
.B(n_797),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_908),
.B(n_575),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1011),
.A2(n_749),
.B(n_736),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_1002),
.B(n_765),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_927),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_888),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_877),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1012),
.A2(n_749),
.B(n_736),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1013),
.A2(n_749),
.B(n_736),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_944),
.B(n_802),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_914),
.A2(n_805),
.B(n_655),
.Y(n_1121)
);

OAI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_872),
.A2(n_413),
.B(n_412),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_991),
.B(n_577),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1020),
.A2(n_751),
.B(n_749),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_905),
.B(n_805),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1023),
.A2(n_780),
.B(n_751),
.Y(n_1126)
);

AOI33xp33_ASAP7_75t_L g1127 ( 
.A1(n_894),
.A2(n_583),
.A3(n_579),
.B1(n_585),
.B2(n_521),
.B3(n_524),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1024),
.A2(n_780),
.B(n_751),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_905),
.B(n_980),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_897),
.B(n_751),
.Y(n_1130)
);

NAND2xp33_ASAP7_75t_L g1131 ( 
.A(n_959),
.B(n_751),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_914),
.A2(n_855),
.B(n_585),
.C(n_583),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_980),
.B(n_780),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1014),
.A2(n_655),
.B(n_666),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_L g1135 ( 
.A(n_959),
.B(n_780),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_975),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1007),
.A2(n_784),
.B1(n_804),
.B2(n_855),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1014),
.A2(n_655),
.B(n_666),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_954),
.A2(n_682),
.B(n_666),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1007),
.B(n_780),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_980),
.B(n_515),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_990),
.A2(n_795),
.B(n_807),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1004),
.B(n_519),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1003),
.A2(n_907),
.B(n_906),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_934),
.A2(n_807),
.B(n_682),
.C(n_718),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1018),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_984),
.B(n_795),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_864),
.B(n_795),
.Y(n_1148)
);

AND2x2_ASAP7_75t_SL g1149 ( 
.A(n_1015),
.B(n_701),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_927),
.B(n_784),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_932),
.B(n_795),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_976),
.B(n_795),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_994),
.A2(n_738),
.B(n_718),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_934),
.A2(n_682),
.B(n_738),
.C(n_377),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_950),
.A2(n_667),
.B(n_665),
.C(n_663),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1000),
.B(n_784),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_938),
.B(n_804),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_957),
.A2(n_804),
.B(n_640),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_979),
.B(n_981),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_963),
.A2(n_659),
.B(n_657),
.Y(n_1160)
);

NOR2xp67_ASAP7_75t_L g1161 ( 
.A(n_952),
.B(n_683),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_SL g1162 ( 
.A(n_1000),
.B(n_763),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_941),
.B(n_637),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1005),
.A2(n_781),
.B(n_763),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_983),
.B(n_948),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_959),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_L g1167 ( 
.A(n_938),
.B(n_683),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_968),
.A2(n_659),
.B(n_657),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_975),
.B(n_763),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_970),
.A2(n_992),
.B(n_987),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_951),
.B(n_683),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_906),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_971),
.A2(n_781),
.B(n_763),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_896),
.A2(n_429),
.B1(n_463),
.B2(n_419),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_900),
.B(n_683),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_901),
.B(n_683),
.Y(n_1176)
);

AOI21xp33_ASAP7_75t_L g1177 ( 
.A1(n_985),
.A2(n_414),
.B(n_413),
.Y(n_1177)
);

NOR2x1p5_ASAP7_75t_L g1178 ( 
.A(n_953),
.B(n_414),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_904),
.B(n_683),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_911),
.A2(n_665),
.B(n_663),
.Y(n_1180)
);

INVx11_ASAP7_75t_L g1181 ( 
.A(n_959),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_973),
.B(n_917),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_939),
.A2(n_419),
.B(n_416),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_973),
.A2(n_781),
.B(n_596),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_978),
.A2(n_781),
.B(n_596),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_930),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_958),
.B(n_416),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_939),
.A2(n_433),
.B1(n_463),
.B2(n_434),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_999),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_978),
.A2(n_596),
.B(n_595),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_958),
.B(n_429),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_998),
.Y(n_1192)
);

AND2x4_ASAP7_75t_SL g1193 ( 
.A(n_919),
.B(n_432),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_962),
.B(n_433),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_995),
.B(n_1010),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_962),
.B(n_434),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_997),
.B(n_667),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_998),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1016),
.B(n_519),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1010),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_989),
.A2(n_597),
.B(n_595),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_989),
.A2(n_597),
.B(n_595),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1021),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_998),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_977),
.A2(n_600),
.B(n_597),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_997),
.B(n_445),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_R g1207 ( 
.A(n_899),
.B(n_246),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_977),
.A2(n_608),
.B(n_600),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1022),
.B(n_521),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1021),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1032),
.A2(n_943),
.B(n_899),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_1041),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1026),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1044),
.A2(n_943),
.B(n_1015),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1087),
.A2(n_931),
.B(n_921),
.C(n_910),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1088),
.A2(n_916),
.B1(n_915),
.B2(n_998),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1123),
.B(n_432),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1083),
.B(n_524),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1050),
.B(n_1009),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1025),
.B(n_1009),
.Y(n_1220)
);

INVx4_ASAP7_75t_L g1221 ( 
.A(n_1029),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1029),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1045),
.A2(n_909),
.B(n_907),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1029),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1047),
.A2(n_912),
.B(n_909),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1082),
.Y(n_1226)
);

OAI21xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1149),
.A2(n_929),
.B(n_912),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1033),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1042),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1159),
.A2(n_936),
.B(n_929),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1087),
.B(n_969),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_SL g1232 ( 
.A(n_1116),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1035),
.A2(n_937),
.B(n_936),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1039),
.B(n_937),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1108),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1129),
.B(n_1030),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1088),
.A2(n_454),
.B(n_394),
.C(n_403),
.Y(n_1237)
);

CKINVDCx16_ASAP7_75t_R g1238 ( 
.A(n_1146),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1141),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1152),
.A2(n_982),
.B(n_940),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1143),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1085),
.B(n_940),
.Y(n_1242)
);

AND2x2_ASAP7_75t_SL g1243 ( 
.A(n_1085),
.B(n_969),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1105),
.B(n_982),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1131),
.A2(n_1135),
.B(n_1052),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1038),
.B(n_1030),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_L g1247 ( 
.A(n_1183),
.B(n_449),
.C(n_446),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1099),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1077),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1038),
.B(n_1001),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1029),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1117),
.Y(n_1252)
);

AOI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1180),
.A2(n_996),
.B(n_993),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1199),
.A2(n_996),
.B1(n_993),
.B2(n_1001),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1182),
.A2(n_372),
.B(n_381),
.C(n_451),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1186),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_1178),
.Y(n_1257)
);

NOR3xp33_ASAP7_75t_SL g1258 ( 
.A(n_1174),
.B(n_254),
.C(n_246),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1080),
.A2(n_382),
.B1(n_389),
.B2(n_407),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1031),
.B(n_998),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1122),
.A2(n_1188),
.B(n_1177),
.C(n_1100),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1130),
.A2(n_608),
.B(n_600),
.Y(n_1262)
);

BUFx4f_ASAP7_75t_L g1263 ( 
.A(n_1037),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1031),
.B(n_254),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1182),
.A2(n_440),
.B(n_430),
.C(n_662),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1034),
.A2(n_1140),
.B1(n_1081),
.B2(n_1069),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1195),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1199),
.A2(n_333),
.B1(n_256),
.B2(n_257),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1130),
.A2(n_608),
.B(n_286),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1127),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1113),
.A2(n_294),
.B(n_238),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1054),
.A2(n_662),
.B1(n_279),
.B2(n_271),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1037),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1112),
.B(n_256),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1034),
.B(n_257),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1103),
.B(n_662),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1120),
.B(n_831),
.Y(n_1277)
);

AO32x1_ASAP7_75t_L g1278 ( 
.A1(n_1209),
.A2(n_831),
.A3(n_664),
.B1(n_658),
.B2(n_13),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1199),
.B(n_10),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1193),
.B(n_10),
.Y(n_1280)
);

OAI22x1_ASAP7_75t_L g1281 ( 
.A1(n_1027),
.A2(n_258),
.B1(n_427),
.B2(n_459),
.Y(n_1281)
);

AOI21xp33_ASAP7_75t_L g1282 ( 
.A1(n_1043),
.A2(n_664),
.B(n_658),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1118),
.A2(n_1124),
.B(n_1119),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1098),
.B(n_258),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1048),
.B(n_1049),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1165),
.B(n_831),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1078),
.A2(n_831),
.B(n_260),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1058),
.Y(n_1288)
);

AND2x2_ASAP7_75t_SL g1289 ( 
.A(n_1149),
.B(n_321),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1065),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1125),
.B(n_1057),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1064),
.A2(n_354),
.B(n_260),
.C(n_261),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1078),
.A2(n_831),
.B(n_261),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1043),
.A2(n_831),
.B1(n_259),
.B2(n_354),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1204),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1079),
.A2(n_259),
.B1(n_262),
.B2(n_464),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1200),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1064),
.A2(n_262),
.B(n_263),
.C(n_264),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1101),
.B(n_658),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1126),
.A2(n_300),
.B(n_299),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1210),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1046),
.B(n_11),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1147),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1128),
.A2(n_366),
.B(n_303),
.Y(n_1304)
);

BUFx8_ASAP7_75t_L g1305 ( 
.A(n_1037),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1046),
.B(n_263),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1081),
.B(n_264),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1074),
.A2(n_265),
.B(n_268),
.C(n_269),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_1204),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1147),
.Y(n_1310)
);

OAI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1187),
.A2(n_265),
.B1(n_268),
.B2(n_464),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1204),
.B(n_658),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1140),
.B(n_658),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1107),
.A2(n_375),
.B(n_308),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1066),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1109),
.B(n_658),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1073),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1191),
.B(n_658),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1091),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1203),
.A2(n_1172),
.B1(n_1095),
.B2(n_1194),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1153),
.A2(n_380),
.B(n_311),
.Y(n_1321)
);

AOI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1040),
.A2(n_664),
.B(n_658),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1037),
.B(n_664),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1092),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1142),
.A2(n_383),
.B(n_312),
.Y(n_1325)
);

AO32x1_ASAP7_75t_L g1326 ( 
.A1(n_1075),
.A2(n_664),
.A3(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_1326)
);

NAND2x1p5_ASAP7_75t_L g1327 ( 
.A(n_1063),
.B(n_664),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1074),
.A2(n_269),
.B(n_271),
.C(n_460),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1181),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1051),
.A2(n_387),
.B(n_314),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1144),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_SL g1332 ( 
.A1(n_1115),
.A2(n_12),
.B(n_14),
.C(n_18),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1161),
.A2(n_1196),
.B(n_1036),
.C(n_1206),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1094),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1096),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1071),
.A2(n_12),
.B(n_20),
.C(n_21),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1111),
.A2(n_279),
.B1(n_410),
.B2(n_460),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1133),
.B(n_664),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1115),
.B(n_1151),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1063),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1063),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1150),
.B(n_1071),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1171),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1063),
.B(n_410),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1150),
.B(n_664),
.Y(n_1345)
);

AOI22x1_ASAP7_75t_L g1346 ( 
.A1(n_1076),
.A2(n_417),
.B1(n_459),
.B2(n_418),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1204),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1132),
.A2(n_21),
.B(n_24),
.C(n_25),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1175),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1102),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_SL g1351 ( 
.A(n_1104),
.B(n_1114),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1176),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1134),
.A2(n_373),
.B(n_457),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1189),
.B(n_1170),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1102),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1138),
.A2(n_365),
.B(n_452),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1145),
.A2(n_1060),
.B(n_1163),
.C(n_1151),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1207),
.B(n_417),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_SL g1359 ( 
.A(n_1104),
.B(n_418),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1160),
.B(n_26),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1056),
.A2(n_1106),
.B(n_1089),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1157),
.A2(n_422),
.B1(n_427),
.B2(n_448),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1197),
.B(n_422),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1179),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1061),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1207),
.B(n_316),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1062),
.B(n_339),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1102),
.B(n_1110),
.Y(n_1368)
);

BUFx5_ASAP7_75t_L g1369 ( 
.A(n_1114),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1102),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1110),
.B(n_26),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1068),
.B(n_339),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1245),
.A2(n_1067),
.B(n_1086),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1237),
.A2(n_1059),
.B(n_1155),
.C(n_1167),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1233),
.A2(n_1283),
.B(n_1361),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1211),
.A2(n_1055),
.B(n_1067),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1322),
.A2(n_1139),
.B(n_1053),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1212),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1213),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1261),
.A2(n_1163),
.B(n_1137),
.C(n_1154),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1253),
.A2(n_1331),
.B(n_1240),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1307),
.A2(n_1070),
.B(n_1084),
.Y(n_1382)
);

OAI22x1_ASAP7_75t_L g1383 ( 
.A1(n_1306),
.A2(n_1166),
.B1(n_1055),
.B2(n_1086),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1231),
.A2(n_1072),
.B(n_1090),
.Y(n_1384)
);

AO31x2_ASAP7_75t_L g1385 ( 
.A1(n_1357),
.A2(n_1333),
.A3(n_1220),
.B(n_1214),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1226),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1223),
.A2(n_1121),
.B(n_1097),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1241),
.A2(n_1166),
.B1(n_1192),
.B2(n_1198),
.Y(n_1388)
);

AOI221xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1336),
.A2(n_1028),
.B1(n_1168),
.B2(n_1202),
.C(n_1201),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1230),
.A2(n_1148),
.A3(n_1190),
.B(n_1205),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1262),
.A2(n_1208),
.B(n_1184),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1239),
.B(n_1267),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1219),
.A2(n_1093),
.B(n_1156),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1236),
.B(n_1110),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1264),
.A2(n_1156),
.B(n_1185),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1225),
.A2(n_1158),
.B(n_1198),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1289),
.A2(n_1192),
.B1(n_1162),
.B2(n_1093),
.Y(n_1397)
);

BUFx2_ASAP7_75t_R g1398 ( 
.A(n_1249),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1367),
.A2(n_1164),
.B(n_1173),
.Y(n_1399)
);

AO22x1_ASAP7_75t_L g1400 ( 
.A1(n_1302),
.A2(n_1279),
.B1(n_1354),
.B2(n_1280),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1295),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1219),
.A2(n_1136),
.B(n_1110),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1291),
.A2(n_1342),
.B(n_1285),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1266),
.B(n_1136),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1291),
.A2(n_1342),
.B(n_1244),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1263),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1238),
.Y(n_1407)
);

AO31x2_ASAP7_75t_L g1408 ( 
.A1(n_1372),
.A2(n_1169),
.A3(n_1136),
.B(n_339),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1234),
.B(n_27),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1299),
.A2(n_338),
.B(n_599),
.Y(n_1410)
);

NOR2x1_ASAP7_75t_R g1411 ( 
.A(n_1347),
.B(n_317),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1305),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1287),
.A2(n_356),
.B(n_450),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1292),
.A2(n_322),
.B(n_328),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1228),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1235),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1305),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1248),
.B(n_28),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1348),
.B(n_1255),
.C(n_1360),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1299),
.A2(n_338),
.B(n_599),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1260),
.A2(n_338),
.B(n_599),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1339),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1263),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1316),
.A2(n_338),
.B(n_599),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1312),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1218),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1217),
.B(n_30),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1363),
.A2(n_329),
.B1(n_332),
.B2(n_443),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1316),
.A2(n_338),
.B(n_599),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1312),
.A2(n_385),
.B(n_435),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1365),
.A2(n_1351),
.B(n_1353),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1284),
.A2(n_401),
.B(n_395),
.C(n_363),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1351),
.A2(n_599),
.B(n_353),
.Y(n_1433)
);

AO32x2_ASAP7_75t_L g1434 ( 
.A1(n_1259),
.A2(n_1272),
.A3(n_1296),
.B1(n_1326),
.B2(n_1227),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1341),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1372),
.A2(n_599),
.B(n_185),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1246),
.B(n_30),
.Y(n_1437)
);

CKINVDCx11_ASAP7_75t_R g1438 ( 
.A(n_1222),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1356),
.A2(n_599),
.B(n_347),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1312),
.A2(n_342),
.B(n_236),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1287),
.A2(n_231),
.B(n_226),
.Y(n_1441)
);

NOR2xp67_ASAP7_75t_L g1442 ( 
.A(n_1368),
.B(n_222),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1222),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1293),
.A2(n_210),
.B(n_203),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1252),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1258),
.B(n_31),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1298),
.A2(n_32),
.B(n_33),
.Y(n_1447)
);

CKINVDCx8_ASAP7_75t_R g1448 ( 
.A(n_1222),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1270),
.B(n_32),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1256),
.B(n_1275),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1259),
.A2(n_1243),
.B1(n_1359),
.B2(n_1281),
.Y(n_1451)
);

O2A1O1Ixp5_ASAP7_75t_L g1452 ( 
.A1(n_1293),
.A2(n_33),
.B(n_34),
.C(n_36),
.Y(n_1452)
);

AO31x2_ASAP7_75t_L g1453 ( 
.A1(n_1343),
.A2(n_201),
.A3(n_197),
.B(n_196),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1277),
.A2(n_194),
.B(n_193),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1277),
.A2(n_189),
.B(n_183),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1313),
.A2(n_178),
.B(n_169),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1290),
.B(n_163),
.Y(n_1457)
);

AOI221x1_ASAP7_75t_L g1458 ( 
.A1(n_1265),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.C(n_44),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1313),
.A2(n_160),
.B(n_159),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1297),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1301),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1363),
.A2(n_46),
.B1(n_48),
.B2(n_52),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1257),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1315),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1286),
.A2(n_141),
.B(n_134),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1359),
.A2(n_48),
.B1(n_54),
.B2(n_55),
.Y(n_1466)
);

AO32x2_ASAP7_75t_L g1467 ( 
.A1(n_1272),
.A2(n_55),
.A3(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1224),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1296),
.B(n_60),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1282),
.A2(n_1286),
.B(n_1269),
.Y(n_1470)
);

O2A1O1Ixp5_ASAP7_75t_SL g1471 ( 
.A1(n_1303),
.A2(n_62),
.B(n_67),
.C(n_70),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_R g1472 ( 
.A(n_1232),
.B(n_121),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1319),
.Y(n_1473)
);

A2O1A1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1247),
.A2(n_62),
.B(n_72),
.C(n_73),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1232),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1349),
.A2(n_117),
.B(n_115),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1268),
.B(n_72),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1352),
.A2(n_111),
.B(n_103),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1250),
.B(n_73),
.Y(n_1479)
);

AO31x2_ASAP7_75t_L g1480 ( 
.A1(n_1364),
.A2(n_96),
.A3(n_93),
.B(n_79),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1311),
.A2(n_74),
.B(n_77),
.C(n_80),
.Y(n_1481)
);

BUFx8_ASAP7_75t_L g1482 ( 
.A(n_1329),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1310),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_1483)
);

INVx8_ASAP7_75t_L g1484 ( 
.A(n_1224),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1324),
.B(n_82),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1334),
.B(n_84),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1274),
.B(n_85),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1224),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1345),
.A2(n_85),
.B(n_86),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1314),
.A2(n_1304),
.B(n_1300),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1345),
.A2(n_1309),
.B(n_1215),
.Y(n_1491)
);

NOR2xp67_ASAP7_75t_L g1492 ( 
.A(n_1370),
.B(n_1221),
.Y(n_1492)
);

CKINVDCx11_ASAP7_75t_R g1493 ( 
.A(n_1251),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1335),
.B(n_1288),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1337),
.B(n_1317),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1358),
.B(n_1366),
.Y(n_1496)
);

BUFx10_ASAP7_75t_L g1497 ( 
.A(n_1251),
.Y(n_1497)
);

OAI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1362),
.A2(n_1216),
.B1(n_1371),
.B2(n_1242),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1318),
.A2(n_1321),
.B(n_1326),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1355),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1276),
.B(n_1350),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1221),
.B(n_1340),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1308),
.A2(n_1328),
.B(n_1330),
.Y(n_1503)
);

OAI21xp33_ASAP7_75t_L g1504 ( 
.A1(n_1346),
.A2(n_1294),
.B(n_1344),
.Y(n_1504)
);

A2O1A1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1254),
.A2(n_1325),
.B(n_1320),
.C(n_1271),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1251),
.Y(n_1506)
);

BUFx12f_ASAP7_75t_L g1507 ( 
.A(n_1273),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1276),
.B(n_1273),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1338),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1326),
.A2(n_1278),
.B(n_1327),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1273),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_1340),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1340),
.B(n_1323),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1278),
.A2(n_1327),
.B(n_1332),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1242),
.A2(n_1369),
.B(n_1282),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1369),
.B(n_1278),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1369),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1369),
.A2(n_1233),
.B(n_1283),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1369),
.B(n_710),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1236),
.B(n_710),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1233),
.A2(n_1283),
.B(n_1361),
.Y(n_1521)
);

AO31x2_ASAP7_75t_L g1522 ( 
.A1(n_1331),
.A2(n_1357),
.A3(n_1283),
.B(n_1333),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1237),
.A2(n_1261),
.B(n_1236),
.C(n_880),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1289),
.A2(n_1088),
.B1(n_1236),
.B2(n_960),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1212),
.Y(n_1525)
);

O2A1O1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1237),
.A2(n_710),
.B(n_730),
.C(n_720),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1289),
.A2(n_1088),
.B1(n_1236),
.B2(n_960),
.Y(n_1527)
);

A2O1A1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1237),
.A2(n_1261),
.B(n_1236),
.C(n_880),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_SL g1529 ( 
.A(n_1289),
.B(n_1243),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1236),
.B(n_710),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1213),
.Y(n_1531)
);

INVx5_ASAP7_75t_L g1532 ( 
.A(n_1312),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1307),
.A2(n_1044),
.B(n_1032),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1236),
.B(n_710),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1237),
.A2(n_1261),
.B(n_1236),
.C(n_880),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1245),
.A2(n_1211),
.B(n_1135),
.Y(n_1536)
);

AO31x2_ASAP7_75t_L g1537 ( 
.A1(n_1331),
.A2(n_1357),
.A3(n_1283),
.B(n_1333),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1213),
.Y(n_1538)
);

INVx3_ASAP7_75t_SL g1539 ( 
.A(n_1238),
.Y(n_1539)
);

BUFx4_ASAP7_75t_SL g1540 ( 
.A(n_1212),
.Y(n_1540)
);

OAI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1307),
.A2(n_1044),
.B(n_1032),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1307),
.A2(n_1044),
.B(n_1032),
.Y(n_1542)
);

AOI221xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1336),
.A2(n_1348),
.B1(n_1261),
.B2(n_1237),
.C(n_698),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1213),
.Y(n_1544)
);

AOI221x1_ASAP7_75t_L g1545 ( 
.A1(n_1255),
.A2(n_1281),
.B1(n_1306),
.B2(n_1236),
.C(n_1259),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1236),
.B(n_710),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1229),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1212),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1524),
.A2(n_1527),
.B1(n_1419),
.B2(n_1469),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_SL g1550 ( 
.A1(n_1529),
.A2(n_1413),
.B1(n_1419),
.B2(n_1477),
.Y(n_1550)
);

CKINVDCx6p67_ASAP7_75t_R g1551 ( 
.A(n_1539),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_1530),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1426),
.B(n_1422),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1524),
.A2(n_1527),
.B1(n_1413),
.B2(n_1451),
.Y(n_1554)
);

BUFx12f_ASAP7_75t_L g1555 ( 
.A(n_1438),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1445),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1529),
.A2(n_1447),
.B1(n_1462),
.B2(n_1409),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1451),
.A2(n_1483),
.B1(n_1466),
.B2(n_1450),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1379),
.Y(n_1559)
);

OAI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1466),
.A2(n_1483),
.B1(n_1545),
.B2(n_1546),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1487),
.A2(n_1533),
.B1(n_1542),
.B2(n_1541),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1534),
.B(n_1392),
.Y(n_1562)
);

BUFx12f_ASAP7_75t_L g1563 ( 
.A(n_1493),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1543),
.A2(n_1523),
.B1(n_1535),
.B2(n_1528),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1532),
.B(n_1423),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1417),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1532),
.Y(n_1567)
);

BUFx2_ASAP7_75t_SL g1568 ( 
.A(n_1512),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_SL g1569 ( 
.A1(n_1481),
.A2(n_1458),
.B(n_1526),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1504),
.A2(n_1437),
.B1(n_1446),
.B2(n_1449),
.Y(n_1570)
);

CKINVDCx14_ASAP7_75t_R g1571 ( 
.A(n_1401),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1415),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1401),
.Y(n_1573)
);

CKINVDCx6p67_ASAP7_75t_R g1574 ( 
.A(n_1386),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1504),
.A2(n_1495),
.B1(n_1427),
.B2(n_1444),
.Y(n_1575)
);

INVx6_ASAP7_75t_L g1576 ( 
.A(n_1482),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1519),
.A2(n_1432),
.B1(n_1394),
.B2(n_1374),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1407),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1472),
.A2(n_1400),
.B1(n_1441),
.B2(n_1467),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1416),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1503),
.A2(n_1405),
.B1(n_1531),
.B2(n_1544),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1538),
.A2(n_1461),
.B1(n_1460),
.B2(n_1494),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1473),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_1482),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1398),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1378),
.B(n_1479),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1485),
.A2(n_1486),
.B1(n_1403),
.B2(n_1457),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1457),
.A2(n_1418),
.B1(n_1547),
.B2(n_1464),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1525),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1448),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1507),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1467),
.A2(n_1543),
.B1(n_1434),
.B2(n_1509),
.Y(n_1592)
);

INVx2_ASAP7_75t_R g1593 ( 
.A(n_1517),
.Y(n_1593)
);

BUFx10_ASAP7_75t_L g1594 ( 
.A(n_1412),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1428),
.A2(n_1474),
.B1(n_1380),
.B2(n_1414),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1452),
.A2(n_1491),
.B(n_1431),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1500),
.Y(n_1597)
);

BUFx10_ASAP7_75t_L g1598 ( 
.A(n_1423),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1467),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1501),
.Y(n_1600)
);

OAI21xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1397),
.A2(n_1471),
.B(n_1404),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1434),
.A2(n_1516),
.B1(n_1489),
.B2(n_1496),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1508),
.Y(n_1603)
);

INVx4_ASAP7_75t_L g1604 ( 
.A(n_1406),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1397),
.A2(n_1498),
.B1(n_1548),
.B2(n_1475),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1434),
.A2(n_1510),
.B1(n_1382),
.B2(n_1499),
.Y(n_1606)
);

BUFx8_ASAP7_75t_L g1607 ( 
.A(n_1463),
.Y(n_1607)
);

INVx6_ASAP7_75t_L g1608 ( 
.A(n_1497),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1506),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1425),
.A2(n_1514),
.B1(n_1470),
.B2(n_1440),
.Y(n_1610)
);

BUFx8_ASAP7_75t_L g1611 ( 
.A(n_1435),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1406),
.A2(n_1511),
.B1(n_1505),
.B2(n_1425),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1513),
.B(n_1443),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1480),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1480),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1430),
.A2(n_1395),
.B1(n_1388),
.B2(n_1384),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_1484),
.Y(n_1617)
);

BUFx12f_ASAP7_75t_L g1618 ( 
.A(n_1497),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1502),
.Y(n_1619)
);

BUFx4_ASAP7_75t_R g1620 ( 
.A(n_1411),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1480),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1484),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1470),
.A2(n_1478),
.B1(n_1476),
.B2(n_1393),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1383),
.A2(n_1459),
.B1(n_1456),
.B2(n_1492),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1502),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1522),
.Y(n_1626)
);

BUFx8_ASAP7_75t_SL g1627 ( 
.A(n_1488),
.Y(n_1627)
);

INVx6_ASAP7_75t_L g1628 ( 
.A(n_1468),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1488),
.B(n_1468),
.Y(n_1629)
);

INVx4_ASAP7_75t_L g1630 ( 
.A(n_1411),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1453),
.Y(n_1631)
);

OAI22x1_ASAP7_75t_L g1632 ( 
.A1(n_1490),
.A2(n_1453),
.B1(n_1385),
.B2(n_1408),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1453),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1385),
.A2(n_1515),
.B1(n_1455),
.B2(n_1454),
.Y(n_1634)
);

NAND2x1p5_ASAP7_75t_L g1635 ( 
.A(n_1492),
.B(n_1442),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1442),
.A2(n_1402),
.B1(n_1387),
.B2(n_1421),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1408),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1522),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1385),
.B(n_1537),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1373),
.A2(n_1376),
.B1(n_1536),
.B2(n_1439),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1433),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1522),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1387),
.A2(n_1396),
.B1(n_1410),
.B2(n_1424),
.Y(n_1643)
);

BUFx12f_ASAP7_75t_L g1644 ( 
.A(n_1389),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1537),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1537),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1465),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1518),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1381),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1420),
.A2(n_1429),
.B1(n_1399),
.B2(n_1436),
.Y(n_1650)
);

CKINVDCx14_ASAP7_75t_R g1651 ( 
.A(n_1389),
.Y(n_1651)
);

OAI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1391),
.A2(n_1390),
.B1(n_1377),
.B2(n_1375),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1521),
.A2(n_1289),
.B1(n_1527),
.B2(n_1524),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1540),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1445),
.Y(n_1656)
);

OAI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1524),
.A2(n_1527),
.B1(n_1466),
.B2(n_1483),
.Y(n_1657)
);

CKINVDCx11_ASAP7_75t_R g1658 ( 
.A(n_1417),
.Y(n_1658)
);

BUFx2_ASAP7_75t_SL g1659 ( 
.A(n_1417),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1540),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1520),
.B(n_1530),
.Y(n_1661)
);

BUFx10_ASAP7_75t_L g1662 ( 
.A(n_1401),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1445),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1512),
.Y(n_1664)
);

BUFx12f_ASAP7_75t_L g1665 ( 
.A(n_1438),
.Y(n_1665)
);

CKINVDCx11_ASAP7_75t_R g1666 ( 
.A(n_1417),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1445),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1445),
.Y(n_1668)
);

BUFx12f_ASAP7_75t_L g1669 ( 
.A(n_1438),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1445),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1445),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1674)
);

CKINVDCx11_ASAP7_75t_R g1675 ( 
.A(n_1417),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1512),
.Y(n_1676)
);

CKINVDCx11_ASAP7_75t_R g1677 ( 
.A(n_1417),
.Y(n_1677)
);

INVx6_ASAP7_75t_L g1678 ( 
.A(n_1482),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1445),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1524),
.A2(n_1527),
.B1(n_1530),
.B2(n_1520),
.Y(n_1680)
);

BUFx8_ASAP7_75t_SL g1681 ( 
.A(n_1417),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1445),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1445),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1686)
);

INVx6_ASAP7_75t_L g1687 ( 
.A(n_1482),
.Y(n_1687)
);

CKINVDCx6p67_ASAP7_75t_R g1688 ( 
.A(n_1539),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1540),
.Y(n_1689)
);

INVx4_ASAP7_75t_L g1690 ( 
.A(n_1423),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1532),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1512),
.Y(n_1692)
);

CKINVDCx20_ASAP7_75t_R g1693 ( 
.A(n_1417),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1524),
.A2(n_1527),
.B1(n_893),
.B2(n_1289),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1445),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1520),
.B(n_1530),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1448),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1698)
);

BUFx2_ASAP7_75t_SL g1699 ( 
.A(n_1417),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1445),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1445),
.Y(n_1701)
);

INVx8_ASAP7_75t_L g1702 ( 
.A(n_1484),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_SL g1703 ( 
.A1(n_1529),
.A2(n_1289),
.B1(n_947),
.B2(n_1302),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1532),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1524),
.A2(n_1527),
.B1(n_1530),
.B2(n_1520),
.Y(n_1705)
);

BUFx8_ASAP7_75t_L g1706 ( 
.A(n_1401),
.Y(n_1706)
);

INVx6_ASAP7_75t_L g1707 ( 
.A(n_1482),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1524),
.A2(n_1527),
.B1(n_1530),
.B2(n_1520),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1524),
.A2(n_1527),
.B1(n_1530),
.B2(n_1520),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1445),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1529),
.A2(n_1289),
.B1(n_947),
.B2(n_1302),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1445),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1512),
.Y(n_1714)
);

BUFx12f_ASAP7_75t_L g1715 ( 
.A(n_1438),
.Y(n_1715)
);

BUFx8_ASAP7_75t_L g1716 ( 
.A(n_1401),
.Y(n_1716)
);

BUFx8_ASAP7_75t_L g1717 ( 
.A(n_1401),
.Y(n_1717)
);

INVx6_ASAP7_75t_L g1718 ( 
.A(n_1482),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1524),
.A2(n_1289),
.B1(n_1527),
.B2(n_1302),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1512),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1445),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1448),
.Y(n_1722)
);

CKINVDCx11_ASAP7_75t_R g1723 ( 
.A(n_1417),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1445),
.B(n_1392),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1651),
.B(n_1559),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1637),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1638),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1596),
.A2(n_1640),
.B(n_1650),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1645),
.Y(n_1729)
);

INVx4_ASAP7_75t_L g1730 ( 
.A(n_1567),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1651),
.B(n_1572),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1580),
.B(n_1583),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1639),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1556),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1656),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1557),
.A2(n_1595),
.B(n_1564),
.Y(n_1736)
);

OA21x2_ASAP7_75t_L g1737 ( 
.A1(n_1631),
.A2(n_1633),
.B(n_1615),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1562),
.B(n_1552),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1626),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1648),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1626),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1700),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1642),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1618),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1602),
.B(n_1642),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1700),
.Y(n_1746)
);

AO21x2_ASAP7_75t_L g1747 ( 
.A1(n_1614),
.A2(n_1621),
.B(n_1652),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1646),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1648),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1646),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1644),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1649),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_L g1753 ( 
.A1(n_1561),
.A2(n_1570),
.B(n_1554),
.C(n_1549),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1599),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1597),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1663),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1581),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1581),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1632),
.Y(n_1759)
);

CKINVDCx20_ASAP7_75t_R g1760 ( 
.A(n_1681),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1667),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1602),
.B(n_1668),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1650),
.A2(n_1643),
.B(n_1636),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1670),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1671),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1679),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1682),
.B(n_1684),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1695),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1724),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1701),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1703),
.A2(n_1711),
.B1(n_1657),
.B2(n_1550),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1703),
.A2(n_1711),
.B1(n_1657),
.B2(n_1550),
.Y(n_1772)
);

OAI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1643),
.A2(n_1636),
.B(n_1624),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1710),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1712),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1721),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1593),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1593),
.Y(n_1778)
);

AO21x1_ASAP7_75t_L g1779 ( 
.A1(n_1560),
.A2(n_1605),
.B(n_1680),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1606),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1606),
.Y(n_1781)
);

OA21x2_ASAP7_75t_L g1782 ( 
.A1(n_1653),
.A2(n_1575),
.B(n_1554),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1652),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1553),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1661),
.B(n_1696),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1654),
.A2(n_1698),
.B1(n_1719),
.B2(n_1713),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1600),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1628),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1654),
.A2(n_1672),
.B1(n_1673),
.B2(n_1686),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1647),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1647),
.Y(n_1791)
);

INVxp33_ASAP7_75t_L g1792 ( 
.A(n_1627),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1582),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1582),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1603),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1635),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1635),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1653),
.B(n_1549),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1705),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1592),
.Y(n_1800)
);

INVx4_ASAP7_75t_L g1801 ( 
.A(n_1567),
.Y(n_1801)
);

BUFx2_ASAP7_75t_SL g1802 ( 
.A(n_1617),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1592),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1708),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1616),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1601),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1624),
.A2(n_1612),
.B(n_1577),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1664),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1605),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1610),
.Y(n_1810)
);

AOI21x1_ASAP7_75t_L g1811 ( 
.A1(n_1709),
.A2(n_1625),
.B(n_1613),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1672),
.B(n_1673),
.Y(n_1812)
);

AOI21x1_ASAP7_75t_L g1813 ( 
.A1(n_1586),
.A2(n_1610),
.B(n_1623),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1608),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1611),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1674),
.B(n_1683),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1623),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1634),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1634),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1561),
.B(n_1570),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1558),
.B(n_1560),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1557),
.A2(n_1569),
.B(n_1575),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1579),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1674),
.A2(n_1719),
.B1(n_1713),
.B2(n_1698),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1579),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1691),
.Y(n_1826)
);

OAI21x1_ASAP7_75t_L g1827 ( 
.A1(n_1587),
.A2(n_1629),
.B(n_1565),
.Y(n_1827)
);

OAI21x1_ASAP7_75t_L g1828 ( 
.A1(n_1587),
.A2(n_1629),
.B(n_1565),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1704),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1704),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1608),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1558),
.B(n_1694),
.Y(n_1832)
);

OAI21x1_ASAP7_75t_L g1833 ( 
.A1(n_1588),
.A2(n_1686),
.B(n_1685),
.Y(n_1833)
);

OAI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1588),
.A2(n_1685),
.B(n_1683),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1704),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1641),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1604),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1604),
.Y(n_1838)
);

INVx2_ASAP7_75t_SL g1839 ( 
.A(n_1608),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1619),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1578),
.A2(n_1589),
.B1(n_1574),
.B2(n_1718),
.Y(n_1841)
);

AOI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1676),
.A2(n_1692),
.B(n_1720),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1622),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1622),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1690),
.Y(n_1845)
);

INVx6_ASAP7_75t_L g1846 ( 
.A(n_1611),
.Y(n_1846)
);

NAND2x1p5_ASAP7_75t_L g1847 ( 
.A(n_1590),
.B(n_1697),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1590),
.Y(n_1848)
);

BUFx3_ASAP7_75t_L g1849 ( 
.A(n_1697),
.Y(n_1849)
);

CKINVDCx11_ASAP7_75t_R g1850 ( 
.A(n_1566),
.Y(n_1850)
);

A2O1A1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1722),
.A2(n_1585),
.B(n_1664),
.C(n_1591),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1568),
.B(n_1714),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1598),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1662),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1598),
.Y(n_1855)
);

OAI21x1_ASAP7_75t_L g1856 ( 
.A1(n_1702),
.A2(n_1662),
.B(n_1571),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1702),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1702),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1594),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1594),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1571),
.B(n_1573),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1576),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1551),
.B(n_1688),
.Y(n_1863)
);

INVx2_ASAP7_75t_SL g1864 ( 
.A(n_1576),
.Y(n_1864)
);

INVx2_ASAP7_75t_SL g1865 ( 
.A(n_1576),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1607),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1630),
.B(n_1609),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1678),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1787),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1769),
.B(n_1699),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1799),
.B(n_1607),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1808),
.B(n_1659),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1786),
.A2(n_1707),
.B1(n_1687),
.B2(n_1678),
.Y(n_1873)
);

OAI21x1_ASAP7_75t_SL g1874 ( 
.A1(n_1779),
.A2(n_1630),
.B(n_1620),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1850),
.B(n_1655),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1808),
.B(n_1784),
.Y(n_1876)
);

OAI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1736),
.A2(n_1660),
.B(n_1584),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1789),
.A2(n_1687),
.B1(n_1718),
.B2(n_1707),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1742),
.B(n_1689),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1822),
.A2(n_1693),
.B(n_1620),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1732),
.B(n_1716),
.Y(n_1881)
);

A2O1A1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1771),
.A2(n_1555),
.B(n_1563),
.C(n_1715),
.Y(n_1882)
);

AOI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1779),
.A2(n_1665),
.B1(n_1669),
.B2(n_1716),
.C(n_1717),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1802),
.B(n_1718),
.Y(n_1884)
);

AOI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1821),
.A2(n_1706),
.B1(n_1717),
.B2(n_1675),
.C(n_1677),
.Y(n_1885)
);

OAI211xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1859),
.A2(n_1658),
.B(n_1666),
.C(n_1723),
.Y(n_1886)
);

OA21x2_ASAP7_75t_L g1887 ( 
.A1(n_1728),
.A2(n_1706),
.B(n_1817),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1746),
.B(n_1756),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1804),
.B(n_1757),
.Y(n_1889)
);

INVxp67_ASAP7_75t_SL g1890 ( 
.A(n_1836),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1725),
.B(n_1731),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1755),
.Y(n_1892)
);

AND2x4_ASAP7_75t_SL g1893 ( 
.A(n_1867),
.B(n_1862),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1802),
.B(n_1849),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1756),
.B(n_1776),
.Y(n_1895)
);

A2O1A1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1772),
.A2(n_1753),
.B(n_1807),
.C(n_1812),
.Y(n_1896)
);

BUFx3_ASAP7_75t_L g1897 ( 
.A(n_1815),
.Y(n_1897)
);

OAI21x1_ASAP7_75t_SL g1898 ( 
.A1(n_1842),
.A2(n_1820),
.B(n_1766),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1852),
.B(n_1762),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1849),
.B(n_1864),
.Y(n_1900)
);

AND4x1_ASAP7_75t_L g1901 ( 
.A(n_1851),
.B(n_1863),
.C(n_1824),
.D(n_1823),
.Y(n_1901)
);

OAI211xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1859),
.A2(n_1860),
.B(n_1806),
.C(n_1805),
.Y(n_1902)
);

OAI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1807),
.A2(n_1805),
.B(n_1809),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1757),
.B(n_1758),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1760),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1809),
.A2(n_1758),
.B(n_1798),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1767),
.B(n_1861),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1864),
.B(n_1865),
.Y(n_1908)
);

O2A1O1Ixp33_ASAP7_75t_L g1909 ( 
.A1(n_1832),
.A2(n_1818),
.B(n_1819),
.C(n_1806),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1861),
.B(n_1761),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1773),
.A2(n_1763),
.B(n_1818),
.Y(n_1911)
);

O2A1O1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1819),
.A2(n_1798),
.B(n_1817),
.C(n_1810),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1766),
.B(n_1749),
.Y(n_1913)
);

CKINVDCx20_ASAP7_75t_R g1914 ( 
.A(n_1815),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1812),
.A2(n_1816),
.B1(n_1823),
.B2(n_1825),
.Y(n_1915)
);

OR2x6_ASAP7_75t_L g1916 ( 
.A(n_1827),
.B(n_1828),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1825),
.A2(n_1816),
.B1(n_1803),
.B2(n_1800),
.Y(n_1917)
);

AOI21xp33_ASAP7_75t_L g1918 ( 
.A1(n_1810),
.A2(n_1782),
.B(n_1781),
.Y(n_1918)
);

A2O1A1Ixp33_ASAP7_75t_L g1919 ( 
.A1(n_1833),
.A2(n_1834),
.B(n_1781),
.C(n_1780),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1744),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1782),
.A2(n_1834),
.B(n_1833),
.Y(n_1921)
);

OR2x6_ASAP7_75t_L g1922 ( 
.A(n_1827),
.B(n_1828),
.Y(n_1922)
);

CKINVDCx6p67_ASAP7_75t_R g1923 ( 
.A(n_1744),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_SL g1924 ( 
.A1(n_1782),
.A2(n_1745),
.B1(n_1803),
.B2(n_1800),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1749),
.B(n_1764),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1780),
.A2(n_1794),
.B(n_1793),
.C(n_1783),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1846),
.Y(n_1927)
);

AOI221xp5_ASAP7_75t_L g1928 ( 
.A1(n_1783),
.A2(n_1785),
.B1(n_1738),
.B2(n_1734),
.C(n_1735),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1765),
.B(n_1768),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1733),
.B(n_1768),
.Y(n_1930)
);

NAND3xp33_ASAP7_75t_L g1931 ( 
.A(n_1759),
.B(n_1782),
.C(n_1848),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1770),
.B(n_1774),
.Y(n_1932)
);

NAND2xp33_ASAP7_75t_R g1933 ( 
.A(n_1863),
.B(n_1867),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1775),
.B(n_1740),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1775),
.B(n_1842),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1848),
.Y(n_1936)
);

AND2x4_ASAP7_75t_SL g1937 ( 
.A(n_1867),
.B(n_1868),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1751),
.B(n_1813),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1754),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1733),
.B(n_1754),
.Y(n_1940)
);

A2O1A1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1759),
.A2(n_1796),
.B(n_1797),
.C(n_1856),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1727),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1740),
.B(n_1868),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1846),
.A2(n_1847),
.B1(n_1866),
.B2(n_1841),
.Y(n_1944)
);

AO32x2_ASAP7_75t_L g1945 ( 
.A1(n_1814),
.A2(n_1839),
.A3(n_1831),
.B1(n_1788),
.B2(n_1801),
.Y(n_1945)
);

OA21x2_ASAP7_75t_L g1946 ( 
.A1(n_1777),
.A2(n_1778),
.B(n_1791),
.Y(n_1946)
);

AOI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1739),
.A2(n_1741),
.B1(n_1743),
.B2(n_1748),
.C(n_1750),
.Y(n_1947)
);

AO32x2_ASAP7_75t_L g1948 ( 
.A1(n_1814),
.A2(n_1839),
.A3(n_1831),
.B1(n_1788),
.B2(n_1801),
.Y(n_1948)
);

AO21x1_ASAP7_75t_L g1949 ( 
.A1(n_1847),
.A2(n_1811),
.B(n_1791),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1727),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1729),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1840),
.B(n_1739),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1811),
.A2(n_1743),
.B(n_1748),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1741),
.B(n_1750),
.Y(n_1954)
);

AO32x2_ASAP7_75t_L g1955 ( 
.A1(n_1730),
.A2(n_1801),
.A3(n_1854),
.B1(n_1795),
.B2(n_1840),
.Y(n_1955)
);

OA21x2_ASAP7_75t_L g1956 ( 
.A1(n_1777),
.A2(n_1778),
.B(n_1726),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1956),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1889),
.B(n_1752),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1954),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1956),
.Y(n_1960)
);

OAI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1896),
.A2(n_1847),
.B1(n_1797),
.B2(n_1796),
.C(n_1853),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1888),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1899),
.B(n_1790),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1954),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1946),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1886),
.B(n_1792),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1939),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1942),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1950),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1883),
.A2(n_1846),
.B1(n_1853),
.B2(n_1855),
.Y(n_1970)
);

BUFx2_ASAP7_75t_L g1971 ( 
.A(n_1945),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1951),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1915),
.A2(n_1846),
.B1(n_1729),
.B2(n_1726),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1935),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1892),
.Y(n_1975)
);

AOI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1915),
.A2(n_1855),
.B1(n_1835),
.B2(n_1826),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1943),
.B(n_1747),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1916),
.B(n_1747),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1946),
.Y(n_1979)
);

NAND2x1_ASAP7_75t_L g1980 ( 
.A(n_1898),
.B(n_1837),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1891),
.B(n_1837),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1930),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1930),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1907),
.B(n_1830),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1940),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1910),
.B(n_1895),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1940),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1893),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1955),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1927),
.B(n_1854),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_1905),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1880),
.A2(n_1829),
.B1(n_1843),
.B2(n_1844),
.Y(n_1992)
);

AOI21xp33_ASAP7_75t_SL g1993 ( 
.A1(n_1933),
.A2(n_1856),
.B(n_1858),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1955),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1955),
.Y(n_1995)
);

INVxp67_ASAP7_75t_SL g1996 ( 
.A(n_1890),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1934),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1925),
.B(n_1845),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1869),
.B(n_1737),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1952),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1913),
.B(n_1934),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1876),
.B(n_1845),
.Y(n_2002)
);

INVxp67_ASAP7_75t_SL g2003 ( 
.A(n_1949),
.Y(n_2003)
);

NOR2xp67_ASAP7_75t_L g2004 ( 
.A(n_1931),
.B(n_1838),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1932),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1929),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1936),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1945),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1945),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1948),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1971),
.B(n_1872),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1980),
.Y(n_2012)
);

OAI33xp33_ASAP7_75t_L g2013 ( 
.A1(n_1970),
.A2(n_1909),
.A3(n_1873),
.B1(n_1878),
.B2(n_1931),
.B3(n_1944),
.Y(n_2013)
);

OAI22xp33_ASAP7_75t_L g2014 ( 
.A1(n_1973),
.A2(n_1880),
.B1(n_1873),
.B2(n_1878),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1971),
.B(n_1938),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1996),
.B(n_1903),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_2004),
.B(n_1916),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1962),
.B(n_1911),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1974),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1999),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1973),
.A2(n_1883),
.B1(n_1944),
.B2(n_1924),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1999),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_2003),
.A2(n_1902),
.B(n_1877),
.Y(n_2023)
);

OAI211xp5_ASAP7_75t_L g2024 ( 
.A1(n_2004),
.A2(n_1877),
.B(n_1885),
.C(n_1902),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1962),
.B(n_1903),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1967),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_SL g2027 ( 
.A1(n_1970),
.A2(n_1885),
.B(n_1901),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1957),
.Y(n_2028)
);

INVxp67_ASAP7_75t_SL g2029 ( 
.A(n_1989),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1957),
.Y(n_2030)
);

OAI221xp5_ASAP7_75t_SL g2031 ( 
.A1(n_1976),
.A2(n_1909),
.B1(n_1912),
.B2(n_1928),
.C(n_1911),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1957),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1960),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1982),
.B(n_1928),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_2000),
.B(n_1904),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1977),
.B(n_1997),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1967),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_2007),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1986),
.B(n_1870),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_2007),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_R g2041 ( 
.A(n_1991),
.B(n_1914),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1960),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1960),
.Y(n_2043)
);

BUFx3_ASAP7_75t_L g2044 ( 
.A(n_1980),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1968),
.Y(n_2045)
);

INVx2_ASAP7_75t_SL g2046 ( 
.A(n_2001),
.Y(n_2046)
);

OAI31xp33_ASAP7_75t_L g2047 ( 
.A1(n_1961),
.A2(n_1926),
.A3(n_1912),
.B(n_1882),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1968),
.Y(n_2048)
);

OAI221xp5_ASAP7_75t_L g2049 ( 
.A1(n_1976),
.A2(n_1919),
.B1(n_1906),
.B2(n_1917),
.C(n_1918),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1969),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2001),
.B(n_1948),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1963),
.B(n_1948),
.Y(n_2052)
);

NAND2xp33_ASAP7_75t_R g2053 ( 
.A(n_1993),
.B(n_1920),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1969),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1972),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_2005),
.B(n_1958),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1972),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1965),
.Y(n_2058)
);

OAI31xp33_ASAP7_75t_L g2059 ( 
.A1(n_1989),
.A2(n_1918),
.A3(n_1941),
.B(n_1871),
.Y(n_2059)
);

AND2x4_ASAP7_75t_L g2060 ( 
.A(n_1977),
.B(n_1922),
.Y(n_2060)
);

OAI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_1992),
.A2(n_1871),
.B1(n_1879),
.B2(n_1881),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1983),
.B(n_1947),
.Y(n_2062)
);

OR2x6_ASAP7_75t_L g2063 ( 
.A(n_1978),
.B(n_1922),
.Y(n_2063)
);

AOI33xp33_ASAP7_75t_L g2064 ( 
.A1(n_1989),
.A2(n_1995),
.A3(n_1994),
.B1(n_2009),
.B2(n_2008),
.B3(n_2010),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_1997),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_1998),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1975),
.Y(n_2067)
);

INVx3_ASAP7_75t_L g2068 ( 
.A(n_1997),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1988),
.Y(n_2069)
);

INVx2_ASAP7_75t_SL g2070 ( 
.A(n_2012),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2026),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2026),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2062),
.B(n_1983),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2052),
.B(n_1994),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2052),
.B(n_1994),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2028),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_2016),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2064),
.B(n_2034),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2028),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2051),
.B(n_1995),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2020),
.B(n_2008),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2051),
.B(n_1995),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2037),
.B(n_1985),
.Y(n_2083)
);

INVxp67_ASAP7_75t_SL g2084 ( 
.A(n_2023),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2015),
.B(n_2009),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2037),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2020),
.B(n_2010),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2045),
.B(n_1985),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2045),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2015),
.B(n_2006),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_2012),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2048),
.B(n_1987),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2065),
.B(n_2006),
.Y(n_2093)
);

BUFx2_ASAP7_75t_L g2094 ( 
.A(n_2044),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_2036),
.B(n_1977),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2065),
.B(n_1998),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2028),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2048),
.B(n_1987),
.Y(n_2098)
);

INVxp67_ASAP7_75t_SL g2099 ( 
.A(n_2018),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2050),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2050),
.B(n_1959),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2054),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2068),
.B(n_1981),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2054),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2055),
.Y(n_2105)
);

OAI321xp33_ASAP7_75t_L g2106 ( 
.A1(n_2031),
.A2(n_1906),
.A3(n_1992),
.B1(n_1921),
.B2(n_1953),
.C(n_1979),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_2036),
.B(n_2017),
.Y(n_2107)
);

INVxp67_ASAP7_75t_SL g2108 ( 
.A(n_2018),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2055),
.B(n_1959),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2068),
.B(n_2002),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_2022),
.B(n_1964),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2068),
.B(n_2002),
.Y(n_2112)
);

OA21x2_ASAP7_75t_L g2113 ( 
.A1(n_2030),
.A2(n_1979),
.B(n_1965),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2030),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_2027),
.B(n_2024),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2030),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2057),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2057),
.B(n_1964),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2011),
.B(n_1984),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2073),
.B(n_2056),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2071),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2084),
.B(n_2025),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2071),
.Y(n_2123)
);

AOI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_2084),
.A2(n_2013),
.B1(n_2021),
.B2(n_2049),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2073),
.B(n_2038),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2078),
.B(n_2056),
.Y(n_2126)
);

INVx2_ASAP7_75t_SL g2127 ( 
.A(n_2094),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_2115),
.B(n_1923),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2119),
.B(n_2044),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2077),
.B(n_2078),
.Y(n_2130)
);

INVx1_ASAP7_75t_SL g2131 ( 
.A(n_2115),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2077),
.B(n_2040),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2071),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2086),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2119),
.B(n_2044),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2086),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2119),
.B(n_2011),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2080),
.B(n_2069),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_2107),
.B(n_2095),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2086),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2080),
.B(n_2069),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2080),
.B(n_2069),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_2099),
.B(n_2022),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2099),
.B(n_2035),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2108),
.B(n_2035),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2108),
.B(n_2019),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2102),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2113),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2083),
.B(n_2067),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2082),
.B(n_2074),
.Y(n_2150)
);

AOI21xp33_ASAP7_75t_SL g2151 ( 
.A1(n_2070),
.A2(n_2053),
.B(n_2061),
.Y(n_2151)
);

INVx2_ASAP7_75t_SL g2152 ( 
.A(n_2094),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2113),
.Y(n_2153)
);

INVx4_ASAP7_75t_L g2154 ( 
.A(n_2094),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2102),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2082),
.B(n_2074),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2082),
.B(n_2074),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2102),
.Y(n_2158)
);

INVx3_ASAP7_75t_L g2159 ( 
.A(n_2107),
.Y(n_2159)
);

INVxp67_ASAP7_75t_L g2160 ( 
.A(n_2070),
.Y(n_2160)
);

INVxp67_ASAP7_75t_SL g2161 ( 
.A(n_2091),
.Y(n_2161)
);

NOR2x1_ASAP7_75t_L g2162 ( 
.A(n_2091),
.B(n_1897),
.Y(n_2162)
);

OAI22xp33_ASAP7_75t_L g2163 ( 
.A1(n_2106),
.A2(n_2014),
.B1(n_1993),
.B2(n_2063),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2104),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2104),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2104),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2075),
.B(n_2012),
.Y(n_2167)
);

NAND3xp33_ASAP7_75t_L g2168 ( 
.A(n_2105),
.B(n_2059),
.C(n_2047),
.Y(n_2168)
);

OAI31xp33_ASAP7_75t_L g2169 ( 
.A1(n_2085),
.A2(n_2047),
.A3(n_2106),
.B(n_2075),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2075),
.B(n_2012),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2083),
.B(n_2067),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2124),
.B(n_2090),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2123),
.Y(n_2173)
);

NOR3xp33_ASAP7_75t_L g2174 ( 
.A(n_2131),
.B(n_2091),
.C(n_2070),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2130),
.B(n_2090),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2150),
.B(n_2085),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2150),
.B(n_2085),
.Y(n_2177)
);

AOI211xp5_ASAP7_75t_SL g2178 ( 
.A1(n_2163),
.A2(n_2122),
.B(n_2159),
.C(n_2128),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2123),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2156),
.B(n_2096),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2169),
.B(n_2090),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_2168),
.B(n_1875),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2156),
.B(n_2096),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_2151),
.B(n_2012),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2157),
.B(n_2096),
.Y(n_2185)
);

INVxp67_ASAP7_75t_L g2186 ( 
.A(n_2126),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2126),
.A2(n_1921),
.B1(n_2017),
.B2(n_2060),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2120),
.B(n_2072),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2134),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2157),
.B(n_2107),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2134),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_2127),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2120),
.B(n_2072),
.Y(n_2193)
);

INVx2_ASAP7_75t_SL g2194 ( 
.A(n_2138),
.Y(n_2194)
);

INVx1_ASAP7_75t_SL g2195 ( 
.A(n_2127),
.Y(n_2195)
);

OAI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2139),
.A2(n_2107),
.B1(n_2046),
.B2(n_2066),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2138),
.B(n_2107),
.Y(n_2197)
);

OAI21xp33_ASAP7_75t_L g2198 ( 
.A1(n_2132),
.A2(n_2087),
.B(n_2081),
.Y(n_2198)
);

INVx2_ASAP7_75t_SL g2199 ( 
.A(n_2141),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_2139),
.B(n_2107),
.Y(n_2200)
);

NAND3xp33_ASAP7_75t_SL g2201 ( 
.A(n_2146),
.B(n_2041),
.C(n_1894),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2125),
.B(n_2089),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2136),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2141),
.B(n_2103),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2136),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2140),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2144),
.B(n_2089),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2148),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_2154),
.B(n_1966),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_2139),
.B(n_2095),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2140),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2144),
.B(n_2100),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2148),
.Y(n_2213)
);

NOR2x1_ASAP7_75t_L g2214 ( 
.A(n_2182),
.B(n_2154),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2190),
.Y(n_2215)
);

HB1xp67_ASAP7_75t_L g2216 ( 
.A(n_2192),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2173),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2197),
.B(n_2200),
.Y(n_2218)
);

AOI22xp33_ASAP7_75t_L g2219 ( 
.A1(n_2172),
.A2(n_2153),
.B1(n_2142),
.B2(n_2017),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_2200),
.B(n_2152),
.Y(n_2220)
);

AOI221xp5_ASAP7_75t_L g2221 ( 
.A1(n_2181),
.A2(n_2153),
.B1(n_2029),
.B2(n_2165),
.C(n_2145),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2186),
.A2(n_2142),
.B1(n_2159),
.B2(n_2137),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2195),
.B(n_2194),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2173),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2195),
.B(n_2137),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2194),
.B(n_2152),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2179),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_L g2228 ( 
.A1(n_2187),
.A2(n_2017),
.B1(n_2170),
.B2(n_2167),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_2200),
.B(n_2154),
.Y(n_2229)
);

OAI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_2200),
.A2(n_2159),
.B1(n_2129),
.B2(n_2135),
.Y(n_2230)
);

AOI21xp33_ASAP7_75t_L g2231 ( 
.A1(n_2209),
.A2(n_2143),
.B(n_2145),
.Y(n_2231)
);

O2A1O1Ixp33_ASAP7_75t_R g2232 ( 
.A1(n_2178),
.A2(n_2143),
.B(n_2087),
.C(n_2081),
.Y(n_2232)
);

OAI221xp5_ASAP7_75t_L g2233 ( 
.A1(n_2198),
.A2(n_2170),
.B1(n_2167),
.B2(n_2087),
.C(n_2081),
.Y(n_2233)
);

INVxp67_ASAP7_75t_SL g2234 ( 
.A(n_2174),
.Y(n_2234)
);

OAI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_2198),
.A2(n_2162),
.B1(n_2079),
.B2(n_2097),
.C(n_2076),
.Y(n_2235)
);

NAND4xp25_ASAP7_75t_L g2236 ( 
.A(n_2201),
.B(n_2129),
.C(n_2135),
.D(n_2160),
.Y(n_2236)
);

O2A1O1Ixp5_ASAP7_75t_L g2237 ( 
.A1(n_2184),
.A2(n_2212),
.B(n_2207),
.C(n_2196),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2199),
.B(n_2175),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_2199),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2179),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2176),
.B(n_2149),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2197),
.B(n_2091),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2190),
.Y(n_2243)
);

AOI21xp33_ASAP7_75t_L g2244 ( 
.A1(n_2234),
.A2(n_2213),
.B(n_2208),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2217),
.Y(n_2245)
);

OAI21xp33_ASAP7_75t_L g2246 ( 
.A1(n_2236),
.A2(n_2193),
.B(n_2188),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2225),
.B(n_2202),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2218),
.B(n_2176),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2217),
.Y(n_2249)
);

OAI21xp33_ASAP7_75t_L g2250 ( 
.A1(n_2219),
.A2(n_2221),
.B(n_2214),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2237),
.A2(n_2213),
.B(n_2208),
.Y(n_2251)
);

AOI22xp33_ASAP7_75t_L g2252 ( 
.A1(n_2231),
.A2(n_2213),
.B1(n_2208),
.B2(n_1874),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2218),
.B(n_2177),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2215),
.B(n_2177),
.Y(n_2254)
);

OAI21xp5_ASAP7_75t_SL g2255 ( 
.A1(n_2232),
.A2(n_2210),
.B(n_2204),
.Y(n_2255)
);

AOI322xp5_ASAP7_75t_L g2256 ( 
.A1(n_2232),
.A2(n_2185),
.A3(n_2180),
.B1(n_2183),
.B2(n_2205),
.C1(n_2206),
.C2(n_2203),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2240),
.Y(n_2257)
);

OAI32xp33_ASAP7_75t_L g2258 ( 
.A1(n_2235),
.A2(n_2211),
.A3(n_2206),
.B1(n_2205),
.B2(n_2189),
.Y(n_2258)
);

AO22x1_ASAP7_75t_L g2259 ( 
.A1(n_2220),
.A2(n_2210),
.B1(n_2161),
.B2(n_1884),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2239),
.B(n_2180),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2220),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2239),
.B(n_2183),
.Y(n_2262)
);

NOR2xp33_ASAP7_75t_L g2263 ( 
.A(n_2216),
.B(n_2210),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2228),
.A2(n_2210),
.B1(n_2042),
.B2(n_2058),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2240),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2223),
.B(n_2185),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2248),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2248),
.Y(n_2268)
);

INVxp67_ASAP7_75t_L g2269 ( 
.A(n_2263),
.Y(n_2269)
);

INVx1_ASAP7_75t_SL g2270 ( 
.A(n_2261),
.Y(n_2270)
);

INVxp67_ASAP7_75t_L g2271 ( 
.A(n_2263),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_L g2272 ( 
.A(n_2261),
.B(n_2229),
.Y(n_2272)
);

AO22x2_ASAP7_75t_L g2273 ( 
.A1(n_2251),
.A2(n_2224),
.B1(n_2227),
.B2(n_2215),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2253),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2255),
.A2(n_2243),
.B1(n_2222),
.B2(n_2230),
.Y(n_2275)
);

AOI21xp5_ASAP7_75t_L g2276 ( 
.A1(n_2258),
.A2(n_2229),
.B(n_2220),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2253),
.B(n_2243),
.Y(n_2277)
);

AOI221xp5_ASAP7_75t_L g2278 ( 
.A1(n_2244),
.A2(n_2233),
.B1(n_2238),
.B2(n_2189),
.C(n_2191),
.Y(n_2278)
);

AOI221xp5_ASAP7_75t_L g2279 ( 
.A1(n_2250),
.A2(n_2191),
.B1(n_2211),
.B2(n_2203),
.C(n_2226),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_2256),
.B(n_2012),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2254),
.B(n_2260),
.Y(n_2281)
);

NOR3xp33_ASAP7_75t_L g2282 ( 
.A(n_2269),
.B(n_2259),
.C(n_2246),
.Y(n_2282)
);

NAND5xp2_ASAP7_75t_L g2283 ( 
.A(n_2272),
.B(n_2262),
.C(n_2266),
.D(n_2249),
.E(n_2265),
.Y(n_2283)
);

NAND3xp33_ASAP7_75t_L g2284 ( 
.A(n_2279),
.B(n_2271),
.C(n_2276),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2267),
.B(n_2247),
.Y(n_2285)
);

AOI21xp5_ASAP7_75t_SL g2286 ( 
.A1(n_2281),
.A2(n_2257),
.B(n_2245),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2268),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2274),
.B(n_2204),
.Y(n_2288)
);

NAND3xp33_ASAP7_75t_SL g2289 ( 
.A(n_2270),
.B(n_2252),
.C(n_2264),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2277),
.B(n_2241),
.Y(n_2290)
);

AOI211xp5_ASAP7_75t_L g2291 ( 
.A1(n_2280),
.A2(n_2242),
.B(n_2252),
.C(n_2165),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_L g2292 ( 
.A(n_2275),
.B(n_2242),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2273),
.B(n_2039),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2273),
.B(n_2039),
.Y(n_2294)
);

NAND3xp33_ASAP7_75t_L g2295 ( 
.A(n_2278),
.B(n_2133),
.C(n_2121),
.Y(n_2295)
);

AOI221xp5_ASAP7_75t_L g2296 ( 
.A1(n_2289),
.A2(n_2147),
.B1(n_2166),
.B2(n_2164),
.C(n_2158),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2288),
.Y(n_2297)
);

AOI222xp33_ASAP7_75t_L g2298 ( 
.A1(n_2284),
.A2(n_2097),
.B1(n_2114),
.B2(n_2079),
.C1(n_2076),
.C2(n_2116),
.Y(n_2298)
);

A2O1A1Ixp33_ASAP7_75t_L g2299 ( 
.A1(n_2291),
.A2(n_2091),
.B(n_2116),
.C(n_2079),
.Y(n_2299)
);

AOI21xp33_ASAP7_75t_L g2300 ( 
.A1(n_2292),
.A2(n_2285),
.B(n_2290),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2287),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2282),
.B(n_2155),
.Y(n_2302)
);

AOI22xp33_ASAP7_75t_SL g2303 ( 
.A1(n_2293),
.A2(n_2095),
.B1(n_2079),
.B2(n_2116),
.Y(n_2303)
);

NOR2x1p5_ASAP7_75t_L g2304 ( 
.A(n_2295),
.B(n_2171),
.Y(n_2304)
);

NAND4xp75_ASAP7_75t_L g2305 ( 
.A(n_2294),
.B(n_1887),
.C(n_2113),
.D(n_1990),
.Y(n_2305)
);

INVxp67_ASAP7_75t_SL g2306 ( 
.A(n_2297),
.Y(n_2306)
);

OR2x2_ASAP7_75t_L g2307 ( 
.A(n_2301),
.B(n_2283),
.Y(n_2307)
);

AOI221xp5_ASAP7_75t_L g2308 ( 
.A1(n_2296),
.A2(n_2283),
.B1(n_2286),
.B2(n_2076),
.C(n_2097),
.Y(n_2308)
);

AOI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2300),
.A2(n_2097),
.B1(n_2076),
.B2(n_2116),
.C(n_2114),
.Y(n_2309)
);

NOR4xp25_ASAP7_75t_L g2310 ( 
.A(n_2302),
.B(n_2105),
.C(n_2117),
.D(n_2100),
.Y(n_2310)
);

AOI211x1_ASAP7_75t_L g2311 ( 
.A1(n_2304),
.A2(n_2105),
.B(n_2117),
.C(n_2098),
.Y(n_2311)
);

NOR2xp67_ASAP7_75t_L g2312 ( 
.A(n_2303),
.B(n_2111),
.Y(n_2312)
);

OAI21xp5_ASAP7_75t_SL g2313 ( 
.A1(n_2299),
.A2(n_1937),
.B(n_2112),
.Y(n_2313)
);

NAND3xp33_ASAP7_75t_L g2314 ( 
.A(n_2307),
.B(n_2298),
.C(n_2305),
.Y(n_2314)
);

AOI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_2306),
.A2(n_2118),
.B(n_2109),
.Y(n_2315)
);

NAND4xp75_ASAP7_75t_L g2316 ( 
.A(n_2308),
.B(n_2113),
.C(n_2093),
.D(n_1887),
.Y(n_2316)
);

NAND4xp75_ASAP7_75t_L g2317 ( 
.A(n_2311),
.B(n_2113),
.C(n_2093),
.D(n_2114),
.Y(n_2317)
);

INVx5_ASAP7_75t_L g2318 ( 
.A(n_2310),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2312),
.Y(n_2319)
);

NOR2xp67_ASAP7_75t_L g2320 ( 
.A(n_2318),
.B(n_2313),
.Y(n_2320)
);

XOR2xp5_ASAP7_75t_L g2321 ( 
.A(n_2314),
.B(n_2095),
.Y(n_2321)
);

NOR3xp33_ASAP7_75t_SL g2322 ( 
.A(n_2319),
.B(n_2309),
.C(n_1900),
.Y(n_2322)
);

OAI22x1_ASAP7_75t_L g2323 ( 
.A1(n_2317),
.A2(n_2095),
.B1(n_2114),
.B2(n_2036),
.Y(n_2323)
);

INVx1_ASAP7_75t_SL g2324 ( 
.A(n_2321),
.Y(n_2324)
);

OAI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2324),
.A2(n_2320),
.B1(n_2316),
.B2(n_2322),
.Y(n_2325)
);

AOI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_2325),
.A2(n_2323),
.B(n_2315),
.Y(n_2326)
);

AO22x2_ASAP7_75t_L g2327 ( 
.A1(n_2325),
.A2(n_2095),
.B1(n_2111),
.B2(n_2088),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2327),
.A2(n_2113),
.B1(n_2111),
.B2(n_2043),
.Y(n_2328)
);

BUFx2_ASAP7_75t_L g2329 ( 
.A(n_2326),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2329),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2328),
.A2(n_2118),
.B(n_2088),
.Y(n_2331)
);

AOI22xp33_ASAP7_75t_L g2332 ( 
.A1(n_2330),
.A2(n_2331),
.B1(n_2033),
.B2(n_2032),
.Y(n_2332)
);

OAI21xp33_ASAP7_75t_SL g2333 ( 
.A1(n_2332),
.A2(n_2112),
.B(n_2110),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2333),
.Y(n_2334)
);

AOI221xp5_ASAP7_75t_L g2335 ( 
.A1(n_2334),
.A2(n_2098),
.B1(n_2092),
.B2(n_2101),
.C(n_2109),
.Y(n_2335)
);

AOI211xp5_ASAP7_75t_L g2336 ( 
.A1(n_2335),
.A2(n_1908),
.B(n_1857),
.C(n_1858),
.Y(n_2336)
);


endmodule