module real_jpeg_12621_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_57;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_58;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_59;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_56;
wire n_30;
wire n_48;
wire n_16;
wire n_15;
wire n_13;

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_11),
.B1(n_20),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_4),
.A2(n_11),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_4),
.A2(n_21),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_5),
.B(n_15),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_5),
.A2(n_11),
.B1(n_20),
.B2(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_5),
.A2(n_25),
.B1(n_44),
.B2(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_11),
.C(n_34),
.Y(n_53)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_37),
.Y(n_7)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_26),
.B(n_36),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_17),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_14),
.Y(n_10)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_16),
.Y(n_23)
);

AO22x1_ASAP7_75t_L g33 ( 
.A1(n_11),
.A2(n_20),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_22),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_35),
.B1(n_44),
.B2(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_59),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_56),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);


endmodule