module fake_jpeg_30371_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

MAJIxp5_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_2),
.C(n_5),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_0),
.C(n_1),
.Y(n_18)
);

NAND2xp67_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_20),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_9),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_15),
.B1(n_9),
.B2(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_10),
.B(n_8),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_29),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_24),
.C(n_20),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_33),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_7),
.C(n_12),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_6),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_27),
.B1(n_6),
.B2(n_4),
.Y(n_39)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_39),
.Y(n_40)
);

AO21x1_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_17),
.B(n_1),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_3),
.C(n_38),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_17),
.C(n_3),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_45),
.C(n_36),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g48 ( 
.A(n_46),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_47),
.B(n_44),
.Y(n_49)
);


endmodule