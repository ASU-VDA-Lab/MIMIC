module real_aes_1020_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_735;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g247 ( .A(n_0), .B(n_154), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_1), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_2), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_3), .B(n_143), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_4), .B(n_152), .Y(n_482) );
INVx1_ASAP7_75t_L g142 ( .A(n_5), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_6), .B(n_143), .Y(n_200) );
NAND2xp33_ASAP7_75t_SL g193 ( .A(n_7), .B(n_149), .Y(n_193) );
INVx1_ASAP7_75t_L g173 ( .A(n_8), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g768 ( .A(n_9), .Y(n_768) );
AND2x2_ASAP7_75t_L g198 ( .A(n_10), .B(n_133), .Y(n_198) );
AND2x2_ASAP7_75t_L g475 ( .A(n_11), .B(n_190), .Y(n_475) );
AND2x2_ASAP7_75t_L g484 ( .A(n_12), .B(n_165), .Y(n_484) );
INVx2_ASAP7_75t_L g134 ( .A(n_13), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_14), .B(n_152), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_15), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g766 ( .A(n_15), .B(n_767), .C(n_769), .Y(n_766) );
AOI221x1_ASAP7_75t_L g187 ( .A1(n_16), .A2(n_137), .B1(n_188), .B2(n_190), .C(n_192), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_17), .B(n_143), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_18), .B(n_143), .Y(n_522) );
INVx1_ASAP7_75t_L g120 ( .A(n_19), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_20), .A2(n_92), .B1(n_143), .B2(n_175), .Y(n_463) );
AOI221xp5_ASAP7_75t_SL g136 ( .A1(n_21), .A2(n_38), .B1(n_137), .B2(n_143), .C(n_150), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_22), .A2(n_137), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_23), .B(n_154), .Y(n_203) );
OR2x2_ASAP7_75t_L g135 ( .A(n_24), .B(n_91), .Y(n_135) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_24), .A2(n_91), .B(n_134), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_25), .B(n_152), .Y(n_164) );
INVxp67_ASAP7_75t_L g186 ( .A(n_26), .Y(n_186) );
AND2x2_ASAP7_75t_L g236 ( .A(n_27), .B(n_132), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_28), .A2(n_137), .B(n_246), .Y(n_245) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_29), .A2(n_190), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_30), .B(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_31), .A2(n_137), .B(n_480), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_32), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_33), .B(n_152), .Y(n_517) );
AND2x2_ASAP7_75t_L g138 ( .A(n_34), .B(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g149 ( .A(n_34), .B(n_142), .Y(n_149) );
INVx1_ASAP7_75t_L g182 ( .A(n_34), .Y(n_182) );
OR2x6_ASAP7_75t_L g118 ( .A(n_35), .B(n_119), .Y(n_118) );
INVxp67_ASAP7_75t_L g769 ( .A(n_35), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_36), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_37), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_37), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_39), .B(n_143), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_40), .A2(n_84), .B1(n_137), .B2(n_180), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_41), .B(n_152), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_42), .B(n_143), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_43), .B(n_154), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_44), .A2(n_137), .B(n_471), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_45), .A2(n_74), .B1(n_739), .B2(n_740), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_45), .Y(n_739) );
AND2x2_ASAP7_75t_L g250 ( .A(n_46), .B(n_132), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_47), .B(n_154), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_48), .B(n_132), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_49), .B(n_143), .Y(n_534) );
INVx1_ASAP7_75t_L g141 ( .A(n_50), .Y(n_141) );
INVx1_ASAP7_75t_L g146 ( .A(n_50), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_51), .B(n_152), .Y(n_473) );
OAI22x1_ASAP7_75t_R g756 ( .A1(n_52), .A2(n_757), .B1(n_760), .B2(n_761), .Y(n_756) );
INVx1_ASAP7_75t_L g760 ( .A(n_52), .Y(n_760) );
AND2x2_ASAP7_75t_L g503 ( .A(n_53), .B(n_132), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_54), .B(n_143), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_55), .B(n_154), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_56), .B(n_154), .Y(n_516) );
AND2x2_ASAP7_75t_L g214 ( .A(n_57), .B(n_132), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_58), .B(n_143), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_59), .B(n_152), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_60), .B(n_143), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_61), .A2(n_137), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_62), .B(n_133), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_63), .B(n_154), .Y(n_211) );
AND2x2_ASAP7_75t_L g528 ( .A(n_64), .B(n_133), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_65), .A2(n_137), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_66), .B(n_152), .Y(n_204) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_67), .B(n_165), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_68), .B(n_154), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_69), .A2(n_72), .B1(n_758), .B2(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_69), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_70), .B(n_154), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_71), .A2(n_94), .B1(n_137), .B2(n_180), .Y(n_464) );
INVx1_ASAP7_75t_L g759 ( .A(n_72), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_73), .B(n_152), .Y(n_525) );
INVx1_ASAP7_75t_L g740 ( .A(n_74), .Y(n_740) );
INVx1_ASAP7_75t_L g139 ( .A(n_75), .Y(n_139) );
INVx1_ASAP7_75t_L g148 ( .A(n_75), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_76), .B(n_154), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_77), .A2(n_137), .B(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_78), .A2(n_137), .B(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_79), .A2(n_137), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g519 ( .A(n_80), .B(n_133), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_81), .B(n_132), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_82), .B(n_143), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_83), .A2(n_86), .B1(n_143), .B2(n_175), .Y(n_219) );
INVx1_ASAP7_75t_L g121 ( .A(n_85), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_87), .B(n_154), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_88), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g496 ( .A(n_89), .B(n_165), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_90), .A2(n_137), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_93), .B(n_152), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_95), .A2(n_137), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_96), .B(n_152), .Y(n_494) );
INVxp67_ASAP7_75t_L g189 ( .A(n_97), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_98), .B(n_143), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_99), .B(n_152), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_100), .A2(n_137), .B(n_162), .Y(n_161) );
BUFx2_ASAP7_75t_L g527 ( .A(n_101), .Y(n_527) );
BUFx2_ASAP7_75t_L g108 ( .A(n_102), .Y(n_108) );
INVx1_ASAP7_75t_SL g749 ( .A(n_102), .Y(n_749) );
AOI21xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_762), .B(n_770), .Y(n_103) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_123), .B(n_748), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AOI21xp33_ASAP7_75t_SL g750 ( .A1(n_110), .A2(n_751), .B(n_754), .Y(n_750) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_122), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_R g753 ( .A(n_115), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AND2x6_ASAP7_75t_SL g446 ( .A(n_116), .B(n_118), .Y(n_446) );
OR2x6_ASAP7_75t_SL g449 ( .A(n_116), .B(n_117), .Y(n_449) );
OR2x2_ASAP7_75t_L g746 ( .A(n_116), .B(n_118), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g765 ( .A(n_119), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
OAI222xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_734), .B1(n_735), .B2(n_741), .C1(n_744), .C2(n_747), .Y(n_123) );
OA22x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_443), .B1(n_447), .B2(n_450), .Y(n_124) );
OAI22x1_ASAP7_75t_L g754 ( .A1(n_125), .A2(n_126), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_126), .A2(n_447), .B1(n_451), .B2(n_743), .Y(n_742) );
OR2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_356), .Y(n_126) );
NAND3xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_266), .C(n_306), .Y(n_127) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_168), .B(n_195), .C(n_222), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_129), .B(n_271), .Y(n_305) );
NOR2x1p5_ASAP7_75t_L g129 ( .A(n_130), .B(n_157), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g241 ( .A(n_131), .Y(n_241) );
INVx2_ASAP7_75t_L g257 ( .A(n_131), .Y(n_257) );
OR2x2_ASAP7_75t_L g269 ( .A(n_131), .B(n_158), .Y(n_269) );
AND2x2_ASAP7_75t_L g283 ( .A(n_131), .B(n_242), .Y(n_283) );
INVx1_ASAP7_75t_L g311 ( .A(n_131), .Y(n_311) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_131), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_131), .B(n_158), .Y(n_417) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_136), .B(n_156), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_132), .Y(n_213) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_132), .A2(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_132), .A2(n_491), .B(n_492), .Y(n_490) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x4_ASAP7_75t_L g174 ( .A(n_134), .B(n_135), .Y(n_174) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
BUFx3_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
AND2x6_ASAP7_75t_L g154 ( .A(n_139), .B(n_145), .Y(n_154) );
INVx2_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
AND2x4_ASAP7_75t_L g180 ( .A(n_140), .B(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x4_ASAP7_75t_L g152 ( .A(n_141), .B(n_147), .Y(n_152) );
INVx2_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx5_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_153), .B(n_155), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_154), .B(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_155), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_155), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_155), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_155), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_155), .A2(n_247), .B(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_155), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_155), .A2(n_481), .B(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_155), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_155), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_155), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_155), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_155), .A2(n_537), .B(n_538), .Y(n_536) );
OR2x2_ASAP7_75t_L g238 ( .A(n_157), .B(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_157), .Y(n_373) );
AND2x2_ASAP7_75t_L g378 ( .A(n_157), .B(n_240), .Y(n_378) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g168 ( .A(n_158), .B(n_169), .Y(n_168) );
OR2x2_ASAP7_75t_L g237 ( .A(n_158), .B(n_170), .Y(n_237) );
OR2x2_ASAP7_75t_L g256 ( .A(n_158), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g285 ( .A(n_158), .Y(n_285) );
AND2x4_ASAP7_75t_SL g324 ( .A(n_158), .B(n_170), .Y(n_324) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_158), .Y(n_328) );
OR2x2_ASAP7_75t_L g345 ( .A(n_158), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g355 ( .A(n_158), .B(n_262), .Y(n_355) );
INVx1_ASAP7_75t_L g384 ( .A(n_158), .Y(n_384) );
OR2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_167), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_165), .Y(n_159) );
INVx2_ASAP7_75t_SL g217 ( .A(n_165), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_165), .A2(n_522), .B(n_523), .Y(n_521) );
BUFx4f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g191 ( .A(n_166), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_168), .B(n_313), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_169), .B(n_242), .Y(n_259) );
AND2x2_ASAP7_75t_L g271 ( .A(n_169), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g289 ( .A(n_169), .B(n_256), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_169), .B(n_310), .Y(n_309) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x4_ASAP7_75t_L g262 ( .A(n_170), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g284 ( .A(n_170), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g319 ( .A(n_170), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_170), .B(n_242), .Y(n_343) );
AND2x4_ASAP7_75t_L g170 ( .A(n_171), .B(n_187), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B1(n_180), .B2(n_185), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_174), .B(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_174), .B(n_189), .Y(n_188) );
NOR3xp33_ASAP7_75t_L g192 ( .A(n_174), .B(n_193), .C(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_174), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_174), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_174), .A2(n_534), .B(n_535), .Y(n_533) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_179), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
NOR2x1p5_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx3_ASAP7_75t_L g512 ( .A(n_190), .Y(n_512) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21x1_ASAP7_75t_L g243 ( .A1(n_191), .A2(n_244), .B(n_250), .Y(n_243) );
AO21x2_ASAP7_75t_L g468 ( .A1(n_191), .A2(n_469), .B(n_475), .Y(n_468) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_205), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_196), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g292 ( .A(n_196), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_196), .B(n_206), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g312 ( .A(n_196), .B(n_313), .C(n_314), .Y(n_312) );
AND2x2_ASAP7_75t_L g360 ( .A(n_196), .B(n_265), .Y(n_360) );
INVx5_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g227 ( .A(n_197), .B(n_228), .Y(n_227) );
AND2x4_ASAP7_75t_SL g264 ( .A(n_197), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
OR2x2_ASAP7_75t_L g303 ( .A(n_197), .B(n_293), .Y(n_303) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_197), .Y(n_320) );
AND2x2_ASAP7_75t_SL g338 ( .A(n_197), .B(n_226), .Y(n_338) );
AND2x4_ASAP7_75t_L g353 ( .A(n_197), .B(n_229), .Y(n_353) );
AND2x2_ASAP7_75t_L g367 ( .A(n_197), .B(n_206), .Y(n_367) );
OR2x2_ASAP7_75t_L g388 ( .A(n_197), .B(n_215), .Y(n_388) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
AND2x2_ASAP7_75t_L g442 ( .A(n_205), .B(n_320), .Y(n_442) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_215), .Y(n_205) );
AND2x4_ASAP7_75t_L g265 ( .A(n_206), .B(n_228), .Y(n_265) );
INVx2_ASAP7_75t_L g276 ( .A(n_206), .Y(n_276) );
AND2x2_ASAP7_75t_L g281 ( .A(n_206), .B(n_226), .Y(n_281) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_206), .Y(n_314) );
OR2x2_ASAP7_75t_L g337 ( .A(n_206), .B(n_229), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_206), .B(n_229), .Y(n_340) );
INVx1_ASAP7_75t_L g349 ( .A(n_206), .Y(n_349) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_213), .B(n_214), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_212), .Y(n_207) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_213), .A2(n_230), .B(n_236), .Y(n_229) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_213), .A2(n_230), .B(n_236), .Y(n_293) );
AOI21x1_ASAP7_75t_L g477 ( .A1(n_213), .A2(n_478), .B(n_484), .Y(n_477) );
AND2x2_ASAP7_75t_L g252 ( .A(n_215), .B(n_229), .Y(n_252) );
BUFx2_ASAP7_75t_L g301 ( .A(n_215), .Y(n_301) );
AND2x2_ASAP7_75t_L g396 ( .A(n_215), .B(n_276), .Y(n_396) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_216), .Y(n_226) );
AOI21x1_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_221), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
OAI221xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_237), .B1(n_238), .B2(n_251), .C(n_253), .Y(n_222) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
NOR2x1_ASAP7_75t_L g298 ( .A(n_225), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_225), .B(n_292), .Y(n_332) );
OR2x2_ASAP7_75t_L g344 ( .A(n_225), .B(n_340), .Y(n_344) );
OR2x2_ASAP7_75t_L g347 ( .A(n_225), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g436 ( .A(n_225), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g275 ( .A(n_226), .B(n_276), .Y(n_275) );
OA33x2_ASAP7_75t_L g308 ( .A1(n_226), .A2(n_269), .A3(n_309), .B1(n_312), .B2(n_315), .B3(n_318), .Y(n_308) );
OR2x2_ASAP7_75t_L g339 ( .A(n_226), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g363 ( .A(n_226), .B(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g371 ( .A(n_226), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g391 ( .A(n_226), .B(n_265), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_226), .B(n_280), .Y(n_429) );
INVx2_ASAP7_75t_L g299 ( .A(n_227), .Y(n_299) );
AOI322xp5_ASAP7_75t_L g369 ( .A1(n_227), .A2(n_282), .A3(n_370), .B1(n_373), .B2(n_374), .C1(n_376), .C2(n_378), .Y(n_369) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_229), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
OR2x2_ASAP7_75t_L g351 ( .A(n_237), .B(n_330), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_237), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g424 ( .A(n_237), .Y(n_424) );
INVx1_ASAP7_75t_SL g290 ( .A(n_238), .Y(n_290) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g323 ( .A(n_240), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g263 ( .A(n_242), .Y(n_263) );
INVx1_ASAP7_75t_L g272 ( .A(n_242), .Y(n_272) );
INVx1_ASAP7_75t_L g313 ( .A(n_242), .Y(n_313) );
OR2x2_ASAP7_75t_L g330 ( .A(n_242), .B(n_257), .Y(n_330) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_242), .Y(n_405) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_249), .Y(n_244) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_252), .B(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_SL g253 ( .A1(n_254), .A2(n_260), .B(n_264), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g327 ( .A1(n_254), .A2(n_328), .B(n_329), .C(n_331), .Y(n_327) );
AND2x4_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g392 ( .A(n_256), .B(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_257), .Y(n_261) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g416 ( .A(n_259), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AND2x2_ASAP7_75t_SL g385 ( .A(n_262), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g393 ( .A(n_262), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_262), .B(n_384), .Y(n_401) );
INVx3_ASAP7_75t_SL g326 ( .A(n_265), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_273), .B1(n_277), .B2(n_282), .C(n_286), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_272), .Y(n_317) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_275), .A2(n_302), .B(n_374), .Y(n_380) );
AND2x2_ASAP7_75t_L g406 ( .A(n_275), .B(n_353), .Y(n_406) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_276), .Y(n_294) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_280), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g415 ( .A(n_280), .B(n_337), .Y(n_415) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g364 ( .A(n_283), .Y(n_364) );
OAI21xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_291), .B(n_295), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx2_ASAP7_75t_L g437 ( .A(n_292), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_293), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g366 ( .A(n_293), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_294), .B(n_316), .Y(n_315) );
OAI31xp33_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_298), .A3(n_300), .B(n_304), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_299), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
OR2x2_ASAP7_75t_L g377 ( .A(n_301), .B(n_303), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_301), .B(n_353), .Y(n_432) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR5xp2_ASAP7_75t_L g306 ( .A(n_307), .B(n_321), .C(n_333), .D(n_342), .E(n_350), .Y(n_306) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_311), .B(n_313), .Y(n_346) );
INVx1_ASAP7_75t_L g386 ( .A(n_311), .Y(n_386) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_311), .Y(n_423) );
INVx1_ASAP7_75t_L g375 ( .A(n_314), .Y(n_375) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp33_ASAP7_75t_SL g318 ( .A(n_319), .B(n_320), .Y(n_318) );
OAI321xp33_ASAP7_75t_L g358 ( .A1(n_319), .A2(n_359), .A3(n_361), .B1(n_365), .B2(n_368), .C(n_369), .Y(n_358) );
INVx1_ASAP7_75t_L g412 ( .A(n_320), .Y(n_412) );
OAI21xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B(n_327), .Y(n_321) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_323), .A2(n_396), .B1(n_403), .B2(n_406), .Y(n_402) );
AND2x2_ASAP7_75t_L g431 ( .A(n_324), .B(n_405), .Y(n_431) );
INVx1_ASAP7_75t_L g341 ( .A(n_329), .Y(n_341) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_339), .B(n_341), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_340), .A2(n_351), .B1(n_352), .B2(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g413 ( .A(n_340), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_345), .B2(n_347), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_349), .B(n_353), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_351), .A2(n_428), .B1(n_430), .B2(n_432), .C(n_433), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_351), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_352), .A2(n_409), .B1(n_416), .B2(n_418), .C(n_419), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_354), .A2(n_380), .B(n_381), .Y(n_379) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_407), .Y(n_356) );
NOR3xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_379), .C(n_397), .Y(n_357) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_360), .Y(n_426) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g425 ( .A(n_368), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_370), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g418 ( .A(n_378), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_387), .B(n_389), .Y(n_381) );
INVxp67_ASAP7_75t_L g439 ( .A(n_382), .Y(n_439) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g394 ( .A(n_385), .Y(n_394) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B1(n_394), .B2(n_395), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI21xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_402), .Y(n_397) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g440 ( .A(n_403), .Y(n_440) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_427), .C(n_438), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_414), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_425), .B(n_426), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_424), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_431), .A2(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI21xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
CKINVDCx6p67_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx4_ASAP7_75t_SL g743 ( .A(n_444), .Y(n_743) );
INVx3_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_448), .Y(n_447) );
CKINVDCx11_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
INVx4_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x6_ASAP7_75t_L g451 ( .A(n_452), .B(n_671), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_587), .C(n_624), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_555), .C(n_570), .Y(n_453) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_500), .B1(n_529), .B2(n_541), .C(n_542), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_457), .B(n_485), .Y(n_456) );
OAI22xp33_ASAP7_75t_SL g615 ( .A1(n_457), .A2(n_579), .B1(n_616), .B2(n_619), .Y(n_615) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_465), .Y(n_457) );
OAI21xp33_ASAP7_75t_SL g625 ( .A1(n_458), .A2(n_626), .B(n_632), .Y(n_625) );
OR2x2_ASAP7_75t_L g654 ( .A(n_458), .B(n_487), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_458), .B(n_574), .Y(n_655) );
INVx2_ASAP7_75t_L g686 ( .A(n_458), .Y(n_686) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_459), .B(n_546), .Y(n_667) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g541 ( .A(n_460), .B(n_468), .Y(n_541) );
BUFx3_ASAP7_75t_L g567 ( .A(n_460), .Y(n_567) );
AND2x2_ASAP7_75t_L g703 ( .A(n_460), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g726 ( .A(n_460), .B(n_488), .Y(n_726) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AND2x4_ASAP7_75t_L g499 ( .A(n_461), .B(n_462), .Y(n_499) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_466), .B(n_488), .Y(n_646) );
INVx1_ASAP7_75t_L g683 ( .A(n_466), .Y(n_683) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_476), .Y(n_466) );
AND2x2_ASAP7_75t_L g498 ( .A(n_467), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g704 ( .A(n_467), .Y(n_704) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g547 ( .A(n_468), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_468), .B(n_476), .Y(n_548) );
AND2x2_ASAP7_75t_L g569 ( .A(n_468), .B(n_489), .Y(n_569) );
AND2x2_ASAP7_75t_L g651 ( .A(n_468), .B(n_477), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
AND2x4_ASAP7_75t_SL g544 ( .A(n_476), .B(n_489), .Y(n_544) );
INVx1_ASAP7_75t_L g575 ( .A(n_476), .Y(n_575) );
INVx2_ASAP7_75t_L g583 ( .A(n_476), .Y(n_583) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_476), .Y(n_607) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_477), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_498), .Y(n_485) );
AND2x2_ASAP7_75t_L g722 ( .A(n_486), .B(n_585), .Y(n_722) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_488), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g633 ( .A(n_488), .B(n_548), .Y(n_633) );
AND2x2_ASAP7_75t_L g650 ( .A(n_488), .B(n_651), .Y(n_650) );
INVx4_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x4_ASAP7_75t_L g574 ( .A(n_489), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g590 ( .A(n_489), .Y(n_590) );
AND2x2_ASAP7_75t_L g634 ( .A(n_489), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g641 ( .A(n_489), .B(n_642), .Y(n_641) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_489), .B(n_547), .Y(n_656) );
BUFx2_ASAP7_75t_L g666 ( .A(n_489), .Y(n_666) );
AND2x2_ASAP7_75t_L g691 ( .A(n_489), .B(n_651), .Y(n_691) );
AND2x2_ASAP7_75t_L g712 ( .A(n_489), .B(n_713), .Y(n_712) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_496), .Y(n_489) );
INVx1_ASAP7_75t_L g643 ( .A(n_497), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_498), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g673 ( .A(n_498), .B(n_544), .Y(n_673) );
INVx3_ASAP7_75t_L g580 ( .A(n_499), .Y(n_580) );
AND2x2_ASAP7_75t_L g713 ( .A(n_499), .B(n_635), .Y(n_713) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_501), .A2(n_543), .B1(n_548), .B2(n_549), .Y(n_542) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
INVx4_ASAP7_75t_L g540 ( .A(n_502), .Y(n_540) );
INVx2_ASAP7_75t_L g577 ( .A(n_502), .Y(n_577) );
NAND2x1_ASAP7_75t_L g603 ( .A(n_502), .B(n_520), .Y(n_603) );
OR2x2_ASAP7_75t_L g618 ( .A(n_502), .B(n_553), .Y(n_618) );
OR2x2_ASAP7_75t_SL g645 ( .A(n_502), .B(n_617), .Y(n_645) );
AND2x2_ASAP7_75t_L g658 ( .A(n_502), .B(n_532), .Y(n_658) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_502), .Y(n_679) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx2_ASAP7_75t_L g558 ( .A(n_510), .Y(n_558) );
AND2x2_ASAP7_75t_L g690 ( .A(n_510), .B(n_664), .Y(n_690) );
NOR2x1_ASAP7_75t_SL g510 ( .A(n_511), .B(n_520), .Y(n_510) );
AND2x2_ASAP7_75t_L g531 ( .A(n_511), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g707 ( .A(n_511), .B(n_630), .Y(n_707) );
AO21x1_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_511) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .Y(n_513) );
OR2x2_ASAP7_75t_L g539 ( .A(n_520), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g550 ( .A(n_520), .B(n_540), .Y(n_550) );
AND2x2_ASAP7_75t_L g596 ( .A(n_520), .B(n_553), .Y(n_596) );
OR2x2_ASAP7_75t_L g617 ( .A(n_520), .B(n_532), .Y(n_617) );
INVx2_ASAP7_75t_SL g623 ( .A(n_520), .Y(n_623) );
AND2x2_ASAP7_75t_L g629 ( .A(n_520), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g639 ( .A(n_520), .B(n_622), .Y(n_639) );
BUFx2_ASAP7_75t_L g661 ( .A(n_520), .Y(n_661) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_528), .Y(n_520) );
INVx2_ASAP7_75t_L g708 ( .A(n_529), .Y(n_708) );
OR2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_539), .Y(n_529) );
OR2x2_ASAP7_75t_L g733 ( .A(n_530), .B(n_577), .Y(n_733) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_531), .B(n_540), .Y(n_599) );
AND2x2_ASAP7_75t_L g670 ( .A(n_531), .B(n_550), .Y(n_670) );
INVx1_ASAP7_75t_L g552 ( .A(n_532), .Y(n_552) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_532), .Y(n_561) );
INVx1_ASAP7_75t_L g594 ( .A(n_532), .Y(n_594) );
INVx2_ASAP7_75t_L g630 ( .A(n_532), .Y(n_630) );
NOR2xp67_ASAP7_75t_L g560 ( .A(n_540), .B(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g620 ( .A(n_540), .Y(n_620) );
INVx2_ASAP7_75t_SL g696 ( .A(n_541), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_543), .A2(n_598), .B1(n_600), .B2(n_604), .Y(n_597) );
AND2x2_ASAP7_75t_SL g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x2_ASAP7_75t_L g724 ( .A(n_544), .B(n_580), .Y(n_724) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_546), .B(n_590), .Y(n_669) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g635 ( .A(n_547), .B(n_583), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_548), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g578 ( .A(n_549), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_549), .A2(n_693), .B1(n_697), .B2(n_699), .C(n_701), .Y(n_692) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x2_ASAP7_75t_L g562 ( .A(n_550), .B(n_563), .Y(n_562) );
INVxp67_ASAP7_75t_SL g586 ( .A(n_550), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_550), .B(n_593), .Y(n_648) );
INVx1_ASAP7_75t_SL g644 ( .A(n_551), .Y(n_644) );
AOI221xp5_ASAP7_75t_SL g672 ( .A1(n_551), .A2(n_562), .B1(n_673), .B2(n_674), .C(n_677), .Y(n_672) );
AOI322xp5_ASAP7_75t_L g705 ( .A1(n_551), .A2(n_623), .A3(n_650), .B1(n_706), .B2(n_708), .C1(n_709), .C2(n_712), .Y(n_705) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
BUFx2_ASAP7_75t_L g572 ( .A(n_552), .Y(n_572) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_553), .Y(n_564) );
INVx2_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
AND2x2_ASAP7_75t_L g663 ( .A(n_553), .B(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OA21x2_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_562), .B(n_565), .Y(n_555) );
AOI211xp5_ASAP7_75t_L g725 ( .A1(n_556), .A2(n_726), .B(n_727), .C(n_731), .Y(n_725) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OR2x2_ASAP7_75t_L g614 ( .A(n_558), .B(n_576), .Y(n_614) );
OR2x2_ASAP7_75t_L g698 ( .A(n_558), .B(n_593), .Y(n_698) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g638 ( .A(n_560), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g716 ( .A(n_563), .Y(n_716) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g602 ( .A(n_564), .Y(n_602) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
OR2x2_ASAP7_75t_L g571 ( .A(n_567), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g606 ( .A(n_569), .B(n_607), .Y(n_606) );
OAI322xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .A3(n_576), .B1(n_578), .B2(n_579), .C1(n_584), .C2(n_586), .Y(n_570) );
INVx1_ASAP7_75t_L g612 ( .A(n_571), .Y(n_612) );
OR2x2_ASAP7_75t_L g584 ( .A(n_573), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_573), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g595 ( .A(n_577), .B(n_596), .Y(n_595) );
OAI32xp33_ASAP7_75t_L g640 ( .A1(n_577), .A2(n_641), .A3(n_644), .B1(n_645), .B2(n_646), .Y(n_640) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx2_ASAP7_75t_L g585 ( .A(n_580), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_580), .B(n_643), .Y(n_642) );
NOR2x1_ASAP7_75t_L g682 ( .A(n_580), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g706 ( .A(n_580), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g627 ( .A(n_581), .Y(n_627) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_585), .B(n_651), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_608), .Y(n_587) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B(n_597), .Y(n_588) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g657 ( .A(n_596), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_599), .A2(n_619), .B1(n_721), .B2(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_601), .A2(n_648), .B(n_649), .C(n_652), .Y(n_647) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx3_ASAP7_75t_L g729 ( .A(n_603), .Y(n_729) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g610 ( .A(n_607), .Y(n_610) );
AO21x1_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_611), .B(n_615), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g675 ( .A(n_610), .Y(n_675) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_616), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g631 ( .A(n_618), .Y(n_631) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g688 ( .A(n_621), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_647), .C(n_659), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OAI21xp5_ASAP7_75t_SL g689 ( .A1(n_628), .A2(n_690), .B(n_691), .Y(n_689) );
AND2x4_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g664 ( .A(n_630), .Y(n_664) );
O2A1O1Ixp5_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_634), .B(n_636), .C(n_640), .Y(n_632) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_642), .Y(n_732) );
INVx2_ASAP7_75t_L g717 ( .A(n_645), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_646), .A2(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g711 ( .A(n_651), .Y(n_711) );
OAI31xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .A3(n_656), .B(n_657), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g730 ( .A(n_658), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_665), .B(n_668), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
BUFx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g680 ( .A(n_663), .Y(n_680) );
AOI21xp33_ASAP7_75t_SL g727 ( .A1(n_665), .A2(n_728), .B(n_730), .Y(n_727) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx2_ASAP7_75t_L g695 ( .A(n_666), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_666), .B(n_686), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_666), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g676 ( .A(n_667), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
NAND5xp2_ASAP7_75t_L g671 ( .A(n_672), .B(n_692), .C(n_705), .D(n_714), .E(n_725), .Y(n_671) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_681), .B1(n_684), .B2(n_687), .C(n_689), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVxp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_718), .B(n_720), .Y(n_714) );
AND2x4_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g761 ( .A(n_757), .Y(n_761) );
INVx3_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g772 ( .A(n_763), .Y(n_772) );
INVx2_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_SL g764 ( .A(n_765), .B(n_766), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
endmodule