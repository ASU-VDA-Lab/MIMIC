module fake_aes_1408_n_697 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_697);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_697;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g78 ( .A(n_31), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_39), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_77), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_67), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_5), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_36), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_17), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
NOR2xp33_ASAP7_75t_L g86 ( .A(n_52), .B(n_28), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_73), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_65), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_63), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_25), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_10), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_34), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_58), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_41), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_57), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_15), .Y(n_96) );
INVx2_ASAP7_75t_SL g97 ( .A(n_50), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_62), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_23), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_35), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_54), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_47), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_45), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_13), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_29), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_48), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_68), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_74), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_66), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_14), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
BUFx10_ASAP7_75t_L g113 ( .A(n_27), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_59), .Y(n_115) );
BUFx10_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_44), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_76), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_30), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_69), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_49), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_51), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_15), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_38), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_3), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_108), .B(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_125), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_108), .Y(n_131) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_78), .A2(n_75), .B(n_72), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_125), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_118), .B(n_0), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_118), .B(n_1), .Y(n_136) );
NAND2xp33_ASAP7_75t_SL g137 ( .A(n_80), .B(n_1), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_102), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_97), .B(n_2), .Y(n_139) );
CKINVDCx8_ASAP7_75t_R g140 ( .A(n_101), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_107), .Y(n_143) );
NAND2xp33_ASAP7_75t_L g144 ( .A(n_90), .B(n_70), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_97), .B(n_2), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_103), .B(n_3), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_81), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_104), .B(n_4), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_83), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_115), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_113), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_124), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_116), .B(n_4), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_125), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_83), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_125), .Y(n_159) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_85), .A2(n_21), .B(n_61), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_85), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_87), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_87), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_88), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_88), .Y(n_165) );
INVxp67_ASAP7_75t_L g166 ( .A(n_116), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_116), .B(n_5), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_89), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_131), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_135), .B(n_109), .Y(n_172) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_135), .B(n_109), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_135), .B(n_91), .Y(n_174) );
AO22x2_ASAP7_75t_L g175 ( .A1(n_135), .A2(n_95), .B1(n_99), .B2(n_122), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_131), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
INVx8_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_139), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_130), .Y(n_182) );
INVx5_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_127), .Y(n_184) );
OAI221xp5_ASAP7_75t_L g185 ( .A1(n_128), .A2(n_123), .B1(n_96), .B2(n_114), .C(n_111), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_126), .Y(n_186) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_127), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_152), .B(n_91), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_144), .B(n_95), .Y(n_190) );
INVxp67_ASAP7_75t_SL g191 ( .A(n_128), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_152), .B(n_113), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_152), .B(n_106), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_157), .B(n_123), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_157), .B(n_92), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_130), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_157), .B(n_94), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_158), .Y(n_201) );
AO22x1_ASAP7_75t_L g202 ( .A1(n_154), .A2(n_93), .B1(n_119), .B2(n_121), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_132), .Y(n_204) );
INVx6_ASAP7_75t_L g205 ( .A(n_130), .Y(n_205) );
AND2x6_ASAP7_75t_L g206 ( .A(n_154), .B(n_100), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_167), .B(n_84), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_167), .B(n_84), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_163), .Y(n_209) );
BUFx10_ASAP7_75t_L g210 ( .A(n_129), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_132), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_163), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_126), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_129), .B(n_90), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_141), .B(n_99), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_136), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_140), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_165), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_141), .B(n_92), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_134), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_147), .B(n_96), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_165), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_140), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_134), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_166), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_147), .B(n_112), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_165), .Y(n_228) );
AND2x2_ASAP7_75t_SL g229 ( .A(n_136), .B(n_89), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_134), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_173), .A2(n_168), .B1(n_164), .B2(n_162), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_191), .B(n_217), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_210), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_177), .B(n_168), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_180), .B(n_162), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_210), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_179), .Y(n_238) );
INVx5_ASAP7_75t_L g239 ( .A(n_210), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_181), .B(n_164), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_179), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_192), .B(n_161), .Y(n_242) );
OR2x6_ASAP7_75t_L g243 ( .A(n_172), .B(n_114), .Y(n_243) );
INVx4_ASAP7_75t_L g244 ( .A(n_178), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_196), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_213), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_213), .Y(n_247) );
BUFx4f_ASAP7_75t_L g248 ( .A(n_172), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_223), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_223), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_228), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_188), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_228), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_193), .Y(n_254) );
AND2x6_ASAP7_75t_L g255 ( .A(n_212), .B(n_98), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_215), .B(n_161), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_171), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_201), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_209), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_173), .A2(n_149), .B1(n_146), .B2(n_148), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_176), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_220), .B(n_149), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_211), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_219), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_207), .B(n_138), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_230), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_178), .Y(n_267) );
OR2x4_ASAP7_75t_L g268 ( .A(n_195), .B(n_105), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_218), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_184), .B(n_117), .Y(n_270) );
BUFx8_ASAP7_75t_L g271 ( .A(n_206), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_230), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_212), .Y(n_273) );
NAND3xp33_ASAP7_75t_SL g274 ( .A(n_218), .B(n_82), .C(n_117), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_206), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_194), .B(n_197), .Y(n_276) );
AND3x1_ASAP7_75t_SL g277 ( .A(n_185), .B(n_98), .C(n_100), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_196), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_194), .B(n_138), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_171), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_229), .B(n_138), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_226), .B(n_110), .Y(n_282) );
AND2x4_ASAP7_75t_SL g283 ( .A(n_196), .B(n_125), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_178), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_229), .B(n_142), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_171), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_207), .B(n_143), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_197), .B(n_142), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_197), .B(n_142), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_178), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_184), .B(n_187), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_169), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_169), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_206), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_169), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_175), .A2(n_137), .B1(n_143), .B2(n_156), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_233), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_239), .B(n_184), .Y(n_298) );
OAI22xp33_ASAP7_75t_L g299 ( .A1(n_243), .A2(n_224), .B1(n_172), .B2(n_187), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_231), .A2(n_208), .B(n_198), .C(n_227), .Y(n_300) );
OR2x6_ASAP7_75t_L g301 ( .A(n_243), .B(n_175), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_269), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_280), .A2(n_187), .B(n_171), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_243), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_238), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_247), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_234), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_236), .A2(n_174), .B(n_222), .C(n_200), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_243), .A2(n_175), .B1(n_206), .B2(n_190), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_247), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_234), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_251), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_235), .A2(n_174), .B(n_222), .C(n_208), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_232), .B(n_206), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_239), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_244), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_269), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
AOI21x1_ASAP7_75t_L g320 ( .A1(n_280), .A2(n_175), .B(n_160), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_244), .B(n_222), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_271), .Y(n_322) );
INVx4_ASAP7_75t_L g323 ( .A(n_244), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_240), .B(n_174), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_241), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_251), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_237), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_242), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_241), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_248), .A2(n_190), .B1(n_224), .B2(n_188), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_253), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_265), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_276), .B(n_206), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_237), .Y(n_334) );
NOR2xp67_ASAP7_75t_SL g335 ( .A(n_239), .B(n_204), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_246), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_256), .A2(n_225), .B(n_221), .C(n_214), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_253), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_248), .A2(n_188), .B1(n_171), .B2(n_204), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_239), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_239), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_248), .A2(n_204), .B1(n_221), .B2(n_186), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_246), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_237), .Y(n_344) );
BUFx12f_ASAP7_75t_L g345 ( .A(n_271), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_237), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_249), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_328), .Y(n_348) );
NOR2xp67_ASAP7_75t_L g349 ( .A(n_303), .B(n_274), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_319), .A2(n_282), .B1(n_260), .B2(n_296), .C(n_262), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_301), .A2(n_276), .B1(n_271), .B2(n_275), .Y(n_351) );
CKINVDCx12_ASAP7_75t_R g352 ( .A(n_301), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_316), .Y(n_353) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_305), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_317), .B(n_276), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_332), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_310), .A2(n_275), .B1(n_294), .B2(n_267), .Y(n_357) );
OR2x6_ASAP7_75t_L g358 ( .A(n_301), .B(n_294), .Y(n_358) );
NOR2xp67_ASAP7_75t_SL g359 ( .A(n_327), .B(n_237), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
BUFx12f_ASAP7_75t_L g361 ( .A(n_303), .Y(n_361) );
INVx6_ASAP7_75t_L g362 ( .A(n_317), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_321), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_301), .B(n_265), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_333), .A2(n_252), .B1(n_216), .B2(n_287), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_297), .A2(n_255), .B1(n_287), .B2(n_284), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_317), .B(n_284), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_302), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_337), .A2(n_273), .B(n_249), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_304), .A2(n_273), .B(n_286), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_333), .A2(n_216), .B1(n_285), .B2(n_281), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_318), .B(n_202), .Y(n_372) );
OR2x6_ASAP7_75t_L g373 ( .A(n_323), .B(n_267), .Y(n_373) );
NOR2x1_ASAP7_75t_SL g374 ( .A(n_323), .B(n_345), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_333), .A2(n_216), .B1(n_254), .B2(n_263), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_306), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_324), .B(n_268), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_306), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_307), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_362), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_379), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_358), .A2(n_299), .B1(n_343), .B2(n_347), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_350), .A2(n_297), .B1(n_324), .B2(n_318), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_364), .B(n_343), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_372), .B(n_330), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_374), .A2(n_345), .B1(n_322), .B2(n_321), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g387 ( .A1(n_377), .A2(n_309), .B1(n_314), .B2(n_300), .C(n_315), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_372), .A2(n_321), .B1(n_325), .B2(n_329), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_364), .A2(n_325), .B1(n_329), .B2(n_336), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_352), .A2(n_277), .B1(n_268), .B2(n_336), .Y(n_390) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_369), .A2(n_320), .B(n_339), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_366), .A2(n_347), .B1(n_268), .B2(n_311), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_362), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_348), .A2(n_216), .B1(n_323), .B2(n_279), .Y(n_394) );
AOI332xp33_ASAP7_75t_L g395 ( .A1(n_356), .A2(n_150), .A3(n_156), .B1(n_153), .B2(n_151), .B3(n_143), .C1(n_120), .C2(n_121), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_360), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_352), .A2(n_255), .B1(n_313), .B2(n_307), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_358), .A2(n_313), .B1(n_326), .B2(n_338), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_368), .B(n_311), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_363), .A2(n_202), .B1(n_288), .B2(n_289), .C(n_263), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_376), .A2(n_378), .B1(n_355), .B2(n_354), .C(n_351), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_362), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_355), .A2(n_216), .B1(n_322), .B2(n_255), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_355), .A2(n_216), .B1(n_255), .B2(n_270), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_367), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_358), .A2(n_255), .B1(n_264), .B2(n_254), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_390), .A2(n_358), .B1(n_373), .B2(n_349), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_406), .B(n_353), .Y(n_409) );
OR2x2_ASAP7_75t_SL g410 ( .A(n_393), .B(n_362), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_383), .B(n_86), .C(n_153), .Y(n_411) );
OAI31xp33_ASAP7_75t_L g412 ( .A1(n_392), .A2(n_367), .A3(n_357), .B(n_365), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_384), .B(n_353), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_396), .Y(n_414) );
OA21x2_ASAP7_75t_L g415 ( .A1(n_382), .A2(n_370), .B(n_286), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_406), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_384), .B(n_326), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_399), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_399), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_385), .A2(n_373), .B1(n_361), .B2(n_312), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_382), .A2(n_373), .B1(n_255), .B2(n_361), .Y(n_423) );
NAND3xp33_ASAP7_75t_SL g424 ( .A(n_395), .B(n_367), .C(n_375), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_406), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_388), .B(n_331), .Y(n_426) );
OR2x6_ASAP7_75t_L g427 ( .A(n_398), .B(n_373), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_390), .B(n_153), .C(n_151), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_403), .B(n_341), .Y(n_429) );
OA21x2_ASAP7_75t_L g430 ( .A1(n_381), .A2(n_320), .B(n_156), .Y(n_430) );
AOI31xp33_ASAP7_75t_L g431 ( .A1(n_386), .A2(n_401), .A3(n_397), .B(n_407), .Y(n_431) );
NOR2x1_ASAP7_75t_SL g432 ( .A(n_393), .B(n_312), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_387), .A2(n_151), .B1(n_150), .B2(n_264), .C(n_250), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_400), .A2(n_371), .B1(n_221), .B2(n_225), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_402), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_403), .B(n_341), .Y(n_437) );
OAI211xp5_ASAP7_75t_SL g438 ( .A1(n_389), .A2(n_120), .B(n_122), .C(n_150), .Y(n_438) );
AOI322xp5_ASAP7_75t_L g439 ( .A1(n_395), .A2(n_186), .A3(n_225), .B1(n_214), .B2(n_9), .C1(n_10), .C2(n_11), .Y(n_439) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_397), .A2(n_338), .B(n_331), .Y(n_440) );
AOI33xp33_ASAP7_75t_L g441 ( .A1(n_394), .A2(n_292), .A3(n_293), .B1(n_295), .B2(n_250), .B3(n_259), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_380), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_425), .Y(n_443) );
NOR2x1p5_ASAP7_75t_L g444 ( .A(n_424), .B(n_393), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_436), .B(n_391), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_422), .B(n_380), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_436), .B(n_391), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_430), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_424), .A2(n_393), .B1(n_404), .B2(n_391), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_430), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_427), .A2(n_393), .B1(n_316), .B2(n_340), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_414), .B(n_160), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_417), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_421), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_411), .B(n_130), .C(n_159), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_433), .B(n_160), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_439), .A2(n_405), .B(n_308), .C(n_340), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_419), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_413), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_420), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_442), .B(n_6), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_418), .B(n_6), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_415), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_415), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_408), .B(n_186), .C(n_214), .Y(n_465) );
INVx5_ASAP7_75t_SL g466 ( .A(n_427), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_412), .A2(n_423), .B1(n_427), .B2(n_438), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_431), .A2(n_259), .B1(n_258), .B2(n_292), .C(n_293), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_416), .B(n_7), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_440), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_440), .Y(n_471) );
AOI33xp33_ASAP7_75t_L g472 ( .A1(n_435), .A2(n_295), .A3(n_8), .B1(n_9), .B2(n_11), .B3(n_12), .Y(n_472) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_426), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_410), .B(n_258), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_432), .B(n_327), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_431), .A2(n_308), .B1(n_342), .B2(n_204), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_441), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_438), .A2(n_308), .B1(n_204), .B2(n_203), .Y(n_478) );
AOI31xp33_ASAP7_75t_L g479 ( .A1(n_409), .A2(n_298), .A3(n_359), .B(n_291), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_429), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_428), .B(n_7), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_437), .B(n_8), .Y(n_482) );
OAI33xp33_ASAP7_75t_L g483 ( .A1(n_434), .A2(n_12), .A3(n_13), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_483) );
INVxp67_ASAP7_75t_L g484 ( .A(n_429), .Y(n_484) );
OAI31xp33_ASAP7_75t_SL g485 ( .A1(n_437), .A2(n_18), .A3(n_19), .B(n_20), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_434), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_414), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_430), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_436), .Y(n_489) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_439), .B(n_203), .C(n_19), .D(n_20), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_430), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_410), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_445), .B(n_159), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_482), .B(n_22), .Y(n_494) );
NAND4xp25_ASAP7_75t_L g495 ( .A(n_485), .B(n_203), .C(n_189), .D(n_199), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_443), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_453), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_490), .A2(n_344), .B(n_335), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_476), .A2(n_334), .B(n_346), .Y(n_499) );
NOR3xp33_ASAP7_75t_SL g500 ( .A(n_490), .B(n_24), .C(n_26), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_453), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_473), .B(n_133), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_445), .B(n_159), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_448), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_448), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_482), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_467), .A2(n_159), .B1(n_155), .B2(n_133), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_487), .Y(n_508) );
OAI33xp33_ASAP7_75t_L g509 ( .A1(n_477), .A2(n_189), .A3(n_199), .B1(n_182), .B2(n_159), .B3(n_155), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_448), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_489), .B(n_159), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_487), .Y(n_512) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_444), .B(n_359), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_458), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_447), .B(n_155), .Y(n_515) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_444), .B(n_335), .Y(n_516) );
NAND2x1_ASAP7_75t_L g517 ( .A(n_450), .B(n_346), .Y(n_517) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_483), .B(n_182), .C(n_344), .Y(n_518) );
NOR2xp33_ASAP7_75t_SL g519 ( .A(n_443), .B(n_346), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_447), .B(n_155), .Y(n_520) );
NOR2x1p5_ASAP7_75t_L g521 ( .A(n_485), .B(n_155), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_450), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_458), .B(n_155), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_454), .Y(n_524) );
NOR2x1_ASAP7_75t_L g525 ( .A(n_474), .B(n_344), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_460), .B(n_133), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_460), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_459), .B(n_133), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_461), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_475), .B(n_346), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_450), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_488), .B(n_133), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_461), .B(n_133), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_488), .B(n_32), .Y(n_534) );
BUFx2_ASAP7_75t_L g535 ( .A(n_480), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_488), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_477), .A2(n_283), .B1(n_266), .B2(n_272), .C(n_183), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_462), .B(n_346), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_491), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_491), .Y(n_540) );
BUFx2_ASAP7_75t_L g541 ( .A(n_480), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_462), .Y(n_542) );
BUFx3_ASAP7_75t_L g543 ( .A(n_475), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_484), .B(n_334), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_491), .B(n_37), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_492), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_466), .B(n_40), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_464), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_466), .B(n_334), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_466), .B(n_42), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_463), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_524), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_524), .B(n_446), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_493), .B(n_470), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_542), .B(n_466), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_512), .Y(n_556) );
NOR2xp67_ASAP7_75t_L g557 ( .A(n_495), .B(n_522), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_529), .B(n_492), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_496), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_514), .B(n_468), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_506), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_535), .B(n_466), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_543), .B(n_471), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_512), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_493), .B(n_471), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_514), .B(n_468), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_497), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_551), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_535), .B(n_474), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_527), .B(n_469), .Y(n_570) );
AOI322xp5_ASAP7_75t_L g571 ( .A1(n_500), .A2(n_469), .A3(n_486), .B1(n_449), .B2(n_451), .C1(n_452), .C2(n_464), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_528), .B(n_472), .C(n_476), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_501), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_546), .B(n_486), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_508), .Y(n_575) );
NOR2x1p5_ASAP7_75t_L g576 ( .A(n_496), .B(n_481), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_519), .B(n_475), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_503), .B(n_452), .Y(n_578) );
NOR2x1p5_ASAP7_75t_L g579 ( .A(n_521), .B(n_481), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_503), .B(n_470), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_528), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_515), .B(n_456), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_511), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_511), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_509), .A2(n_455), .B(n_475), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_515), .B(n_471), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_522), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_520), .B(n_470), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_543), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_520), .B(n_456), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_548), .B(n_463), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_523), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_548), .B(n_463), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_541), .B(n_457), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_541), .B(n_465), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_523), .B(n_478), .Y(n_596) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_522), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_502), .B(n_479), .Y(n_598) );
AND3x2_ASAP7_75t_L g599 ( .A(n_547), .B(n_479), .C(n_455), .Y(n_599) );
NOR2xp67_ASAP7_75t_L g600 ( .A(n_536), .B(n_43), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_526), .B(n_46), .Y(n_601) );
NAND3xp33_ASAP7_75t_SL g602 ( .A(n_494), .B(n_53), .C(n_55), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_526), .B(n_183), .C(n_327), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_567), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_573), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_552), .B(n_502), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_575), .Y(n_607) );
OAI31xp33_ASAP7_75t_SL g608 ( .A1(n_561), .A2(n_550), .A3(n_547), .B(n_525), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_556), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_587), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_574), .B(n_526), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_564), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_553), .B(n_574), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_583), .B(n_539), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_557), .A2(n_513), .B1(n_516), .B2(n_549), .Y(n_615) );
XNOR2xp5_ASAP7_75t_L g616 ( .A(n_579), .B(n_550), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_584), .Y(n_617) );
OAI21xp5_ASAP7_75t_SL g618 ( .A1(n_599), .A2(n_571), .B(n_572), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_581), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_554), .B(n_540), .Y(n_620) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_587), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_578), .B(n_539), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_570), .B(n_540), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_589), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_558), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_598), .A2(n_513), .B1(n_516), .B2(n_545), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_591), .B(n_540), .Y(n_627) );
OAI32xp33_ASAP7_75t_L g628 ( .A1(n_559), .A2(n_516), .A3(n_513), .B1(n_549), .B2(n_538), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_568), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_594), .A2(n_533), .B1(n_507), .B2(n_498), .C(n_518), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_582), .B(n_551), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_568), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_555), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_560), .B(n_544), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_591), .B(n_593), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_566), .A2(n_499), .B1(n_537), .B2(n_536), .C(n_504), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_593), .B(n_536), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_592), .B(n_504), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_554), .B(n_505), .Y(n_639) );
XOR2xp5_ASAP7_75t_SL g640 ( .A(n_562), .B(n_545), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_590), .B(n_531), .Y(n_641) );
XOR2x2_ASAP7_75t_L g642 ( .A(n_599), .B(n_530), .Y(n_642) );
XOR2x2_ASAP7_75t_L g643 ( .A(n_577), .B(n_530), .Y(n_643) );
AOI221x1_ASAP7_75t_L g644 ( .A1(n_585), .A2(n_532), .B1(n_534), .B2(n_531), .C(n_505), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_569), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_576), .A2(n_510), .B1(n_534), .B2(n_530), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_595), .A2(n_532), .B(n_510), .C(n_517), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_577), .A2(n_517), .B1(n_283), .B2(n_327), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_602), .B(n_266), .C(n_272), .Y(n_649) );
NOR2xp67_ASAP7_75t_L g650 ( .A(n_603), .B(n_56), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_565), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_565), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_580), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_580), .B(n_64), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_586), .B(n_588), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_586), .Y(n_656) );
NAND2xp33_ASAP7_75t_L g657 ( .A(n_588), .B(n_334), .Y(n_657) );
AOI321xp33_ASAP7_75t_L g658 ( .A1(n_597), .A2(n_278), .A3(n_245), .B1(n_205), .B2(n_257), .C(n_183), .Y(n_658) );
XNOR2x1_ASAP7_75t_L g659 ( .A(n_563), .B(n_334), .Y(n_659) );
NAND4xp25_ASAP7_75t_SL g660 ( .A(n_601), .B(n_327), .C(n_290), .D(n_257), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_563), .B(n_257), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_596), .A2(n_183), .B1(n_257), .B2(n_245), .C(n_278), .Y(n_662) );
XNOR2xp5_ASAP7_75t_L g663 ( .A(n_616), .B(n_642), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_624), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_617), .B(n_619), .Y(n_665) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_618), .A2(n_608), .B1(n_616), .B2(n_626), .C(n_613), .Y(n_666) );
AOI22x1_ASAP7_75t_L g667 ( .A1(n_658), .A2(n_621), .B1(n_610), .B2(n_633), .Y(n_667) );
OA22x2_ASAP7_75t_L g668 ( .A1(n_646), .A2(n_625), .B1(n_644), .B2(n_645), .Y(n_668) );
OAI211xp5_ASAP7_75t_L g669 ( .A1(n_628), .A2(n_630), .B(n_634), .C(n_658), .Y(n_669) );
NOR4xp25_ASAP7_75t_SL g670 ( .A(n_636), .B(n_605), .C(n_604), .D(n_607), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_646), .A2(n_615), .B1(n_656), .B2(n_611), .Y(n_671) );
XNOR2xp5_ASAP7_75t_L g672 ( .A(n_643), .B(n_640), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_622), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_647), .A2(n_650), .B(n_648), .Y(n_674) );
AOI321xp33_ASAP7_75t_L g675 ( .A1(n_613), .A2(n_634), .A3(n_628), .B1(n_606), .B2(n_623), .C(n_620), .Y(n_675) );
NOR2xp67_ASAP7_75t_L g676 ( .A(n_648), .B(n_660), .Y(n_676) );
OR3x2_ASAP7_75t_L g677 ( .A(n_666), .B(n_654), .C(n_622), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_673), .Y(n_678) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_669), .B(n_600), .Y(n_679) );
OAI21xp33_ASAP7_75t_SL g680 ( .A1(n_668), .A2(n_659), .B(n_655), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_663), .B(n_652), .Y(n_681) );
AOI32xp33_ASAP7_75t_L g682 ( .A1(n_671), .A2(n_657), .A3(n_620), .B1(n_639), .B2(n_651), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_664), .A2(n_649), .B(n_612), .C(n_609), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_667), .A2(n_662), .B(n_614), .C(n_627), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_680), .A2(n_675), .B1(n_672), .B2(n_668), .C(n_674), .Y(n_685) );
AOI22xp5_ASAP7_75t_SL g686 ( .A1(n_681), .A2(n_664), .B1(n_670), .B2(n_665), .Y(n_686) );
NAND3xp33_ASAP7_75t_SL g687 ( .A(n_682), .B(n_676), .C(n_631), .Y(n_687) );
OAI22xp5_ASAP7_75t_SL g688 ( .A1(n_679), .A2(n_665), .B1(n_653), .B2(n_635), .Y(n_688) );
AND3x4_ASAP7_75t_L g689 ( .A(n_685), .B(n_677), .C(n_684), .Y(n_689) );
OR4x2_ASAP7_75t_L g690 ( .A(n_687), .B(n_683), .C(n_678), .D(n_631), .Y(n_690) );
AOI22x1_ASAP7_75t_L g691 ( .A1(n_686), .A2(n_641), .B1(n_629), .B2(n_632), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_689), .A2(n_688), .B1(n_563), .B2(n_629), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_691), .A2(n_637), .B1(n_638), .B2(n_632), .Y(n_693) );
INVx4_ASAP7_75t_L g694 ( .A(n_692), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_694), .A2(n_693), .B(n_690), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_695), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_696), .A2(n_661), .B1(n_639), .B2(n_290), .C(n_183), .Y(n_697) );
endmodule