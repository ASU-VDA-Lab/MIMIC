module fake_jpeg_22874_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_38),
.Y(n_45)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_20),
.B1(n_16),
.B2(n_22),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_53),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_58),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_17),
.Y(n_53)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_16),
.B1(n_22),
.B2(n_26),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_31),
.B1(n_32),
.B2(n_26),
.Y(n_82)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_34),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_80),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_46),
.Y(n_107)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_23),
.A3(n_30),
.B1(n_18),
.B2(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_48),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_27),
.B1(n_60),
.B2(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_66),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_46),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_42),
.B1(n_27),
.B2(n_26),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_42),
.B1(n_60),
.B2(n_51),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_47),
.B(n_52),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_55),
.B(n_43),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_92),
.B1(n_75),
.B2(n_67),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_93),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_95),
.B1(n_105),
.B2(n_50),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_45),
.B1(n_49),
.B2(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_51),
.B1(n_60),
.B2(n_36),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_56),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_48),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_73),
.C(n_77),
.Y(n_109)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_39),
.B1(n_43),
.B2(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_57),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_78),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_124),
.C(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_116),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_77),
.B(n_81),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_118),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_91),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_125),
.Y(n_141)
);

XOR2x1_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_94),
.B(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_85),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_117),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_132),
.B1(n_133),
.B2(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_103),
.B1(n_124),
.B2(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_90),
.B1(n_107),
.B2(n_95),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_139),
.C(n_147),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_137),
.B(n_142),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_106),
.B1(n_75),
.B2(n_102),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_83),
.C(n_66),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_120),
.Y(n_144)
);

INVxp33_ASAP7_75t_SL g152 ( 
.A(n_144),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_39),
.B1(n_18),
.B2(n_23),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_114),
.B1(n_135),
.B2(n_127),
.Y(n_158)
);

AO221x1_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_99),
.B1(n_33),
.B2(n_25),
.C(n_24),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_30),
.C(n_28),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

FAx1_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_118),
.CI(n_114),
.CON(n_154),
.SN(n_154)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_19),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_110),
.C(n_125),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_149),
.C(n_154),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_24),
.B1(n_25),
.B2(n_15),
.Y(n_171)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_112),
.B(n_111),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_136),
.B1(n_141),
.B2(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

AOI321xp33_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_141),
.A3(n_134),
.B1(n_139),
.B2(n_147),
.C(n_117),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_171),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_24),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_173),
.C(n_152),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_15),
.C(n_14),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_174),
.A2(n_159),
.B1(n_162),
.B2(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_179),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_171),
.B1(n_166),
.B2(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_159),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_182),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_170),
.A2(n_148),
.B(n_149),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_162),
.C(n_157),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_3),
.C(n_4),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_181),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_163),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_190),
.C(n_8),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_189),
.C(n_10),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_164),
.B1(n_173),
.B2(n_14),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_191),
.B(n_192),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_180),
.B1(n_13),
.B2(n_12),
.Y(n_192)
);

OAI221xp5_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_5),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_196),
.C(n_190),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_186),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_8),
.C(n_9),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_199),
.B(n_202),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_10),
.C(n_195),
.Y(n_205)
);


endmodule