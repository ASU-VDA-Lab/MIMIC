module fake_jpeg_20177_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVxp67_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVxp33_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_17),
.Y(n_25)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_9),
.B(n_8),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_10),
.B1(n_14),
.B2(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_8),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_17),
.B1(n_23),
.B2(n_11),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_33),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_16),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_11),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_16),
.C(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

OA21x2_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_28),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_7),
.Y(n_44)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_34),
.C(n_35),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_46),
.C(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_48),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_49),
.B(n_47),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_53),
.B(n_6),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_42),
.B(n_6),
.C(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

AOI321xp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_55),
.C(n_49),
.Y(n_57)
);

BUFx24_ASAP7_75t_SL g58 ( 
.A(n_57),
.Y(n_58)
);


endmodule