module fake_jpeg_17978_n_32 (n_3, n_2, n_1, n_0, n_4, n_5, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_32;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

AOI22xp33_ASAP7_75t_L g11 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_11),
.A2(n_9),
.B1(n_5),
.B2(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_0),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_14),
.C(n_9),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_6),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_16),
.B1(n_8),
.B2(n_4),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_8),
.A2(n_9),
.B1(n_10),
.B2(n_5),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_20),
.B1(n_14),
.B2(n_11),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_23),
.Y(n_25)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_19),
.B1(n_20),
.B2(n_15),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_22),
.B2(n_23),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.C(n_27),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_10),
.Y(n_29)
);

A2O1A1O1Ixp25_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_26),
.B(n_10),
.C(n_9),
.D(n_3),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_26),
.Y(n_32)
);


endmodule