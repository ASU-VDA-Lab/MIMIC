module fake_aes_12429_n_693 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_693);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_693;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx10_ASAP7_75t_L g89 ( .A(n_1), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_16), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_79), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_75), .Y(n_92) );
INVx1_ASAP7_75t_SL g93 ( .A(n_71), .Y(n_93) );
BUFx5_ASAP7_75t_L g94 ( .A(n_49), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_86), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_69), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_70), .Y(n_97) );
BUFx2_ASAP7_75t_L g98 ( .A(n_24), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_62), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_65), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_51), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_59), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_88), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_77), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_47), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_33), .B(n_57), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_3), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_34), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_40), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_37), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
BUFx2_ASAP7_75t_SL g112 ( .A(n_7), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_22), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_44), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_55), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_87), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_58), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_50), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_52), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_45), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_41), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_15), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_78), .Y(n_123) );
CKINVDCx14_ASAP7_75t_R g124 ( .A(n_68), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_85), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_53), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_72), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_9), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_73), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_2), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_66), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_84), .Y(n_132) );
INVxp67_ASAP7_75t_SL g133 ( .A(n_54), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_130), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_94), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_118), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_130), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_98), .B(n_0), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_94), .Y(n_139) );
CKINVDCx6p67_ASAP7_75t_R g140 ( .A(n_91), .Y(n_140) );
INVxp33_ASAP7_75t_SL g141 ( .A(n_122), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_92), .B(n_21), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_94), .B(n_1), .Y(n_143) );
NOR2x1_ASAP7_75t_L g144 ( .A(n_95), .B(n_2), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_90), .B(n_3), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_118), .Y(n_148) );
INVx6_ASAP7_75t_L g149 ( .A(n_94), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_122), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_99), .B(n_4), .Y(n_151) );
INVx6_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_124), .B(n_4), .Y(n_153) );
NOR3xp33_ASAP7_75t_L g154 ( .A(n_150), .B(n_111), .C(n_107), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_138), .B(n_128), .Y(n_156) );
INVx1_ASAP7_75t_SL g157 ( .A(n_150), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_147), .B(n_96), .Y(n_158) );
BUFx10_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
INVx4_ASAP7_75t_L g160 ( .A(n_142), .Y(n_160) );
OR2x6_ASAP7_75t_L g161 ( .A(n_153), .B(n_112), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_151), .A2(n_124), .B1(n_89), .B2(n_131), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_141), .B(n_96), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_140), .B(n_115), .Y(n_165) );
NAND3xp33_ASAP7_75t_L g166 ( .A(n_138), .B(n_125), .C(n_132), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
INVx2_ASAP7_75t_SL g168 ( .A(n_149), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_145), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_138), .B(n_125), .Y(n_171) );
NAND2xp33_ASAP7_75t_L g172 ( .A(n_142), .B(n_127), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_151), .A2(n_89), .B1(n_110), .B2(n_129), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_136), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_153), .B(n_89), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_139), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_140), .B(n_100), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_138), .B(n_132), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_165), .B(n_140), .Y(n_184) );
AO22x1_ASAP7_75t_L g185 ( .A1(n_156), .A2(n_142), .B1(n_138), .B2(n_151), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_159), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_180), .Y(n_187) );
NAND2x1_ASAP7_75t_L g188 ( .A(n_180), .B(n_149), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_163), .B(n_147), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_158), .B(n_151), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_181), .B(n_148), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_182), .A2(n_121), .B1(n_136), .B2(n_146), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_180), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_175), .B(n_139), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_175), .B(n_134), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_157), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_180), .B(n_144), .Y(n_198) );
BUFx6f_ASAP7_75t_SL g199 ( .A(n_161), .Y(n_199) );
NOR2x1p5_ASAP7_75t_L g200 ( .A(n_166), .B(n_146), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_154), .A2(n_142), .B1(n_149), .B2(n_152), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_156), .A2(n_142), .B1(n_149), .B2(n_152), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_182), .B(n_134), .Y(n_203) );
OR2x6_ASAP7_75t_L g204 ( .A(n_161), .B(n_144), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_156), .B(n_134), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_155), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_156), .B(n_134), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_155), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_173), .B(n_134), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_171), .B(n_137), .Y(n_210) );
NOR2xp67_ASAP7_75t_L g211 ( .A(n_160), .B(n_137), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_161), .B(n_137), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
OR2x6_ASAP7_75t_L g214 ( .A(n_161), .B(n_143), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_164), .Y(n_215) );
INVx4_ASAP7_75t_L g216 ( .A(n_159), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_183), .B(n_93), .Y(n_217) );
INVx8_ASAP7_75t_L g218 ( .A(n_161), .Y(n_218) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_174), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_160), .A2(n_142), .B1(n_149), .B2(n_152), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_160), .A2(n_142), .B1(n_152), .B2(n_143), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
AND2x6_ASAP7_75t_SL g223 ( .A(n_162), .B(n_106), .Y(n_223) );
NAND2x1_ASAP7_75t_L g224 ( .A(n_187), .B(n_142), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_218), .A2(n_121), .B1(n_160), .B2(n_167), .Y(n_225) );
OR2x2_ASAP7_75t_L g226 ( .A(n_197), .B(n_137), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_216), .B(n_159), .Y(n_227) );
OAI21xp33_ASAP7_75t_L g228 ( .A1(n_197), .A2(n_172), .B(n_169), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_192), .A2(n_169), .B(n_177), .C(n_176), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_185), .A2(n_167), .B(n_178), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_185), .A2(n_167), .B(n_178), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_196), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_216), .B(n_159), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_195), .B(n_167), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_189), .B(n_170), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_190), .A2(n_179), .B(n_178), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_188), .A2(n_179), .B(n_168), .Y(n_237) );
NAND3xp33_ASAP7_75t_L g238 ( .A(n_201), .B(n_202), .C(n_191), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_187), .A2(n_179), .B(n_177), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_218), .A2(n_152), .B1(n_137), .B2(n_170), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_200), .B(n_177), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_216), .B(n_170), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_186), .B(n_176), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_200), .B(n_176), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_186), .B(n_168), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_194), .A2(n_109), .B(n_133), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_188), .A2(n_101), .B(n_102), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_184), .B(n_152), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_218), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_218), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_219), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_212), .B(n_103), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_194), .A2(n_116), .B(n_126), .Y(n_253) );
NOR3xp33_ASAP7_75t_L g254 ( .A(n_217), .B(n_113), .C(n_123), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_212), .B(n_142), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_204), .B(n_104), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_220), .B(n_105), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_209), .A2(n_205), .B(n_207), .Y(n_258) );
AOI21xp5_ASAP7_75t_SL g259 ( .A1(n_225), .A2(n_199), .B(n_214), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_230), .A2(n_211), .B(n_210), .Y(n_260) );
AO32x2_ASAP7_75t_L g261 ( .A1(n_240), .A2(n_223), .A3(n_198), .B1(n_204), .B2(n_214), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_232), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_239), .A2(n_193), .B(n_222), .Y(n_263) );
CKINVDCx11_ASAP7_75t_R g264 ( .A(n_249), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_231), .A2(n_211), .B(n_203), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_234), .A2(n_214), .B(n_222), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_SL g267 ( .A1(n_224), .A2(n_108), .B(n_120), .C(n_117), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_258), .A2(n_214), .B(n_193), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_241), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_249), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_229), .A2(n_204), .B(n_119), .C(n_215), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_256), .B(n_204), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_256), .B(n_198), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_226), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_SL g275 ( .A1(n_258), .A2(n_106), .B(n_206), .C(n_215), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_236), .A2(n_206), .B(n_213), .Y(n_276) );
BUFx12f_ASAP7_75t_L g277 ( .A(n_249), .Y(n_277) );
AO32x2_ASAP7_75t_L g278 ( .A1(n_228), .A2(n_223), .A3(n_198), .B1(n_199), .B2(n_221), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_251), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_254), .B(n_198), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_238), .A2(n_199), .B1(n_208), .B2(n_213), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_250), .B(n_198), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_237), .A2(n_208), .B(n_198), .Y(n_283) );
NOR2xp67_ASAP7_75t_L g284 ( .A(n_246), .B(n_5), .Y(n_284) );
NOR2x1_ASAP7_75t_L g285 ( .A(n_259), .B(n_244), .Y(n_285) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_283), .A2(n_247), .B(n_253), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_275), .A2(n_255), .B(n_257), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_262), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_262), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_269), .B(n_242), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_263), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_277), .Y(n_292) );
AO31x2_ASAP7_75t_L g293 ( .A1(n_268), .A2(n_246), .A3(n_235), .B(n_198), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_277), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_261), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_266), .A2(n_252), .B(n_248), .Y(n_296) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_265), .A2(n_243), .B(n_245), .Y(n_297) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_276), .A2(n_233), .B(n_227), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_269), .B(n_114), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_280), .B(n_5), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_271), .A2(n_6), .B(n_7), .Y(n_301) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_260), .A2(n_114), .B(n_48), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_278), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_275), .A2(n_114), .B(n_8), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_274), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_273), .B(n_114), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_288), .Y(n_308) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_303), .A2(n_281), .B(n_282), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_299), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_288), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_289), .B(n_272), .Y(n_312) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_304), .A2(n_267), .B(n_278), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_289), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_299), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_299), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_306), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_293), .B(n_270), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_299), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_291), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_305), .B(n_279), .Y(n_321) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_299), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_294), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_306), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_295), .B(n_261), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_293), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_290), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_293), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_293), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_293), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_293), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_295), .B(n_261), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_293), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_295), .B(n_261), .Y(n_335) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_303), .A2(n_291), .B(n_287), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_319), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_327), .B(n_303), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_325), .B(n_304), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_308), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_308), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_325), .B(n_304), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_327), .B(n_291), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_326), .B(n_300), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_325), .B(n_304), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_326), .B(n_300), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_333), .B(n_304), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_333), .B(n_290), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_319), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_333), .B(n_290), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_311), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_321), .B(n_294), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_328), .B(n_294), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_310), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_335), .B(n_290), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_314), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_335), .B(n_290), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_328), .B(n_305), .Y(n_364) );
INVx2_ASAP7_75t_SL g365 ( .A(n_310), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_327), .B(n_285), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_310), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_329), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_327), .B(n_285), .Y(n_369) );
NAND2x1_ASAP7_75t_L g370 ( .A(n_316), .B(n_302), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_329), .B(n_301), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_336), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_331), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_336), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_331), .B(n_301), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_335), .B(n_278), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_332), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_332), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_336), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_334), .B(n_298), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_334), .B(n_278), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_322), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_336), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_330), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_372), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_364), .B(n_317), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_340), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_364), .B(n_317), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_341), .B(n_324), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_344), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_366), .B(n_330), .Y(n_391) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_337), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_342), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_384), .B(n_318), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_384), .B(n_318), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_372), .Y(n_397) );
AND2x2_ASAP7_75t_SL g398 ( .A(n_351), .B(n_302), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_354), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_372), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_350), .B(n_324), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_354), .B(n_312), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_374), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_355), .B(n_361), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_350), .B(n_322), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_357), .B(n_353), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_366), .B(n_315), .Y(n_408) );
NAND2x1p5_ASAP7_75t_SL g409 ( .A(n_358), .B(n_316), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_361), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_357), .B(n_312), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_353), .B(n_336), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_366), .B(n_315), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_337), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_368), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_368), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_360), .B(n_336), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_356), .A2(n_315), .B1(n_316), .B2(n_312), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_360), .B(n_315), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_373), .B(n_323), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_363), .B(n_309), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_377), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_363), .B(n_309), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_376), .B(n_309), .Y(n_428) );
NAND2x1_ASAP7_75t_L g429 ( .A(n_367), .B(n_302), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_374), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_379), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_378), .B(n_292), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_376), .B(n_309), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_339), .B(n_309), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_352), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_339), .B(n_313), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_382), .B(n_313), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_343), .B(n_313), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_352), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_379), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_343), .B(n_292), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_352), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_347), .B(n_313), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_359), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_359), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_379), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_359), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_362), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_344), .B(n_264), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_383), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_344), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_347), .B(n_313), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_393), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_412), .B(n_349), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_441), .B(n_346), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_412), .B(n_381), .Y(n_456) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_449), .B(n_370), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_417), .B(n_381), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_417), .B(n_380), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_398), .A2(n_370), .B(n_371), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_395), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_402), .B(n_380), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_422), .B(n_380), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_422), .B(n_380), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_427), .B(n_338), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_431), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_427), .B(n_338), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_428), .B(n_338), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_428), .B(n_338), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_433), .B(n_383), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_433), .B(n_383), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_434), .B(n_345), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_426), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_407), .B(n_346), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_414), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_407), .B(n_348), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_434), .B(n_345), .Y(n_477) );
AND2x4_ASAP7_75t_SL g478 ( .A(n_408), .B(n_367), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_402), .B(n_348), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_410), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_414), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_436), .B(n_345), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_421), .B(n_6), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_391), .B(n_367), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_386), .B(n_375), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_394), .B(n_375), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_436), .B(n_345), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_438), .B(n_367), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_388), .B(n_371), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_394), .B(n_396), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_431), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_401), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_438), .B(n_362), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_443), .B(n_362), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_432), .B(n_358), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_387), .B(n_358), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_443), .B(n_365), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_452), .B(n_365), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_396), .B(n_365), .Y(n_499) );
INVx2_ASAP7_75t_SL g500 ( .A(n_390), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_452), .B(n_366), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_431), .B(n_369), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_399), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_385), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_411), .B(n_369), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_406), .B(n_302), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_406), .B(n_302), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_391), .B(n_297), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_425), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_405), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_401), .B(n_8), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_392), .B(n_9), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_391), .B(n_297), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_420), .B(n_297), .Y(n_514) );
AND2x2_ASAP7_75t_SL g515 ( .A(n_398), .B(n_286), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_420), .B(n_297), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_385), .B(n_297), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_397), .B(n_286), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_397), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_451), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_400), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_451), .B(n_307), .Y(n_522) );
INVx3_ASAP7_75t_L g523 ( .A(n_400), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_403), .B(n_10), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_437), .B(n_10), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_415), .B(n_11), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_408), .B(n_298), .Y(n_527) );
NOR2x1p5_ASAP7_75t_L g528 ( .A(n_429), .B(n_11), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_404), .B(n_286), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_404), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_490), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_510), .B(n_416), .Y(n_532) );
NAND2x1_ASAP7_75t_L g533 ( .A(n_457), .B(n_424), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_456), .B(n_408), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_474), .B(n_424), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_473), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_524), .A2(n_418), .B1(n_413), .B2(n_389), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_483), .B(n_413), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_454), .B(n_419), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_523), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_500), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_456), .B(n_413), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_528), .A2(n_423), .B1(n_450), .B2(n_430), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_458), .B(n_430), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_458), .B(n_454), .Y(n_545) );
NOR2x1_ASAP7_75t_L g546 ( .A(n_511), .B(n_429), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_503), .Y(n_547) );
OAI21xp33_ASAP7_75t_L g548 ( .A1(n_511), .A2(n_437), .B(n_440), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_523), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_500), .B(n_440), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_501), .B(n_446), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_474), .B(n_450), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_501), .B(n_435), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_515), .A2(n_448), .B1(n_447), .B2(n_445), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_459), .B(n_435), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_459), .B(n_439), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_476), .B(n_409), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_486), .B(n_442), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_520), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_472), .B(n_445), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_472), .B(n_447), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_475), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_470), .B(n_409), .Y(n_563) );
AND2x2_ASAP7_75t_SL g564 ( .A(n_478), .B(n_448), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_453), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_523), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_477), .B(n_444), .Y(n_567) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_484), .B(n_307), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_478), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_477), .B(n_307), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_463), .B(n_307), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_461), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_485), .B(n_12), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_479), .B(n_13), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_489), .B(n_13), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_470), .B(n_14), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_481), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_499), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_493), .B(n_14), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_484), .B(n_15), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_493), .B(n_16), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_455), .B(n_525), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_494), .B(n_17), .Y(n_583) );
OAI21xp33_ASAP7_75t_L g584 ( .A1(n_525), .A2(n_296), .B(n_287), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_463), .B(n_286), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_530), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_471), .B(n_17), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_494), .B(n_18), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_515), .A2(n_296), .B1(n_286), .B2(n_267), .Y(n_589) );
CKINVDCx16_ASAP7_75t_R g590 ( .A(n_484), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_471), .B(n_18), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_455), .B(n_19), .Y(n_592) );
OR2x6_ASAP7_75t_L g593 ( .A(n_522), .B(n_19), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_464), .B(n_497), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_530), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_531), .B(n_464), .Y(n_597) );
AOI21xp33_ASAP7_75t_SL g598 ( .A1(n_564), .A2(n_512), .B(n_492), .Y(n_598) );
OAI32xp33_ASAP7_75t_L g599 ( .A1(n_590), .A2(n_557), .A3(n_559), .B1(n_577), .B2(n_563), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_593), .A2(n_460), .B(n_495), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_537), .A2(n_512), .B1(n_462), .B2(n_505), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_535), .B(n_488), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_552), .B(n_488), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_546), .B(n_543), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_593), .A2(n_496), .B(n_526), .Y(n_605) );
AOI21xp33_ASAP7_75t_SL g606 ( .A1(n_569), .A2(n_506), .B(n_507), .Y(n_606) );
NAND4xp25_ASAP7_75t_L g607 ( .A(n_537), .B(n_527), .C(n_506), .D(n_507), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_SL g608 ( .A1(n_541), .A2(n_509), .B(n_480), .C(n_466), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_592), .A2(n_527), .B(n_491), .C(n_466), .Y(n_609) );
OR4x1_ASAP7_75t_L g610 ( .A(n_536), .B(n_527), .C(n_498), .D(n_502), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_545), .B(n_482), .Y(n_611) );
INVxp67_ASAP7_75t_L g612 ( .A(n_562), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_558), .Y(n_613) );
AOI211x1_ASAP7_75t_L g614 ( .A1(n_548), .A2(n_465), .B(n_467), .C(n_468), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_593), .A2(n_487), .B1(n_482), .B2(n_465), .Y(n_615) );
NAND3xp33_ASAP7_75t_SL g616 ( .A(n_559), .B(n_513), .C(n_508), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_532), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_550), .A2(n_502), .B(n_514), .Y(n_618) );
AOI221xp5_ASAP7_75t_SL g619 ( .A1(n_582), .A2(n_487), .B1(n_468), .B2(n_469), .C(n_467), .Y(n_619) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_575), .A2(n_529), .B(n_518), .Y(n_620) );
AND2x4_ASAP7_75t_L g621 ( .A(n_534), .B(n_469), .Y(n_621) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_580), .B(n_504), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_577), .B(n_516), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_576), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_548), .A2(n_508), .B1(n_521), .B2(n_519), .C(n_504), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_554), .B(n_521), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_547), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_533), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_573), .B(n_519), .C(n_529), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_581), .A2(n_517), .B(n_20), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_539), .B(n_517), .Y(n_631) );
NAND3xp33_ASAP7_75t_SL g632 ( .A(n_587), .B(n_20), .C(n_23), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_542), .B(n_25), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_594), .B(n_26), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_539), .B(n_27), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_544), .B(n_28), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_555), .B(n_29), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_578), .Y(n_638) );
AOI31xp33_ASAP7_75t_L g639 ( .A1(n_619), .A2(n_538), .A3(n_591), .B(n_583), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_614), .A2(n_574), .B1(n_581), .B2(n_583), .C(n_579), .Y(n_640) );
NAND4xp75_ASAP7_75t_L g641 ( .A(n_619), .B(n_588), .C(n_554), .D(n_585), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_598), .A2(n_568), .B(n_556), .C(n_560), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_599), .A2(n_595), .B1(n_571), .B2(n_570), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_632), .B(n_584), .C(n_595), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_617), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_618), .A2(n_561), .B(n_567), .C(n_553), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_624), .B(n_572), .Y(n_647) );
AOI31xp33_ASAP7_75t_L g648 ( .A1(n_604), .A2(n_584), .A3(n_551), .B(n_589), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_600), .A2(n_589), .B1(n_565), .B2(n_586), .C(n_566), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_616), .A2(n_596), .B(n_549), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_607), .A2(n_540), .B1(n_30), .B2(n_31), .C(n_32), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_601), .A2(n_35), .B1(n_36), .B2(n_38), .C(n_39), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_615), .A2(n_42), .B1(n_43), .B2(n_46), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_606), .A2(n_630), .B(n_609), .C(n_629), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_638), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_610), .A2(n_56), .B1(n_60), .B2(n_61), .C(n_63), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_627), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_608), .A2(n_64), .B(n_67), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_626), .A2(n_74), .B(n_76), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_613), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_625), .A2(n_80), .B1(n_81), .B2(n_82), .C(n_83), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_605), .A2(n_620), .B(n_634), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_628), .A2(n_623), .B1(n_635), .B2(n_597), .C(n_631), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_628), .A2(n_611), .B1(n_621), .B2(n_602), .C(n_603), .Y(n_664) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_633), .B(n_630), .C(n_614), .D(n_537), .Y(n_665) );
OAI322xp33_ASAP7_75t_L g666 ( .A1(n_637), .A2(n_612), .A3(n_601), .B1(n_604), .B2(n_615), .C1(n_624), .C2(n_582), .Y(n_666) );
NOR4xp25_ASAP7_75t_L g667 ( .A(n_636), .B(n_604), .C(n_612), .D(n_624), .Y(n_667) );
NAND3x1_ASAP7_75t_L g668 ( .A(n_622), .B(n_600), .C(n_628), .Y(n_668) );
NAND3xp33_ASAP7_75t_SL g669 ( .A(n_667), .B(n_654), .C(n_656), .Y(n_669) );
NOR2x2_ASAP7_75t_L g670 ( .A(n_641), .B(n_668), .Y(n_670) );
NAND4xp25_ASAP7_75t_SL g671 ( .A(n_643), .B(n_642), .C(n_664), .D(n_640), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_655), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_657), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_662), .B(n_646), .Y(n_674) );
AOI211xp5_ASAP7_75t_L g675 ( .A1(n_666), .A2(n_651), .B(n_665), .C(n_644), .Y(n_675) );
NAND4xp25_ASAP7_75t_SL g676 ( .A(n_658), .B(n_649), .C(n_639), .D(n_653), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_672), .B(n_648), .Y(n_677) );
NOR3xp33_ASAP7_75t_L g678 ( .A(n_669), .B(n_652), .C(n_661), .Y(n_678) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_673), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_675), .B(n_647), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_677), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_680), .B(n_676), .Y(n_682) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_679), .B(n_676), .Y(n_683) );
OAI21x1_ASAP7_75t_SL g684 ( .A1(n_682), .A2(n_670), .B(n_650), .Y(n_684) );
CKINVDCx16_ASAP7_75t_R g685 ( .A(n_681), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_685), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_684), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_686), .B(n_671), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_687), .A2(n_683), .B1(n_674), .B2(n_678), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_689), .B(n_660), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_690), .B(n_688), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_691), .B(n_645), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_692), .A2(n_663), .B(n_659), .Y(n_693) );
endmodule