module real_jpeg_28948_n_17 (n_5, n_4, n_8, n_0, n_12, n_318, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_318;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_0),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_28),
.B1(n_63),
.B2(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_0),
.A2(n_28),
.B1(n_48),
.B2(n_50),
.Y(n_242)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_53),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_3),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_3),
.A2(n_48),
.B1(n_50),
.B2(n_135),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_135),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_135),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_5),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_69),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_69),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_6),
.A2(n_40),
.B1(n_48),
.B2(n_50),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_66),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_8),
.A2(n_48),
.B1(n_50),
.B2(n_66),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_66),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_10),
.B(n_35),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_10),
.A2(n_35),
.B(n_43),
.C(n_149),
.D(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_10),
.B(n_32),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_10),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_10),
.A2(n_82),
.B(n_166),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_10),
.A2(n_30),
.B(n_31),
.C(n_199),
.D(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_10),
.B(n_30),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_10),
.B(n_59),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_10),
.A2(n_61),
.B(n_64),
.C(n_244),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_181),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_11),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_97),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_97),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_97),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_12),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_12),
.A2(n_48),
.B1(n_50),
.B2(n_161),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_161),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_161),
.Y(n_272)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_13),
.A2(n_35),
.B(n_44),
.C(n_47),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_13),
.B(n_48),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_113),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_98),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_21),
.B(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.C(n_79),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_22),
.A2(n_23),
.B1(n_71),
.B2(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_56),
.B2(n_70),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_26),
.B(n_55),
.C(n_56),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_29),
.A2(n_30),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g209 ( 
.A1(n_29),
.A2(n_35),
.A3(n_199),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_30),
.A2(n_60),
.B(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_31),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_31),
.A2(n_32),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_33),
.Y(n_211)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_34),
.A2(n_46),
.A3(n_50),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_34),
.B(n_211),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_39),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_41),
.A2(n_55),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_51),
.B(n_52),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_42),
.A2(n_51),
.B1(n_92),
.B2(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_42),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_42),
.A2(n_51),
.B1(n_129),
.B2(n_258),
.Y(n_277)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_47),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_43),
.A2(n_47),
.B1(n_74),
.B2(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_43),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_43),
.A2(n_47),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_83),
.Y(n_82)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_50),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_51),
.B(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_51),
.A2(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_51),
.B(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_51),
.A2(n_162),
.B(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_70),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_57),
.A2(n_67),
.B1(n_68),
.B2(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_57),
.A2(n_133),
.B(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_58),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_58),
.A2(n_59),
.B1(n_134),
.B2(n_272),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_59),
.B(n_96),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_67),
.B(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_67),
.A2(n_95),
.B(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_73),
.B(n_76),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_107),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_79),
.A2(n_80),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_88),
.B(n_93),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_93),
.B1(n_94),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_81),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_81),
.A2(n_89),
.B1(n_90),
.B2(n_119),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_87),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_87),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_82),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_82),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_82),
.B(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_82),
.A2(n_86),
.B1(n_208),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_82),
.A2(n_86),
.B1(n_126),
.B2(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_84),
.A2(n_173),
.B(n_183),
.Y(n_182)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_SL g127 ( 
.A(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_85),
.B(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_85),
.A2(n_184),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_85),
.A2(n_174),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_111),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_107),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_109),
.B(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_109),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_109),
.A2(n_131),
.B(n_220),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_140),
.B(n_316),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_137),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_115),
.B(n_137),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_304)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_122),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.C(n_132),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_123),
.A2(n_124),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_125),
.B(n_128),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_130),
.B(n_132),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_136),
.Y(n_250)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI321xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_296),
.A3(n_305),
.B1(n_310),
.B2(n_315),
.C(n_318),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_260),
.C(n_292),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_234),
.B(n_259),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_214),
.B(n_233),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_194),
.B(n_213),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_169),
.B(n_193),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_147),
.B(n_154),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_151),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_152),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_159),
.C(n_164),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_178),
.B(n_192),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_177),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_185),
.B(n_191),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_180),
.B(n_182),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_195),
.B(n_196),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_205),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_202),
.C(n_205),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_200),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_204),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_209),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_215),
.B(n_216),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_228),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_229),
.C(n_230),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_223),
.C(n_226),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_219),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_227),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_236),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_247),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_238),
.B(n_239),
.C(n_247),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_242),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_245),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_253),
.C(n_256),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_257),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_255),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_261),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_279),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_262),
.B(n_279),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_274),
.C(n_278),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_266),
.C(n_273),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_270),
.B2(n_273),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_270),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_278),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_277),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_288),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_288),
.C(n_291),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_285),
.C(n_286),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_294),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_303),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_303),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.C(n_302),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_301),
.Y(n_309)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_311),
.B(n_314),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_307),
.B(n_308),
.Y(n_314)
);


endmodule