module fake_ibex_576_n_3763 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_768, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_592, n_495, n_762, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_3763);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_768;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_3763;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_3750;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_3458;
wire n_2955;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_3211;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3395;
wire n_3242;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_2436;
wire n_1663;
wire n_2333;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3097;
wire n_2906;
wire n_3030;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3667;
wire n_3221;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_2373;
wire n_1927;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3023;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_1969;
wire n_1296;
wire n_3060;
wire n_1326;
wire n_971;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_3217;
wire n_1787;
wire n_2782;
wire n_2401;
wire n_2511;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_3471;
wire n_3320;
wire n_3117;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_3524;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_2176;
wire n_1884;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_3357;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_2252;
wire n_1982;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_2294;
wire n_1977;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_3236;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_998;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_3587;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3401;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_3070;
wire n_2842;
wire n_2711;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_991;
wire n_1331;
wire n_1223;
wire n_961;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_3585;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_3512;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_3538;
wire n_2299;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2675;
wire n_2576;
wire n_2417;
wire n_2348;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_3066;
wire n_2714;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_3102;
wire n_2872;
wire n_3173;
wire n_2790;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3305;
wire n_1635;
wire n_1572;
wire n_3051;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3742;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_3430;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_2689;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_849;
wire n_1193;
wire n_2928;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3380;
wire n_1074;
wire n_3557;
wire n_3067;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3622;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2302;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3550;
wire n_3261;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_364),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_286),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_111),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_176),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_508),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_737),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_96),
.Y(n_800)
);

CKINVDCx16_ASAP7_75t_R g801 ( 
.A(n_553),
.Y(n_801)
);

BUFx5_ASAP7_75t_L g802 ( 
.A(n_133),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_9),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_774),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_142),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_670),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_757),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_411),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_460),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_549),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_657),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_272),
.Y(n_812)
);

BUFx2_ASAP7_75t_SL g813 ( 
.A(n_307),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_241),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_583),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_359),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_554),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_36),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_410),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_687),
.B(n_363),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_359),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_581),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_557),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_39),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_660),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_757),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_660),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_191),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_687),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_725),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_630),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_388),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_70),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_373),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_608),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_79),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_66),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_469),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_678),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_762),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_403),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_80),
.Y(n_842)
);

CKINVDCx14_ASAP7_75t_R g843 ( 
.A(n_25),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_179),
.B(n_166),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_473),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_691),
.Y(n_846)
);

BUFx5_ASAP7_75t_L g847 ( 
.A(n_232),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_742),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_390),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_397),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_589),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_334),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_679),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_290),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_353),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_316),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_217),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_61),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_200),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_588),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_425),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_232),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_134),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_347),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_349),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_83),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_419),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_337),
.Y(n_868)
);

BUFx10_ASAP7_75t_L g869 ( 
.A(n_345),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_707),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_451),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_545),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_407),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_706),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_77),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_187),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_680),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_542),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_624),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_559),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_740),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_364),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_396),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_632),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_728),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_120),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_587),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_655),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_303),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_57),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_63),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_739),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_210),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_589),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_314),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_127),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_636),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_418),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_637),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_167),
.Y(n_900)
);

BUFx2_ASAP7_75t_SL g901 ( 
.A(n_534),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_501),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_714),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_507),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_551),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_142),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_111),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_385),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_62),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_536),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_517),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_469),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_580),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_635),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_312),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_598),
.Y(n_916)
);

CKINVDCx16_ASAP7_75t_R g917 ( 
.A(n_628),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_484),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_670),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_172),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_583),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_681),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_258),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_477),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_680),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_450),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_758),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_29),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_245),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_570),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_L g931 ( 
.A(n_524),
.B(n_522),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_153),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_68),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_134),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_705),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_790),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_629),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_30),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_249),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_258),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_12),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_633),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_336),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_293),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_132),
.Y(n_945)
);

BUFx8_ASAP7_75t_SL g946 ( 
.A(n_283),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_60),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_603),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_236),
.Y(n_949)
);

BUFx2_ASAP7_75t_SL g950 ( 
.A(n_74),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_714),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_786),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_120),
.B(n_65),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_265),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_6),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_91),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_450),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_598),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_783),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_742),
.B(n_83),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_326),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_275),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_18),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_117),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_260),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_72),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_651),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_82),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_148),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_567),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_444),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_780),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_114),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_380),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_315),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_242),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_673),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_329),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_724),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_474),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_572),
.Y(n_981)
);

CKINVDCx16_ASAP7_75t_R g982 ( 
.A(n_705),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_198),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_160),
.B(n_681),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_97),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_707),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_630),
.Y(n_987)
);

NOR2xp67_ASAP7_75t_L g988 ( 
.A(n_245),
.B(n_382),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_754),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_762),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_419),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_21),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_711),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_734),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_787),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_625),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_266),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_26),
.Y(n_998)
);

CKINVDCx16_ASAP7_75t_R g999 ( 
.A(n_221),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_152),
.Y(n_1000)
);

CKINVDCx14_ASAP7_75t_R g1001 ( 
.A(n_606),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_392),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_81),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_628),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_485),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_225),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_684),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_518),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_656),
.Y(n_1009)
);

INVxp33_ASAP7_75t_L g1010 ( 
.A(n_597),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_252),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_421),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_743),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_585),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_698),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_793),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_764),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_193),
.Y(n_1018)
);

CKINVDCx16_ASAP7_75t_R g1019 ( 
.A(n_22),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_785),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_235),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_139),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_141),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_90),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_709),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_435),
.Y(n_1026)
);

BUFx10_ASAP7_75t_L g1027 ( 
.A(n_502),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_644),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_284),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_505),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_548),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_9),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_285),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_222),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_483),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_31),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_265),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_353),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_720),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_702),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_170),
.Y(n_1041)
);

CKINVDCx16_ASAP7_75t_R g1042 ( 
.A(n_389),
.Y(n_1042)
);

CKINVDCx16_ASAP7_75t_R g1043 ( 
.A(n_343),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_234),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_164),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_77),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_732),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_616),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_584),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_127),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_588),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_414),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_468),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_236),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_750),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_487),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_725),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_392),
.B(n_612),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_778),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_324),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_325),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_357),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_367),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_604),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_275),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_577),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_298),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_76),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_382),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_381),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_198),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_235),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_164),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_268),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_166),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_603),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_728),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_108),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_547),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_643),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_259),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_148),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_299),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_791),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_640),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_354),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_402),
.Y(n_1087)
);

BUFx10_ASAP7_75t_L g1088 ( 
.A(n_349),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_692),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_33),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_281),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_194),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_789),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_34),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_605),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_25),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_618),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_101),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_51),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_172),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_226),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_304),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_323),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_49),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_609),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_665),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_644),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_29),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_729),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_492),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_640),
.Y(n_1111)
);

BUFx5_ASAP7_75t_L g1112 ( 
.A(n_205),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_222),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_461),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_613),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_480),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_412),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_467),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_68),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_467),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_242),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_343),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_586),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_620),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_596),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_633),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_98),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_407),
.Y(n_1128)
);

BUFx2_ASAP7_75t_SL g1129 ( 
.A(n_623),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_318),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_116),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_465),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_462),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_197),
.Y(n_1134)
);

CKINVDCx14_ASAP7_75t_R g1135 ( 
.A(n_145),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_496),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_658),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_228),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_523),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_321),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_720),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_521),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_770),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_446),
.Y(n_1144)
);

BUFx10_ASAP7_75t_L g1145 ( 
.A(n_437),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_183),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_776),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_335),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_215),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_472),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_746),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_226),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_112),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_400),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_529),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_426),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_188),
.Y(n_1157)
);

INVxp33_ASAP7_75t_L g1158 ( 
.A(n_463),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_684),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_721),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_200),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_145),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_135),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_619),
.B(n_413),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_360),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_735),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_750),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_180),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_648),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_317),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_495),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_459),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_530),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_319),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_411),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_L g1176 ( 
.A(n_110),
.B(n_590),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_23),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_370),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_624),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_453),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_6),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_217),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_386),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_632),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_280),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_645),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_214),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_128),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_510),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_400),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_90),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_189),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_362),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_673),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_711),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_432),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_795),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_829),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_843),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_843),
.Y(n_1200)
);

CKINVDCx6p67_ASAP7_75t_R g1201 ( 
.A(n_869),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1001),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_802),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1001),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_839),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_802),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_952),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_795),
.Y(n_1208)
);

INVxp33_ASAP7_75t_SL g1209 ( 
.A(n_797),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_802),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_795),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_802),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_802),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_869),
.Y(n_1214)
);

INVx5_ASAP7_75t_L g1215 ( 
.A(n_952),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_802),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_795),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1135),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_839),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_869),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1010),
.B(n_3),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_806),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_856),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_802),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1027),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1020),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_806),
.Y(n_1227)
);

BUFx8_ASAP7_75t_L g1228 ( 
.A(n_942),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1016),
.A2(n_782),
.B(n_781),
.Y(n_1229)
);

BUFx8_ASAP7_75t_SL g1230 ( 
.A(n_946),
.Y(n_1230)
);

BUFx8_ASAP7_75t_L g1231 ( 
.A(n_969),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_870),
.B(n_926),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_870),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_875),
.B(n_4),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_927),
.B(n_4),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1027),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_926),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_936),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1016),
.A2(n_995),
.B(n_959),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1027),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_965),
.B(n_5),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_847),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_806),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1135),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_965),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1010),
.Y(n_1246)
);

AND2x6_ASAP7_75t_L g1247 ( 
.A(n_1093),
.B(n_784),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1088),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_980),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_847),
.Y(n_1250)
);

INVx5_ASAP7_75t_L g1251 ( 
.A(n_806),
.Y(n_1251)
);

BUFx8_ASAP7_75t_SL g1252 ( 
.A(n_946),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_847),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1158),
.B(n_5),
.Y(n_1254)
);

CKINVDCx6p67_ASAP7_75t_R g1255 ( 
.A(n_1088),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_847),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_975),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1088),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1158),
.B(n_7),
.Y(n_1259)
);

OAI22x1_ASAP7_75t_L g1260 ( 
.A1(n_892),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_SL g1261 ( 
.A(n_1084),
.B(n_788),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_799),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1078),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_871),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1078),
.B(n_10),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_871),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1120),
.B(n_11),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1120),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1146),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_847),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_871),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_878),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_847),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_878),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_957),
.B(n_981),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1146),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_985),
.B(n_12),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_929),
.Y(n_1278)
);

CKINVDCx16_ASAP7_75t_R g1279 ( 
.A(n_801),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1174),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1112),
.Y(n_1281)
);

BUFx8_ASAP7_75t_L g1282 ( 
.A(n_1127),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1145),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_917),
.Y(n_1284)
);

OAI22x1_ASAP7_75t_R g1285 ( 
.A1(n_794),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1174),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1186),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1145),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1186),
.B(n_14),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_933),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_878),
.Y(n_1291)
);

INVx4_ASAP7_75t_L g1292 ( 
.A(n_878),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1153),
.Y(n_1293)
);

BUFx8_ASAP7_75t_L g1294 ( 
.A(n_1112),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_804),
.B(n_15),
.Y(n_1295)
);

INVx5_ASAP7_75t_L g1296 ( 
.A(n_883),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1203),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1206),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1294),
.B(n_1112),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1295),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1280),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1294),
.B(n_1112),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1295),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1280),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1232),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1246),
.B(n_982),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1238),
.B(n_1009),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1214),
.B(n_1026),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1210),
.B(n_1112),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1232),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1212),
.B(n_1213),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1246),
.B(n_999),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1207),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1216),
.B(n_1112),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1224),
.B(n_1112),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1207),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1200),
.B(n_1244),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1242),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1250),
.B(n_883),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1253),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1256),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1270),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1201),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1241),
.Y(n_1324)
);

AND3x2_ASAP7_75t_L g1325 ( 
.A(n_1257),
.B(n_1178),
.C(n_1105),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1265),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1273),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1281),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1239),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1239),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1197),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1265),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1220),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1267),
.B(n_883),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1267),
.B(n_883),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1197),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1197),
.Y(n_1337)
);

NAND2xp33_ASAP7_75t_L g1338 ( 
.A(n_1247),
.B(n_902),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1208),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1209),
.A2(n_1019),
.B1(n_1042),
.B2(n_1040),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1208),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1289),
.Y(n_1342)
);

CKINVDCx6p67_ASAP7_75t_R g1343 ( 
.A(n_1255),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1208),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1211),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1211),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1217),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1217),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1217),
.Y(n_1349)
);

INVx6_ASAP7_75t_L g1350 ( 
.A(n_1240),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1229),
.A2(n_820),
.B(n_809),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1225),
.B(n_1043),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1198),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1205),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1222),
.Y(n_1355)
);

AND3x2_ASAP7_75t_L g1356 ( 
.A(n_1262),
.B(n_984),
.C(n_838),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1215),
.B(n_902),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1222),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1227),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1284),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1226),
.Y(n_1361)
);

NAND2xp33_ASAP7_75t_L g1362 ( 
.A(n_1247),
.B(n_925),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1219),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1230),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1236),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1202),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1262),
.B(n_836),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1209),
.A2(n_798),
.B1(n_803),
.B2(n_800),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1283),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1234),
.A2(n_810),
.B(n_807),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1292),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1223),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1292),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1283),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1233),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1251),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1237),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1215),
.B(n_925),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1251),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1278),
.B(n_1153),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1296),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1234),
.A2(n_814),
.B(n_812),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1245),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1249),
.Y(n_1384)
);

CKINVDCx6p67_ASAP7_75t_R g1385 ( 
.A(n_1279),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1293),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1290),
.B(n_1202),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1278),
.B(n_1153),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1263),
.B(n_1268),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1290),
.A2(n_805),
.B1(n_815),
.B2(n_808),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1276),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1286),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1284),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1287),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1227),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1247),
.Y(n_1396)
);

NAND2xp33_ASAP7_75t_L g1397 ( 
.A(n_1218),
.B(n_930),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1235),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1235),
.Y(n_1399)
);

NAND3x1_ASAP7_75t_L g1400 ( 
.A(n_1204),
.B(n_984),
.C(n_811),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1248),
.B(n_930),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1227),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1243),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1243),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1218),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1277),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1258),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1243),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1275),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1275),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1288),
.B(n_816),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1254),
.B(n_817),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1264),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1264),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1261),
.B(n_1259),
.Y(n_1415)
);

NOR2x1p5_ASAP7_75t_L g1416 ( 
.A(n_1230),
.B(n_834),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1221),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_SL g1418 ( 
.A(n_1252),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1264),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1266),
.Y(n_1420)
);

CKINVDCx6p67_ASAP7_75t_R g1421 ( 
.A(n_1260),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1266),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1271),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1271),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1271),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1272),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1274),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1274),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1274),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1291),
.B(n_930),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1204),
.B(n_804),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1228),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1291),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1252),
.Y(n_1434)
);

AND3x2_ASAP7_75t_L g1435 ( 
.A(n_1285),
.B(n_1282),
.C(n_1231),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1199),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1199),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1228),
.B(n_838),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1231),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1282),
.B(n_958),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_L g1441 ( 
.A(n_1247),
.B(n_958),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1295),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1295),
.Y(n_1443)
);

INVxp33_ASAP7_75t_L g1444 ( 
.A(n_1246),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1203),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1294),
.B(n_958),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1295),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1269),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1269),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_1246),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1409),
.B(n_818),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1410),
.B(n_1398),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1312),
.B(n_1367),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1305),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1399),
.B(n_821),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1450),
.Y(n_1456)
);

NOR2xp67_ASAP7_75t_L g1457 ( 
.A(n_1406),
.B(n_792),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1417),
.B(n_1444),
.Y(n_1458)
);

NOR2xp67_ASAP7_75t_L g1459 ( 
.A(n_1299),
.B(n_1302),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1450),
.B(n_824),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1306),
.B(n_890),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1431),
.A2(n_1195),
.B1(n_825),
.B2(n_827),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1350),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1310),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1380),
.B(n_826),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1388),
.B(n_828),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1412),
.B(n_831),
.Y(n_1467)
);

INVxp67_ASAP7_75t_SL g1468 ( 
.A(n_1329),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1437),
.A2(n_1164),
.B1(n_953),
.B2(n_835),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1323),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1432),
.B(n_813),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1391),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_SL g1473 ( 
.A(n_1439),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1390),
.B(n_852),
.C(n_851),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1365),
.B(n_854),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1342),
.B(n_855),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1352),
.A2(n_1184),
.B1(n_1187),
.B2(n_1182),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1350),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1396),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1342),
.B(n_857),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1330),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1391),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1365),
.B(n_860),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1301),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1369),
.B(n_1374),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1369),
.B(n_863),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1304),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1392),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1392),
.Y(n_1489)
);

INVxp33_ASAP7_75t_L g1490 ( 
.A(n_1352),
.Y(n_1490)
);

A2O1A1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1303),
.A2(n_822),
.B(n_823),
.C(n_819),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1374),
.B(n_865),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1330),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1350),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1300),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1387),
.B(n_1333),
.Y(n_1496)
);

AO221x1_ASAP7_75t_L g1497 ( 
.A1(n_1340),
.A2(n_811),
.B1(n_833),
.B2(n_830),
.C(n_794),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1407),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1386),
.B(n_866),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1407),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1324),
.B(n_872),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1326),
.B(n_879),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1436),
.A2(n_1188),
.B1(n_1191),
.B2(n_1179),
.Y(n_1503)
);

OR2x6_ASAP7_75t_L g1504 ( 
.A(n_1407),
.B(n_901),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1332),
.B(n_1008),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1300),
.B(n_880),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1370),
.A2(n_845),
.B1(n_848),
.B2(n_832),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1382),
.A2(n_849),
.B1(n_853),
.B2(n_850),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1368),
.B(n_884),
.C(n_882),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1447),
.B(n_887),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1317),
.Y(n_1512)
);

NOR3xp33_ASAP7_75t_L g1513 ( 
.A(n_1437),
.B(n_1054),
.C(n_949),
.Y(n_1513)
);

NOR3xp33_ASAP7_75t_L g1514 ( 
.A(n_1440),
.B(n_1393),
.C(n_1360),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1307),
.B(n_893),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1307),
.B(n_898),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1448),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1366),
.B(n_905),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1308),
.B(n_906),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1353),
.A2(n_862),
.B(n_867),
.C(n_859),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1343),
.B(n_909),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1385),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1383),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1308),
.B(n_912),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1382),
.B(n_913),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1440),
.B(n_1405),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1384),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1438),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1449),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1351),
.Y(n_1530)
);

OAI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1421),
.A2(n_830),
.B1(n_837),
.B2(n_833),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1334),
.B(n_918),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1313),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1334),
.B(n_923),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1335),
.B(n_924),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1354),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1316),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1361),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1363),
.B(n_935),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1372),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1375),
.B(n_937),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_SL g1542 ( 
.A(n_1418),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1377),
.B(n_938),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1394),
.B(n_940),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1411),
.B(n_941),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1411),
.A2(n_876),
.B1(n_877),
.B2(n_874),
.C(n_873),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1415),
.A2(n_945),
.B1(n_951),
.B2(n_943),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1299),
.B(n_954),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1389),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1302),
.B(n_956),
.Y(n_1550)
);

NOR3xp33_ASAP7_75t_L g1551 ( 
.A(n_1434),
.B(n_1059),
.C(n_1057),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1446),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1415),
.B(n_1072),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1389),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1401),
.B(n_964),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1401),
.B(n_1371),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1376),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1325),
.B(n_973),
.Y(n_1558)
);

BUFx4_ASAP7_75t_L g1559 ( 
.A(n_1418),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1373),
.B(n_1072),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1356),
.B(n_977),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1397),
.B(n_978),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1325),
.B(n_979),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1356),
.B(n_983),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1338),
.B(n_986),
.Y(n_1565)
);

NOR3xp33_ASAP7_75t_L g1566 ( 
.A(n_1364),
.B(n_1070),
.C(n_1061),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1400),
.A2(n_987),
.B1(n_996),
.B2(n_991),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1445),
.B(n_1297),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1445),
.B(n_998),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1435),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1416),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1379),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1338),
.A2(n_885),
.B(n_886),
.C(n_881),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1357),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1298),
.B(n_1079),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1357),
.Y(n_1576)
);

INVxp33_ASAP7_75t_L g1577 ( 
.A(n_1378),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1362),
.B(n_1441),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1381),
.Y(n_1579)
);

INVx4_ASAP7_75t_L g1580 ( 
.A(n_1318),
.Y(n_1580)
);

INVxp33_ASAP7_75t_L g1581 ( 
.A(n_1435),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1320),
.B(n_1002),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1320),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1311),
.B(n_1007),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1321),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1321),
.B(n_1011),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1322),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1309),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1314),
.A2(n_889),
.B(n_891),
.C(n_888),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1322),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1327),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1327),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1328),
.B(n_1079),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1328),
.B(n_1013),
.Y(n_1594)
);

OR2x6_ASAP7_75t_L g1595 ( 
.A(n_1314),
.B(n_950),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1311),
.B(n_1014),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1315),
.B(n_1021),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1315),
.B(n_1086),
.Y(n_1598)
);

AO21x2_ASAP7_75t_L g1599 ( 
.A1(n_1319),
.A2(n_931),
.B(n_844),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1408),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1408),
.B(n_1022),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1430),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1420),
.B(n_1102),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1420),
.B(n_1024),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1428),
.B(n_1025),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1428),
.B(n_1030),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1402),
.Y(n_1607)
);

NAND2xp33_ASAP7_75t_L g1608 ( 
.A(n_1402),
.B(n_1102),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1423),
.A2(n_896),
.B1(n_897),
.B2(n_894),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1426),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1402),
.B(n_1102),
.Y(n_1611)
);

NAND2xp33_ASAP7_75t_L g1612 ( 
.A(n_1433),
.B(n_1102),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1395),
.B(n_1031),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1403),
.B(n_1032),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1331),
.A2(n_1036),
.B1(n_1037),
.B2(n_1034),
.Y(n_1615)
);

OR2x6_ASAP7_75t_L g1616 ( 
.A(n_1336),
.B(n_1129),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1419),
.B(n_1044),
.Y(n_1617)
);

NAND2x1p5_ASAP7_75t_L g1618 ( 
.A(n_1337),
.B(n_1134),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1422),
.B(n_1045),
.Y(n_1619)
);

NOR3xp33_ASAP7_75t_L g1620 ( 
.A(n_1424),
.B(n_1154),
.C(n_1141),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1429),
.B(n_1047),
.Y(n_1621)
);

INVx4_ASAP7_75t_L g1622 ( 
.A(n_1404),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1339),
.A2(n_1049),
.B1(n_1051),
.B2(n_1048),
.Y(n_1623)
);

NOR3xp33_ASAP7_75t_L g1624 ( 
.A(n_1425),
.B(n_1060),
.C(n_1052),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1427),
.B(n_1063),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_L g1626 ( 
.A(n_1341),
.B(n_1069),
.C(n_1066),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1344),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1344),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1345),
.B(n_1071),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1346),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1347),
.A2(n_900),
.B(n_907),
.C(n_899),
.Y(n_1631)
);

O2A1O1Ixp5_ASAP7_75t_L g1632 ( 
.A1(n_1347),
.A2(n_864),
.B(n_868),
.C(n_858),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1348),
.A2(n_1076),
.B1(n_1077),
.B2(n_1074),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1349),
.B(n_1080),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1349),
.B(n_1081),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1355),
.B(n_1082),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1358),
.B(n_1083),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1359),
.B(n_1085),
.Y(n_1638)
);

OAI21xp33_ASAP7_75t_L g1639 ( 
.A1(n_1452),
.A2(n_1090),
.B(n_1089),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1471),
.B(n_960),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1512),
.B(n_796),
.Y(n_1641)
);

INVx4_ASAP7_75t_L g1642 ( 
.A(n_1504),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1586),
.B(n_1091),
.Y(n_1643)
);

O2A1O1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1458),
.A2(n_908),
.B(n_911),
.C(n_910),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1457),
.A2(n_914),
.B(n_921),
.C(n_920),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1632),
.A2(n_1414),
.B(n_1413),
.Y(n_1646)
);

OAI22x1_ASAP7_75t_L g1647 ( 
.A1(n_1567),
.A2(n_841),
.B1(n_842),
.B2(n_840),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1491),
.A2(n_922),
.B(n_932),
.C(n_928),
.Y(n_1648)
);

O2A1O1Ixp33_ASAP7_75t_L g1649 ( 
.A1(n_1520),
.A2(n_947),
.B(n_948),
.C(n_939),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1585),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1513),
.A2(n_1490),
.B1(n_1451),
.B2(n_1525),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1580),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1455),
.A2(n_962),
.B(n_961),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1568),
.A2(n_970),
.B(n_968),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1469),
.A2(n_972),
.B(n_976),
.C(n_971),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1457),
.A2(n_1578),
.B(n_1554),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1508),
.A2(n_990),
.B(n_989),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1495),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1549),
.A2(n_993),
.B(n_992),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1588),
.A2(n_1000),
.B(n_997),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1465),
.A2(n_1096),
.B1(n_1098),
.B2(n_1094),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1536),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1459),
.A2(n_1005),
.B(n_1004),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1540),
.A2(n_1006),
.B(n_1015),
.C(n_1012),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1456),
.B(n_1103),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1580),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1459),
.A2(n_1017),
.B(n_1028),
.C(n_1018),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1453),
.B(n_846),
.Y(n_1668)
);

NOR3xp33_ASAP7_75t_L g1669 ( 
.A(n_1531),
.B(n_1111),
.C(n_1107),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1461),
.B(n_861),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1556),
.A2(n_1035),
.B(n_1029),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1548),
.A2(n_1039),
.B(n_1038),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_1481),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1496),
.B(n_1114),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1466),
.B(n_1115),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1528),
.B(n_1189),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1550),
.A2(n_1053),
.B(n_1046),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1460),
.B(n_840),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1518),
.Y(n_1679)
);

AO21x1_ASAP7_75t_L g1680 ( 
.A1(n_1485),
.A2(n_1056),
.B(n_1055),
.Y(n_1680)
);

OAI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1470),
.A2(n_842),
.B1(n_919),
.B2(n_841),
.Y(n_1681)
);

AOI21xp33_ASAP7_75t_L g1682 ( 
.A1(n_1545),
.A2(n_1125),
.B(n_1121),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1454),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1504),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1507),
.B(n_1131),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1509),
.B(n_1133),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1547),
.B(n_1136),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1478),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1462),
.A2(n_934),
.B1(n_944),
.B2(n_919),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1515),
.B(n_1137),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1504),
.B(n_934),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1493),
.A2(n_1065),
.B(n_1064),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1464),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1523),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1589),
.A2(n_1075),
.B(n_1073),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1516),
.B(n_1138),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1573),
.A2(n_1097),
.B(n_1092),
.Y(n_1697)
);

INVx4_ASAP7_75t_L g1698 ( 
.A(n_1471),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1530),
.A2(n_1101),
.B(n_1100),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1471),
.Y(n_1700)
);

A2O1A1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1472),
.A2(n_1106),
.B(n_1108),
.C(n_1104),
.Y(n_1701)
);

CKINVDCx20_ASAP7_75t_R g1702 ( 
.A(n_1522),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1467),
.A2(n_1110),
.B(n_1109),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1583),
.A2(n_1116),
.B(n_1113),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1482),
.A2(n_1118),
.B(n_1117),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1510),
.B(n_895),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1587),
.A2(n_1126),
.B(n_1123),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1552),
.B(n_1142),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1488),
.A2(n_1130),
.B(n_1128),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1511),
.B(n_1143),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1479),
.Y(n_1711)
);

A2O1A1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1489),
.A2(n_1140),
.B(n_1144),
.C(n_1139),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1501),
.A2(n_955),
.B1(n_963),
.B2(n_944),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1502),
.A2(n_1148),
.B(n_1147),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1616),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1527),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1597),
.A2(n_1157),
.B(n_1150),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1506),
.A2(n_1162),
.B(n_1161),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1477),
.B(n_955),
.Y(n_1719)
);

OAI321xp33_ASAP7_75t_L g1720 ( 
.A1(n_1546),
.A2(n_1168),
.A3(n_1166),
.B1(n_1169),
.B2(n_1167),
.C(n_1163),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1514),
.A2(n_1474),
.B1(n_1626),
.B2(n_1497),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1526),
.B(n_1177),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1476),
.A2(n_1171),
.B(n_1170),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1607),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_L g1725 ( 
.A(n_1521),
.B(n_963),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1590),
.A2(n_1173),
.B(n_1172),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1480),
.A2(n_1180),
.B(n_1175),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1519),
.B(n_903),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1607),
.Y(n_1729)
);

OAI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1591),
.A2(n_1183),
.B(n_1181),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1592),
.A2(n_1192),
.B(n_1185),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1539),
.A2(n_1543),
.B(n_1541),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1544),
.A2(n_1196),
.B(n_967),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1475),
.B(n_1149),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1569),
.A2(n_967),
.B(n_966),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1616),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1607),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1486),
.B(n_1151),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1532),
.B(n_1152),
.Y(n_1739)
);

O2A1O1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1631),
.A2(n_994),
.B(n_1023),
.C(n_974),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1598),
.A2(n_1033),
.B1(n_1041),
.B2(n_1003),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1463),
.Y(n_1742)
);

OAI21xp33_ASAP7_75t_L g1743 ( 
.A1(n_1503),
.A2(n_1160),
.B(n_1159),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1494),
.B(n_1498),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1524),
.B(n_1155),
.Y(n_1745)
);

OA22x2_ASAP7_75t_L g1746 ( 
.A1(n_1570),
.A2(n_1033),
.B1(n_1041),
.B2(n_1003),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1500),
.B(n_1165),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_SL g1748 ( 
.A(n_1542),
.B(n_1050),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1561),
.B(n_904),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1582),
.A2(n_1095),
.B(n_1062),
.Y(n_1750)
);

OAI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1594),
.A2(n_1099),
.B(n_1095),
.Y(n_1751)
);

OAI21xp33_ASAP7_75t_L g1752 ( 
.A1(n_1499),
.A2(n_1067),
.B(n_1050),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1618),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1483),
.A2(n_1119),
.B(n_1099),
.Y(n_1754)
);

A2O1A1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1565),
.A2(n_1058),
.B(n_1176),
.C(n_988),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1534),
.B(n_1119),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1492),
.A2(n_1132),
.B(n_1122),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1535),
.B(n_1122),
.Y(n_1758)
);

NOR2x1p5_ASAP7_75t_SL g1759 ( 
.A(n_1602),
.B(n_1132),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1484),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1624),
.B(n_1067),
.Y(n_1761)
);

O2A1O1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1564),
.A2(n_1087),
.B(n_1190),
.C(n_1124),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1616),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1622),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1487),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1517),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1595),
.B(n_1068),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1595),
.Y(n_1768)
);

INVx4_ASAP7_75t_L g1769 ( 
.A(n_1473),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1574),
.A2(n_1193),
.B(n_1124),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1576),
.A2(n_1190),
.B(n_1087),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1566),
.A2(n_1194),
.B(n_1068),
.C(n_916),
.Y(n_1772)
);

A2O1A1Ixp33_ASAP7_75t_L g1773 ( 
.A1(n_1562),
.A2(n_1156),
.B(n_915),
.C(n_18),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1529),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1595),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1584),
.A2(n_20),
.B1(n_16),
.B2(n_19),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1596),
.B(n_20),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1555),
.B(n_21),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_SL g1779 ( 
.A(n_1542),
.B(n_1581),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1571),
.B(n_24),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1609),
.B(n_27),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1615),
.B(n_27),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1533),
.A2(n_1538),
.B(n_1537),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1634),
.A2(n_28),
.B(n_30),
.Y(n_1784)
);

AOI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1610),
.A2(n_28),
.B(n_31),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1557),
.A2(n_32),
.B(n_33),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1623),
.B(n_32),
.Y(n_1787)
);

OAI21xp33_ASAP7_75t_L g1788 ( 
.A1(n_1558),
.A2(n_34),
.B(n_35),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1563),
.B(n_771),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1473),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1635),
.A2(n_35),
.B(n_36),
.Y(n_1791)
);

BUFx6f_ASAP7_75t_L g1792 ( 
.A(n_1622),
.Y(n_1792)
);

OAI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1572),
.A2(n_37),
.B(n_38),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1636),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1637),
.A2(n_37),
.B(n_39),
.Y(n_1795)
);

AO21x1_ASAP7_75t_L g1796 ( 
.A1(n_1575),
.A2(n_40),
.B(n_41),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1551),
.B(n_778),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1638),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1620),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1633),
.B(n_43),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1577),
.B(n_44),
.Y(n_1801)
);

BUFx4f_ASAP7_75t_L g1802 ( 
.A(n_1559),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1601),
.B(n_45),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1579),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1604),
.B(n_48),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1605),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1600),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1606),
.B(n_769),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1599),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1505),
.A2(n_50),
.B(n_51),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1613),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1599),
.B(n_50),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1614),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1617),
.B(n_52),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1621),
.B(n_53),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1625),
.Y(n_1816)
);

NOR3xp33_ASAP7_75t_L g1817 ( 
.A(n_1619),
.B(n_53),
.C(n_54),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1629),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1560),
.B(n_58),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1630),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1593),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_R g1822 ( 
.A(n_1603),
.B(n_64),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1627),
.A2(n_66),
.B(n_67),
.Y(n_1823)
);

OR2x2_ASAP7_75t_SL g1824 ( 
.A(n_1628),
.B(n_69),
.Y(n_1824)
);

AND2x4_ASAP7_75t_SL g1825 ( 
.A(n_1611),
.B(n_766),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1608),
.B(n_768),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1612),
.B(n_71),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1585),
.Y(n_1828)
);

OAI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1468),
.A2(n_73),
.B(n_74),
.Y(n_1829)
);

CKINVDCx20_ASAP7_75t_R g1830 ( 
.A(n_1470),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1468),
.A2(n_75),
.B(n_76),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1452),
.B(n_75),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1468),
.A2(n_78),
.B(n_79),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1452),
.B(n_78),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1452),
.B(n_80),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1468),
.A2(n_81),
.B(n_82),
.Y(n_1836)
);

AO21x1_ASAP7_75t_L g1837 ( 
.A1(n_1553),
.A2(n_84),
.B(n_85),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1452),
.B(n_86),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1452),
.Y(n_1839)
);

AOI21x1_ASAP7_75t_L g1840 ( 
.A1(n_1457),
.A2(n_86),
.B(n_87),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1468),
.A2(n_87),
.B(n_88),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1580),
.Y(n_1842)
);

INVxp67_ASAP7_75t_L g1843 ( 
.A(n_1452),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1452),
.A2(n_92),
.B1(n_88),
.B2(n_89),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1580),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1452),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1512),
.B(n_768),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1452),
.B(n_89),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1585),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1468),
.A2(n_93),
.B(n_94),
.Y(n_1850)
);

NOR3xp33_ASAP7_75t_L g1851 ( 
.A(n_1531),
.B(n_95),
.C(n_96),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1452),
.B(n_95),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1452),
.B(n_97),
.Y(n_1853)
);

INVxp67_ASAP7_75t_SL g1854 ( 
.A(n_1452),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1468),
.A2(n_98),
.B(n_99),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1522),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1512),
.B(n_100),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1452),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1452),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1481),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1468),
.A2(n_105),
.B(n_106),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1453),
.B(n_767),
.Y(n_1862)
);

AO21x1_ASAP7_75t_L g1863 ( 
.A1(n_1553),
.A2(n_106),
.B(n_107),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1452),
.B(n_109),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1854),
.A2(n_113),
.B(n_115),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1843),
.B(n_115),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1732),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1839),
.B(n_118),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1846),
.B(n_119),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1651),
.B(n_119),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1662),
.B(n_121),
.Y(n_1871)
);

AOI21x1_ASAP7_75t_L g1872 ( 
.A1(n_1840),
.A2(n_122),
.B(n_123),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1656),
.A2(n_123),
.B(n_124),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1641),
.B(n_767),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1832),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1668),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1698),
.B(n_125),
.Y(n_1877)
);

AO31x2_ASAP7_75t_L g1878 ( 
.A1(n_1645),
.A2(n_129),
.A3(n_126),
.B(n_128),
.Y(n_1878)
);

A2O1A1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1653),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1659),
.B(n_130),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1802),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1830),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1834),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_1883)
);

AOI21xp33_ASAP7_75t_L g1884 ( 
.A1(n_1777),
.A2(n_138),
.B(n_139),
.Y(n_1884)
);

OAI21x1_ASAP7_75t_L g1885 ( 
.A1(n_1646),
.A2(n_140),
.B(n_143),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1657),
.B(n_144),
.Y(n_1886)
);

AO21x1_ASAP7_75t_L g1887 ( 
.A1(n_1829),
.A2(n_146),
.B(n_147),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1670),
.B(n_775),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1794),
.B(n_149),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1798),
.B(n_149),
.Y(n_1890)
);

INVxp67_ASAP7_75t_L g1891 ( 
.A(n_1748),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1698),
.B(n_150),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1811),
.B(n_151),
.Y(n_1893)
);

CKINVDCx11_ASAP7_75t_R g1894 ( 
.A(n_1702),
.Y(n_1894)
);

AOI221x1_ASAP7_75t_L g1895 ( 
.A1(n_1788),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.C(n_157),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1783),
.A2(n_155),
.B(n_156),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1673),
.A2(n_157),
.B(n_158),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1802),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_SL g1899 ( 
.A(n_1673),
.B(n_159),
.Y(n_1899)
);

AO31x2_ASAP7_75t_L g1900 ( 
.A1(n_1837),
.A2(n_163),
.A3(n_161),
.B(n_162),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1719),
.B(n_163),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1676),
.Y(n_1902)
);

AOI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1655),
.A2(n_168),
.B1(n_165),
.B2(n_167),
.C(n_169),
.Y(n_1903)
);

AOI21x1_ASAP7_75t_L g1904 ( 
.A1(n_1785),
.A2(n_171),
.B(n_173),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1813),
.B(n_173),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1699),
.A2(n_1703),
.B(n_1677),
.Y(n_1906)
);

A2O1A1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1644),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1692),
.A2(n_174),
.B(n_175),
.Y(n_1908)
);

O2A1O1Ixp33_ASAP7_75t_L g1909 ( 
.A1(n_1667),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1694),
.B(n_177),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1835),
.Y(n_1911)
);

A2O1A1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1740),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1652),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1716),
.B(n_181),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1664),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.C(n_187),
.Y(n_1915)
);

INVx5_ASAP7_75t_L g1916 ( 
.A(n_1642),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1672),
.A2(n_185),
.B(n_186),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1683),
.Y(n_1918)
);

A2O1A1Ixp33_ASAP7_75t_L g1919 ( 
.A1(n_1717),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_1919)
);

AO31x2_ASAP7_75t_L g1920 ( 
.A1(n_1863),
.A2(n_1755),
.A3(n_1818),
.B(n_1796),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1660),
.A2(n_190),
.B(n_191),
.Y(n_1921)
);

OAI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1671),
.A2(n_192),
.B(n_193),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1856),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1838),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1847),
.B(n_195),
.Y(n_1925)
);

OAI21x1_ASAP7_75t_SL g1926 ( 
.A1(n_1855),
.A2(n_195),
.B(n_196),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1679),
.B(n_196),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1862),
.B(n_197),
.Y(n_1928)
);

INVx6_ASAP7_75t_L g1929 ( 
.A(n_1769),
.Y(n_1929)
);

OA21x2_ASAP7_75t_L g1930 ( 
.A1(n_1823),
.A2(n_199),
.B(n_201),
.Y(n_1930)
);

AND2x6_ASAP7_75t_L g1931 ( 
.A(n_1736),
.B(n_199),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1753),
.B(n_202),
.Y(n_1932)
);

HAxp5_ASAP7_75t_L g1933 ( 
.A(n_1746),
.B(n_1681),
.CON(n_1933),
.SN(n_1933)
);

AO31x2_ASAP7_75t_L g1934 ( 
.A1(n_1735),
.A2(n_205),
.A3(n_203),
.B(n_204),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1693),
.B(n_204),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1860),
.A2(n_206),
.B(n_207),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1724),
.Y(n_1937)
);

AO31x2_ASAP7_75t_L g1938 ( 
.A1(n_1750),
.A2(n_210),
.A3(n_208),
.B(n_209),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1704),
.B(n_211),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1860),
.A2(n_212),
.B(n_213),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1652),
.Y(n_1941)
);

NAND2x1p5_ASAP7_75t_L g1942 ( 
.A(n_1642),
.B(n_213),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1767),
.B(n_764),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1767),
.B(n_765),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1806),
.B(n_216),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1666),
.Y(n_1946)
);

AOI21xp33_ASAP7_75t_L g1947 ( 
.A1(n_1803),
.A2(n_218),
.B(n_219),
.Y(n_1947)
);

AO31x2_ASAP7_75t_L g1948 ( 
.A1(n_1754),
.A2(n_221),
.A3(n_218),
.B(n_220),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1707),
.B(n_220),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1724),
.A2(n_223),
.B(n_224),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1691),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1769),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1715),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1678),
.B(n_225),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1741),
.B(n_227),
.Y(n_1955)
);

AOI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1729),
.A2(n_229),
.B(n_230),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1848),
.Y(n_1957)
);

OAI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1733),
.A2(n_1714),
.B(n_1654),
.Y(n_1958)
);

AO31x2_ASAP7_75t_L g1959 ( 
.A1(n_1757),
.A2(n_237),
.A3(n_231),
.B(n_233),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1729),
.A2(n_231),
.B(n_233),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1726),
.B(n_237),
.Y(n_1961)
);

INVx4_ASAP7_75t_L g1962 ( 
.A(n_1666),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1730),
.B(n_1718),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1728),
.B(n_238),
.Y(n_1964)
);

NAND3xp33_ASAP7_75t_L g1965 ( 
.A(n_1817),
.B(n_238),
.C(n_239),
.Y(n_1965)
);

NAND2x1p5_ASAP7_75t_L g1966 ( 
.A(n_1842),
.B(n_239),
.Y(n_1966)
);

INVx1_ASAP7_75t_SL g1967 ( 
.A(n_1842),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1723),
.B(n_240),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1845),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1727),
.B(n_243),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1729),
.A2(n_243),
.B(n_244),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1737),
.A2(n_244),
.B(n_246),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1663),
.B(n_247),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1857),
.B(n_248),
.Y(n_1974)
);

AND3x4_ASAP7_75t_L g1975 ( 
.A(n_1669),
.B(n_248),
.C(n_249),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1816),
.B(n_250),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1701),
.B(n_251),
.Y(n_1977)
);

INVxp67_ASAP7_75t_L g1978 ( 
.A(n_1713),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_R g1979 ( 
.A(n_1761),
.B(n_253),
.Y(n_1979)
);

BUFx2_ASAP7_75t_L g1980 ( 
.A(n_1684),
.Y(n_1980)
);

OAI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1852),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1712),
.B(n_256),
.Y(n_1982)
);

OAI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1864),
.A2(n_257),
.B(n_259),
.Y(n_1983)
);

OA21x2_ASAP7_75t_L g1984 ( 
.A1(n_1786),
.A2(n_257),
.B(n_260),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1737),
.A2(n_261),
.B(n_262),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1745),
.B(n_261),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1689),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1705),
.B(n_263),
.Y(n_1988)
);

NAND3xp33_ASAP7_75t_L g1989 ( 
.A(n_1721),
.B(n_1851),
.C(n_1793),
.Y(n_1989)
);

AOI21xp33_ASAP7_75t_L g1990 ( 
.A1(n_1805),
.A2(n_264),
.B(n_266),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1764),
.Y(n_1991)
);

AOI21x1_ASAP7_75t_L g1992 ( 
.A1(n_1814),
.A2(n_267),
.B(n_269),
.Y(n_1992)
);

AO31x2_ASAP7_75t_L g1993 ( 
.A1(n_1831),
.A2(n_271),
.A3(n_269),
.B(n_270),
.Y(n_1993)
);

OAI21xp5_ASAP7_75t_L g1994 ( 
.A1(n_1709),
.A2(n_270),
.B(n_271),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1658),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1751),
.B(n_1808),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1784),
.A2(n_276),
.B(n_273),
.C(n_274),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_SL g1998 ( 
.A1(n_1647),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1752),
.B(n_277),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1790),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1760),
.Y(n_2001)
);

A2O1A1Ixp33_ASAP7_75t_L g2002 ( 
.A1(n_1791),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_2002)
);

OAI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1833),
.A2(n_282),
.B(n_284),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1756),
.B(n_282),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1765),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1711),
.A2(n_287),
.B(n_288),
.Y(n_2006)
);

NAND2x1_ASAP7_75t_SL g2007 ( 
.A(n_1725),
.B(n_289),
.Y(n_2007)
);

OAI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1824),
.A2(n_1776),
.B1(n_1778),
.B2(n_1853),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1758),
.B(n_1731),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1685),
.B(n_291),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1686),
.B(n_292),
.Y(n_2011)
);

BUFx2_ASAP7_75t_L g2012 ( 
.A(n_1700),
.Y(n_2012)
);

NAND2x1p5_ASAP7_75t_L g2013 ( 
.A(n_1736),
.B(n_294),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1815),
.B(n_294),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1815),
.B(n_295),
.Y(n_2015)
);

OR2x6_ASAP7_75t_L g2016 ( 
.A(n_1780),
.B(n_780),
.Y(n_2016)
);

AO31x2_ASAP7_75t_L g2017 ( 
.A1(n_1836),
.A2(n_298),
.A3(n_296),
.B(n_297),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1688),
.Y(n_2018)
);

AOI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1749),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_2019)
);

NAND2x1p5_ASAP7_75t_L g2020 ( 
.A(n_1763),
.B(n_301),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1766),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1722),
.B(n_302),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1710),
.A2(n_305),
.B(n_306),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1747),
.B(n_308),
.Y(n_2024)
);

OAI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_1841),
.A2(n_309),
.B(n_310),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1768),
.B(n_311),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1774),
.Y(n_2027)
);

OAI22x1_ASAP7_75t_L g2028 ( 
.A1(n_1780),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_2028)
);

OAI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1850),
.A2(n_313),
.B(n_315),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1781),
.Y(n_2030)
);

AOI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1771),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_2031)
);

BUFx3_ASAP7_75t_L g2032 ( 
.A(n_1744),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1770),
.B(n_320),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1764),
.Y(n_2034)
);

AOI21xp33_ASAP7_75t_L g2035 ( 
.A1(n_1801),
.A2(n_322),
.B(n_323),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1734),
.A2(n_327),
.B(n_328),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1797),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1648),
.B(n_329),
.Y(n_2038)
);

OAI22x1_ASAP7_75t_L g2039 ( 
.A1(n_1812),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_SL g2040 ( 
.A(n_1711),
.B(n_330),
.Y(n_2040)
);

BUFx2_ASAP7_75t_SL g2041 ( 
.A(n_1764),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1643),
.B(n_331),
.Y(n_2042)
);

NOR2xp67_ASAP7_75t_L g2043 ( 
.A(n_1789),
.B(n_332),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1649),
.B(n_333),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1800),
.Y(n_2045)
);

INVx3_ASAP7_75t_L g2046 ( 
.A(n_1792),
.Y(n_2046)
);

OAI22x1_ASAP7_75t_L g2047 ( 
.A1(n_1812),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1650),
.B(n_336),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1828),
.B(n_337),
.Y(n_2049)
);

OAI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_1861),
.A2(n_338),
.B(n_339),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1661),
.B(n_338),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1849),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1792),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1807),
.Y(n_2054)
);

A2O1A1Ixp33_ASAP7_75t_L g2055 ( 
.A1(n_1795),
.A2(n_342),
.B(n_340),
.C(n_341),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1738),
.A2(n_344),
.B(n_346),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_1675),
.B(n_348),
.Y(n_2057)
);

INVx8_ASAP7_75t_L g2058 ( 
.A(n_1744),
.Y(n_2058)
);

NOR2x1_ASAP7_75t_SL g2059 ( 
.A(n_1711),
.B(n_350),
.Y(n_2059)
);

NAND3xp33_ASAP7_75t_SL g2060 ( 
.A(n_1799),
.B(n_351),
.C(n_352),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1690),
.B(n_354),
.Y(n_2061)
);

INVxp67_ASAP7_75t_SL g2062 ( 
.A(n_1762),
.Y(n_2062)
);

AOI21xp33_ASAP7_75t_L g2063 ( 
.A1(n_1782),
.A2(n_355),
.B(n_356),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1696),
.B(n_358),
.Y(n_2064)
);

AOI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_1739),
.A2(n_361),
.B(n_362),
.Y(n_2065)
);

A2O1A1Ixp33_ASAP7_75t_L g2066 ( 
.A1(n_1759),
.A2(n_1695),
.B(n_1787),
.C(n_1697),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1674),
.B(n_361),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1773),
.B(n_363),
.Y(n_2068)
);

NAND3xp33_ASAP7_75t_L g2069 ( 
.A(n_1640),
.B(n_365),
.C(n_366),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1687),
.A2(n_1708),
.B(n_1639),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1706),
.B(n_365),
.Y(n_2071)
);

OAI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1720),
.A2(n_366),
.B(n_368),
.Y(n_2072)
);

A2O1A1Ixp33_ASAP7_75t_L g2073 ( 
.A1(n_1682),
.A2(n_371),
.B(n_369),
.C(n_370),
.Y(n_2073)
);

AO31x2_ASAP7_75t_L g2074 ( 
.A1(n_1844),
.A2(n_373),
.A3(n_371),
.B(n_372),
.Y(n_2074)
);

OAI22x1_ASAP7_75t_L g2075 ( 
.A1(n_1640),
.A2(n_375),
.B1(n_372),
.B2(n_374),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1743),
.B(n_374),
.Y(n_2076)
);

AOI221xp5_ASAP7_75t_L g2077 ( 
.A1(n_1772),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.C(n_379),
.Y(n_2077)
);

BUFx3_ASAP7_75t_L g2078 ( 
.A(n_1742),
.Y(n_2078)
);

NAND2xp33_ASAP7_75t_L g2079 ( 
.A(n_1807),
.B(n_377),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1665),
.B(n_378),
.Y(n_2080)
);

AOI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1775),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.Y(n_2081)
);

A2O1A1Ixp33_ASAP7_75t_L g2082 ( 
.A1(n_1819),
.A2(n_387),
.B(n_384),
.C(n_386),
.Y(n_2082)
);

A2O1A1Ixp33_ASAP7_75t_L g2083 ( 
.A1(n_1810),
.A2(n_389),
.B(n_387),
.C(n_388),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1859),
.B(n_390),
.Y(n_2084)
);

NAND3x1_ASAP7_75t_L g2085 ( 
.A(n_1779),
.B(n_391),
.C(n_393),
.Y(n_2085)
);

AO21x2_ASAP7_75t_L g2086 ( 
.A1(n_1804),
.A2(n_391),
.B(n_393),
.Y(n_2086)
);

OAI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_1858),
.A2(n_394),
.B(n_395),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1820),
.B(n_398),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1822),
.Y(n_2089)
);

A2O1A1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_1827),
.A2(n_402),
.B(n_399),
.C(n_401),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1826),
.Y(n_2091)
);

OAI21x1_ASAP7_75t_L g2092 ( 
.A1(n_1821),
.A2(n_403),
.B(n_404),
.Y(n_2092)
);

NAND2x1p5_ASAP7_75t_L g2093 ( 
.A(n_1825),
.B(n_404),
.Y(n_2093)
);

AOI21x1_ASAP7_75t_L g2094 ( 
.A1(n_1840),
.A2(n_405),
.B(n_406),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_1846),
.Y(n_2095)
);

AOI21x1_ASAP7_75t_L g2096 ( 
.A1(n_1840),
.A2(n_408),
.B(n_409),
.Y(n_2096)
);

A2O1A1Ixp33_ASAP7_75t_L g2097 ( 
.A1(n_1732),
.A2(n_410),
.B(n_408),
.C(n_409),
.Y(n_2097)
);

NAND2x1p5_ASAP7_75t_L g2098 ( 
.A(n_1839),
.B(n_412),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_1854),
.A2(n_415),
.B(n_416),
.Y(n_2099)
);

AOI21x1_ASAP7_75t_L g2100 ( 
.A1(n_1840),
.A2(n_415),
.B(n_416),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1843),
.B(n_417),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1854),
.A2(n_420),
.B1(n_417),
.B2(n_418),
.Y(n_2102)
);

INVxp67_ASAP7_75t_SL g2103 ( 
.A(n_1854),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1846),
.Y(n_2104)
);

AOI21xp33_ASAP7_75t_L g2105 ( 
.A1(n_1777),
.A2(n_422),
.B(n_423),
.Y(n_2105)
);

BUFx12f_ASAP7_75t_L g2106 ( 
.A(n_1769),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1846),
.B(n_424),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_1854),
.A2(n_426),
.B(n_427),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1843),
.B(n_427),
.Y(n_2109)
);

A2O1A1Ixp33_ASAP7_75t_L g2110 ( 
.A1(n_1732),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_1843),
.B(n_428),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1843),
.B(n_431),
.Y(n_2112)
);

BUFx2_ASAP7_75t_L g2113 ( 
.A(n_1830),
.Y(n_2113)
);

OAI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_1732),
.A2(n_433),
.B(n_434),
.Y(n_2114)
);

OAI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_1732),
.A2(n_436),
.B(n_437),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_1843),
.B(n_436),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1846),
.B(n_438),
.Y(n_2117)
);

INVx3_ASAP7_75t_SL g2118 ( 
.A(n_1830),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1846),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1843),
.B(n_439),
.Y(n_2120)
);

BUFx2_ASAP7_75t_SL g2121 ( 
.A(n_1830),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1846),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_SL g2123 ( 
.A1(n_1854),
.A2(n_440),
.B(n_441),
.Y(n_2123)
);

O2A1O1Ixp33_ASAP7_75t_L g2124 ( 
.A1(n_1843),
.A2(n_443),
.B(n_441),
.C(n_442),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1839),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1839),
.B(n_442),
.Y(n_2126)
);

AO21x1_ASAP7_75t_L g2127 ( 
.A1(n_1840),
.A2(n_443),
.B(n_444),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1854),
.A2(n_445),
.B(n_446),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_1846),
.A2(n_448),
.B1(n_445),
.B2(n_447),
.Y(n_2129)
);

BUFx2_ASAP7_75t_L g2130 ( 
.A(n_1830),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1839),
.B(n_447),
.Y(n_2131)
);

OA21x2_ASAP7_75t_L g2132 ( 
.A1(n_1656),
.A2(n_448),
.B(n_449),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_1724),
.Y(n_2133)
);

BUFx4f_ASAP7_75t_L g2134 ( 
.A(n_1839),
.Y(n_2134)
);

NAND3xp33_ASAP7_75t_SL g2135 ( 
.A(n_1830),
.B(n_452),
.C(n_453),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_1846),
.B(n_452),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1854),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_1652),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1839),
.B(n_454),
.Y(n_2139)
);

BUFx4_ASAP7_75t_SL g2140 ( 
.A(n_1702),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_1854),
.A2(n_455),
.B(n_456),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_1846),
.B(n_457),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_1724),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1839),
.Y(n_2144)
);

AO21x1_ASAP7_75t_L g2145 ( 
.A1(n_1840),
.A2(n_458),
.B(n_459),
.Y(n_2145)
);

AOI21xp33_ASAP7_75t_L g2146 ( 
.A1(n_1777),
.A2(n_460),
.B(n_461),
.Y(n_2146)
);

O2A1O1Ixp5_ASAP7_75t_L g2147 ( 
.A1(n_1680),
.A2(n_468),
.B(n_464),
.C(n_466),
.Y(n_2147)
);

AOI221xp5_ASAP7_75t_L g2148 ( 
.A1(n_1655),
.A2(n_471),
.B1(n_466),
.B2(n_470),
.C(n_472),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1843),
.B(n_471),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1843),
.B(n_473),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1843),
.B(n_475),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1854),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1843),
.B(n_476),
.Y(n_2153)
);

A2O1A1Ixp33_ASAP7_75t_L g2154 ( 
.A1(n_1732),
.A2(n_480),
.B(n_478),
.C(n_479),
.Y(n_2154)
);

AOI21xp33_ASAP7_75t_L g2155 ( 
.A1(n_1777),
.A2(n_478),
.B(n_479),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1846),
.Y(n_2156)
);

AND2x2_ASAP7_75t_SL g2157 ( 
.A(n_1802),
.B(n_481),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1843),
.B(n_482),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1846),
.B(n_482),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1843),
.B(n_483),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_1652),
.Y(n_2161)
);

NAND2x1p5_ASAP7_75t_L g2162 ( 
.A(n_1839),
.B(n_484),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_1843),
.B(n_485),
.Y(n_2163)
);

O2A1O1Ixp5_ASAP7_75t_L g2164 ( 
.A1(n_1680),
.A2(n_488),
.B(n_486),
.C(n_487),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_1854),
.A2(n_486),
.B(n_488),
.Y(n_2165)
);

AO31x2_ASAP7_75t_L g2166 ( 
.A1(n_1809),
.A2(n_491),
.A3(n_489),
.B(n_490),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1839),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_1854),
.A2(n_492),
.B(n_493),
.Y(n_2168)
);

OAI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_1732),
.A2(n_493),
.B(n_494),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1846),
.Y(n_2170)
);

BUFx2_ASAP7_75t_L g2171 ( 
.A(n_1830),
.Y(n_2171)
);

A2O1A1Ixp33_ASAP7_75t_L g2172 ( 
.A1(n_1732),
.A2(n_497),
.B(n_494),
.C(n_496),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1843),
.B(n_497),
.Y(n_2173)
);

OAI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_1732),
.A2(n_498),
.B(n_499),
.Y(n_2174)
);

AOI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_1854),
.A2(n_499),
.B(n_500),
.Y(n_2175)
);

OAI21x1_ASAP7_75t_SL g2176 ( 
.A1(n_1698),
.A2(n_503),
.B(n_504),
.Y(n_2176)
);

OAI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_1732),
.A2(n_503),
.B(n_505),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1839),
.B(n_506),
.Y(n_2178)
);

HB1xp67_ASAP7_75t_L g2179 ( 
.A(n_1846),
.Y(n_2179)
);

AOI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_1854),
.A2(n_506),
.B(n_508),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1843),
.B(n_509),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1843),
.B(n_509),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1839),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1843),
.B(n_510),
.Y(n_2184)
);

INVx2_ASAP7_75t_SL g2185 ( 
.A(n_1846),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1843),
.B(n_511),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1843),
.B(n_512),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1846),
.Y(n_2188)
);

NOR2x1_ASAP7_75t_L g2189 ( 
.A(n_1769),
.B(n_513),
.Y(n_2189)
);

OAI21x1_ASAP7_75t_SL g2190 ( 
.A1(n_1698),
.A2(n_514),
.B(n_515),
.Y(n_2190)
);

AOI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_1854),
.A2(n_515),
.B(n_516),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_1854),
.A2(n_518),
.B(n_519),
.Y(n_2192)
);

AO21x1_ASAP7_75t_L g2193 ( 
.A1(n_1840),
.A2(n_519),
.B(n_520),
.Y(n_2193)
);

OAI22x1_ASAP7_75t_L g2194 ( 
.A1(n_1767),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_2194)
);

AO21x1_ASAP7_75t_L g2195 ( 
.A1(n_1840),
.A2(n_523),
.B(n_524),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_1741),
.B(n_525),
.Y(n_2196)
);

OAI21xp5_ASAP7_75t_L g2197 ( 
.A1(n_1732),
.A2(n_525),
.B(n_526),
.Y(n_2197)
);

A2O1A1Ixp33_ASAP7_75t_L g2198 ( 
.A1(n_1732),
.A2(n_528),
.B(n_526),
.C(n_527),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_1843),
.B(n_527),
.Y(n_2199)
);

BUFx4_ASAP7_75t_SL g2200 ( 
.A(n_1702),
.Y(n_2200)
);

AND2x4_ASAP7_75t_L g2201 ( 
.A(n_1843),
.B(n_530),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1846),
.B(n_531),
.Y(n_2202)
);

AOI21xp5_ASAP7_75t_L g2203 ( 
.A1(n_1854),
.A2(n_531),
.B(n_532),
.Y(n_2203)
);

OAI21xp5_ASAP7_75t_L g2204 ( 
.A1(n_1732),
.A2(n_533),
.B(n_534),
.Y(n_2204)
);

OAI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_1732),
.A2(n_535),
.B(n_537),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1843),
.B(n_538),
.Y(n_2206)
);

INVx3_ASAP7_75t_SL g2207 ( 
.A(n_1830),
.Y(n_2207)
);

INVxp67_ASAP7_75t_SL g2208 ( 
.A(n_1854),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_1846),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_1641),
.B(n_539),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1846),
.Y(n_2211)
);

OAI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_1732),
.A2(n_540),
.B(n_541),
.Y(n_2212)
);

HB1xp67_ASAP7_75t_L g2213 ( 
.A(n_1846),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1839),
.B(n_542),
.Y(n_2214)
);

AO21x1_ASAP7_75t_L g2215 ( 
.A1(n_1840),
.A2(n_543),
.B(n_544),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_L g2216 ( 
.A(n_1724),
.Y(n_2216)
);

AOI21x1_ASAP7_75t_L g2217 ( 
.A1(n_1840),
.A2(n_546),
.B(n_547),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1846),
.Y(n_2218)
);

AND2x4_ASAP7_75t_L g2219 ( 
.A(n_1843),
.B(n_550),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1839),
.B(n_552),
.Y(n_2220)
);

AND2x2_ASAP7_75t_SL g2221 ( 
.A(n_1802),
.B(n_554),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_1830),
.Y(n_2222)
);

AO21x2_ASAP7_75t_L g2223 ( 
.A1(n_1809),
.A2(n_555),
.B(n_556),
.Y(n_2223)
);

CKINVDCx16_ASAP7_75t_R g2224 ( 
.A(n_1830),
.Y(n_2224)
);

BUFx8_ASAP7_75t_SL g2225 ( 
.A(n_1802),
.Y(n_2225)
);

AOI221xp5_ASAP7_75t_SL g2226 ( 
.A1(n_1740),
.A2(n_558),
.B1(n_559),
.B2(n_560),
.C(n_561),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1846),
.B(n_558),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1843),
.B(n_561),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1843),
.B(n_562),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1846),
.Y(n_2230)
);

BUFx2_ASAP7_75t_L g2231 ( 
.A(n_1830),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_1724),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1846),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_1846),
.B(n_563),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_SL g2235 ( 
.A(n_1881),
.Y(n_2235)
);

OAI21x1_ASAP7_75t_SL g2236 ( 
.A1(n_1926),
.A2(n_564),
.B(n_565),
.Y(n_2236)
);

OA21x2_ASAP7_75t_L g2237 ( 
.A1(n_1885),
.A2(n_564),
.B(n_565),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2185),
.B(n_566),
.Y(n_2238)
);

AO21x2_ASAP7_75t_L g2239 ( 
.A1(n_2114),
.A2(n_566),
.B(n_567),
.Y(n_2239)
);

AO21x2_ASAP7_75t_L g2240 ( 
.A1(n_2114),
.A2(n_568),
.B(n_569),
.Y(n_2240)
);

AOI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_2103),
.A2(n_2208),
.B1(n_1987),
.B2(n_1902),
.Y(n_2241)
);

BUFx3_ASAP7_75t_L g2242 ( 
.A(n_2034),
.Y(n_2242)
);

INVx4_ASAP7_75t_L g2243 ( 
.A(n_2225),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_2134),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2125),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2144),
.B(n_571),
.Y(n_2246)
);

OAI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_2066),
.A2(n_573),
.B(n_574),
.Y(n_2247)
);

OR2x6_ASAP7_75t_L g2248 ( 
.A(n_2016),
.B(n_2121),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2167),
.B(n_2183),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_1989),
.B(n_575),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_1978),
.B(n_576),
.Y(n_2251)
);

AO21x1_ASAP7_75t_L g2252 ( 
.A1(n_2008),
.A2(n_2162),
.B(n_2098),
.Y(n_2252)
);

NAND2x1p5_ASAP7_75t_L g2253 ( 
.A(n_2134),
.B(n_578),
.Y(n_2253)
);

OAI21x1_ASAP7_75t_SL g2254 ( 
.A1(n_2115),
.A2(n_578),
.B(n_579),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2104),
.Y(n_2255)
);

AOI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_2070),
.A2(n_580),
.B(n_581),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2045),
.B(n_582),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1918),
.Y(n_2258)
);

BUFx8_ASAP7_75t_L g2259 ( 
.A(n_2113),
.Y(n_2259)
);

OA21x2_ASAP7_75t_L g2260 ( 
.A1(n_2169),
.A2(n_591),
.B(n_592),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2119),
.Y(n_2261)
);

BUFx2_ASAP7_75t_SL g2262 ( 
.A(n_1898),
.Y(n_2262)
);

INVx1_ASAP7_75t_SL g2263 ( 
.A(n_2095),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2122),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2156),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_SL g2266 ( 
.A1(n_2169),
.A2(n_593),
.B(n_594),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2170),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_2140),
.Y(n_2268)
);

OR2x6_ASAP7_75t_L g2269 ( 
.A(n_2016),
.B(n_1942),
.Y(n_2269)
);

CKINVDCx11_ASAP7_75t_R g2270 ( 
.A(n_2118),
.Y(n_2270)
);

OR2x6_ASAP7_75t_L g2271 ( 
.A(n_2016),
.B(n_594),
.Y(n_2271)
);

CKINVDCx20_ASAP7_75t_R g2272 ( 
.A(n_1894),
.Y(n_2272)
);

NAND2x1p5_ASAP7_75t_L g2273 ( 
.A(n_1916),
.B(n_595),
.Y(n_2273)
);

OR2x6_ASAP7_75t_L g2274 ( 
.A(n_1942),
.B(n_599),
.Y(n_2274)
);

AO21x2_ASAP7_75t_L g2275 ( 
.A1(n_2174),
.A2(n_600),
.B(n_601),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_1916),
.B(n_602),
.Y(n_2276)
);

OR2x6_ASAP7_75t_L g2277 ( 
.A(n_2106),
.B(n_602),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_2062),
.B(n_604),
.Y(n_2278)
);

NOR2xp33_ASAP7_75t_L g2279 ( 
.A(n_2188),
.B(n_606),
.Y(n_2279)
);

OAI21x1_ASAP7_75t_SL g2280 ( 
.A1(n_2174),
.A2(n_607),
.B(n_609),
.Y(n_2280)
);

AOI21x1_ASAP7_75t_L g2281 ( 
.A1(n_1872),
.A2(n_607),
.B(n_610),
.Y(n_2281)
);

AOI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2009),
.A2(n_610),
.B(n_611),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2211),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2005),
.Y(n_2284)
);

BUFx2_ASAP7_75t_SL g2285 ( 
.A(n_1916),
.Y(n_2285)
);

INVx3_ASAP7_75t_L g2286 ( 
.A(n_1962),
.Y(n_2286)
);

OA21x2_ASAP7_75t_L g2287 ( 
.A1(n_2177),
.A2(n_614),
.B(n_615),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_L g2288 ( 
.A1(n_1955),
.A2(n_616),
.B1(n_617),
.B2(n_618),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2179),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_1937),
.Y(n_2290)
);

AO21x2_ASAP7_75t_L g2291 ( 
.A1(n_2177),
.A2(n_617),
.B(n_619),
.Y(n_2291)
);

AOI221xp5_ASAP7_75t_L g2292 ( 
.A1(n_1888),
.A2(n_2077),
.B1(n_1944),
.B2(n_1943),
.C(n_2008),
.Y(n_2292)
);

AOI22xp33_ASAP7_75t_SL g2293 ( 
.A1(n_2157),
.A2(n_621),
.B1(n_622),
.B2(n_623),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2218),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2209),
.B(n_625),
.Y(n_2295)
);

OAI21xp5_ASAP7_75t_L g2296 ( 
.A1(n_1996),
.A2(n_626),
.B(n_627),
.Y(n_2296)
);

BUFx2_ASAP7_75t_L g2297 ( 
.A(n_2207),
.Y(n_2297)
);

AND2x4_ASAP7_75t_L g2298 ( 
.A(n_2230),
.B(n_629),
.Y(n_2298)
);

AOI21x1_ASAP7_75t_L g2299 ( 
.A1(n_2094),
.A2(n_631),
.B(n_634),
.Y(n_2299)
);

BUFx12f_ASAP7_75t_L g2300 ( 
.A(n_2130),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2213),
.B(n_631),
.Y(n_2301)
);

INVx3_ASAP7_75t_L g2302 ( 
.A(n_1962),
.Y(n_2302)
);

BUFx2_ASAP7_75t_R g2303 ( 
.A(n_2171),
.Y(n_2303)
);

INVxp67_ASAP7_75t_L g2304 ( 
.A(n_2111),
.Y(n_2304)
);

BUFx12f_ASAP7_75t_L g2305 ( 
.A(n_2222),
.Y(n_2305)
);

AOI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_1963),
.A2(n_638),
.B(n_639),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_2200),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2233),
.Y(n_2308)
);

BUFx2_ASAP7_75t_L g2309 ( 
.A(n_2231),
.Y(n_2309)
);

AOI21xp5_ASAP7_75t_L g2310 ( 
.A1(n_1958),
.A2(n_638),
.B(n_639),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1868),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2126),
.Y(n_2312)
);

OAI21xp5_ASAP7_75t_L g2313 ( 
.A1(n_1989),
.A2(n_641),
.B(n_642),
.Y(n_2313)
);

INVx4_ASAP7_75t_L g2314 ( 
.A(n_2058),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2126),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2131),
.Y(n_2316)
);

AO21x2_ASAP7_75t_L g2317 ( 
.A1(n_2197),
.A2(n_2205),
.B(n_2204),
.Y(n_2317)
);

AO31x2_ASAP7_75t_L g2318 ( 
.A1(n_2127),
.A2(n_2145),
.A3(n_2195),
.B(n_2193),
.Y(n_2318)
);

CKINVDCx20_ASAP7_75t_R g2319 ( 
.A(n_2224),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2131),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2139),
.Y(n_2321)
);

AND2x4_ASAP7_75t_L g2322 ( 
.A(n_1995),
.B(n_646),
.Y(n_2322)
);

AO21x2_ASAP7_75t_L g2323 ( 
.A1(n_2197),
.A2(n_647),
.B(n_649),
.Y(n_2323)
);

INVx8_ASAP7_75t_L g2324 ( 
.A(n_2058),
.Y(n_2324)
);

BUFx3_ASAP7_75t_L g2325 ( 
.A(n_2034),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_1899),
.B(n_650),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2139),
.Y(n_2327)
);

HB1xp67_ASAP7_75t_L g2328 ( 
.A(n_2034),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_2037),
.B(n_651),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2178),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2178),
.Y(n_2331)
);

INVxp67_ASAP7_75t_SL g2332 ( 
.A(n_2048),
.Y(n_2332)
);

OA21x2_ASAP7_75t_L g2333 ( 
.A1(n_2204),
.A2(n_652),
.B(n_653),
.Y(n_2333)
);

NAND2x1p5_ASAP7_75t_L g2334 ( 
.A(n_2053),
.B(n_652),
.Y(n_2334)
);

OAI21x1_ASAP7_75t_SL g2335 ( 
.A1(n_2205),
.A2(n_653),
.B(n_654),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2214),
.Y(n_2336)
);

OA21x2_ASAP7_75t_L g2337 ( 
.A1(n_2212),
.A2(n_654),
.B(n_655),
.Y(n_2337)
);

INVxp67_ASAP7_75t_SL g2338 ( 
.A(n_2048),
.Y(n_2338)
);

BUFx10_ASAP7_75t_L g2339 ( 
.A(n_1932),
.Y(n_2339)
);

OA21x2_ASAP7_75t_L g2340 ( 
.A1(n_2212),
.A2(n_659),
.B(n_661),
.Y(n_2340)
);

AO21x2_ASAP7_75t_L g2341 ( 
.A1(n_2096),
.A2(n_659),
.B(n_661),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2214),
.Y(n_2342)
);

INVx5_ASAP7_75t_L g2343 ( 
.A(n_2053),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2021),
.Y(n_2344)
);

OAI21xp5_ASAP7_75t_L g2345 ( 
.A1(n_2030),
.A2(n_1958),
.B(n_1906),
.Y(n_2345)
);

BUFx12f_ASAP7_75t_L g2346 ( 
.A(n_1923),
.Y(n_2346)
);

OA21x2_ASAP7_75t_L g2347 ( 
.A1(n_1895),
.A2(n_662),
.B(n_663),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_L g2348 ( 
.A1(n_2100),
.A2(n_664),
.B(n_665),
.Y(n_2348)
);

INVx2_ASAP7_75t_SL g2349 ( 
.A(n_2058),
.Y(n_2349)
);

CKINVDCx20_ASAP7_75t_R g2350 ( 
.A(n_1882),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_1899),
.B(n_666),
.Y(n_2351)
);

NAND3xp33_ASAP7_75t_L g2352 ( 
.A(n_2226),
.B(n_667),
.C(n_668),
.Y(n_2352)
);

AOI22xp33_ASAP7_75t_L g2353 ( 
.A1(n_2060),
.A2(n_667),
.B1(n_668),
.B2(n_669),
.Y(n_2353)
);

BUFx3_ASAP7_75t_L g2354 ( 
.A(n_2053),
.Y(n_2354)
);

NAND3xp33_ASAP7_75t_L g2355 ( 
.A(n_2226),
.B(n_669),
.C(n_671),
.Y(n_2355)
);

NAND2x1p5_ASAP7_75t_L g2356 ( 
.A(n_1877),
.B(n_671),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_1991),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2220),
.Y(n_2358)
);

AO21x2_ASAP7_75t_L g2359 ( 
.A1(n_2217),
.A2(n_672),
.B(n_674),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2220),
.Y(n_2360)
);

BUFx12f_ASAP7_75t_L g2361 ( 
.A(n_1929),
.Y(n_2361)
);

INVxp67_ASAP7_75t_SL g2362 ( 
.A(n_2049),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_1901),
.B(n_675),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1910),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1910),
.Y(n_2365)
);

NAND2x1p5_ASAP7_75t_L g2366 ( 
.A(n_1877),
.B(n_676),
.Y(n_2366)
);

AO21x2_ASAP7_75t_L g2367 ( 
.A1(n_2215),
.A2(n_676),
.B(n_677),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_1933),
.B(n_679),
.Y(n_2368)
);

INVx8_ASAP7_75t_L g2369 ( 
.A(n_1931),
.Y(n_2369)
);

BUFx2_ASAP7_75t_SL g2370 ( 
.A(n_1932),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1914),
.Y(n_2371)
);

AO21x2_ASAP7_75t_L g2372 ( 
.A1(n_1887),
.A2(n_682),
.B(n_683),
.Y(n_2372)
);

AND2x4_ASAP7_75t_L g2373 ( 
.A(n_2001),
.B(n_682),
.Y(n_2373)
);

CKINVDCx6p67_ASAP7_75t_R g2374 ( 
.A(n_2221),
.Y(n_2374)
);

AND2x4_ASAP7_75t_L g2375 ( 
.A(n_2027),
.B(n_683),
.Y(n_2375)
);

OAI222xp33_ASAP7_75t_L g2376 ( 
.A1(n_2137),
.A2(n_685),
.B1(n_686),
.B2(n_688),
.C1(n_689),
.C2(n_690),
.Y(n_2376)
);

HB1xp67_ASAP7_75t_L g2377 ( 
.A(n_1945),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1914),
.Y(n_2378)
);

INVx2_ASAP7_75t_SL g2379 ( 
.A(n_1929),
.Y(n_2379)
);

HB1xp67_ASAP7_75t_L g2380 ( 
.A(n_1945),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_2196),
.A2(n_2111),
.B1(n_2163),
.B2(n_2116),
.Y(n_2381)
);

BUFx3_ASAP7_75t_L g2382 ( 
.A(n_1991),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_1875),
.A2(n_688),
.B(n_689),
.Y(n_2383)
);

INVx6_ASAP7_75t_L g2384 ( 
.A(n_2000),
.Y(n_2384)
);

AND2x4_ASAP7_75t_L g2385 ( 
.A(n_2091),
.B(n_692),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1889),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2089),
.B(n_2107),
.Y(n_2387)
);

BUFx2_ASAP7_75t_SL g2388 ( 
.A(n_1931),
.Y(n_2388)
);

AND2x4_ASAP7_75t_L g2389 ( 
.A(n_2117),
.B(n_693),
.Y(n_2389)
);

BUFx2_ASAP7_75t_SL g2390 ( 
.A(n_1931),
.Y(n_2390)
);

AO21x2_ASAP7_75t_L g2391 ( 
.A1(n_1904),
.A2(n_693),
.B(n_694),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1889),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_2136),
.B(n_695),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_1911),
.B(n_696),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2142),
.B(n_2159),
.Y(n_2395)
);

AOI21x1_ASAP7_75t_L g2396 ( 
.A1(n_1992),
.A2(n_697),
.B(n_699),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_1924),
.B(n_699),
.Y(n_2397)
);

BUFx2_ASAP7_75t_L g2398 ( 
.A(n_2018),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1890),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_1890),
.Y(n_2400)
);

NAND2x1_ASAP7_75t_L g2401 ( 
.A(n_2133),
.B(n_700),
.Y(n_2401)
);

OAI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_1906),
.A2(n_700),
.B(n_701),
.Y(n_2402)
);

INVx1_ASAP7_75t_SL g2403 ( 
.A(n_2041),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1893),
.Y(n_2404)
);

OA21x2_ASAP7_75t_L g2405 ( 
.A1(n_1915),
.A2(n_703),
.B(n_704),
.Y(n_2405)
);

NAND4xp25_ASAP7_75t_L g2406 ( 
.A(n_1998),
.B(n_708),
.C(n_709),
.D(n_710),
.Y(n_2406)
);

AO21x2_ASAP7_75t_L g2407 ( 
.A1(n_1873),
.A2(n_708),
.B(n_710),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_1951),
.B(n_712),
.Y(n_2408)
);

NAND2x1p5_ASAP7_75t_L g2409 ( 
.A(n_2046),
.B(n_712),
.Y(n_2409)
);

A2O1A1Ixp33_ASAP7_75t_L g2410 ( 
.A1(n_2087),
.A2(n_713),
.B(n_715),
.C(n_716),
.Y(n_2410)
);

AO21x2_ASAP7_75t_L g2411 ( 
.A1(n_2003),
.A2(n_713),
.B(n_716),
.Y(n_2411)
);

AO21x2_ASAP7_75t_L g2412 ( 
.A1(n_2003),
.A2(n_717),
.B(n_718),
.Y(n_2412)
);

INVx6_ASAP7_75t_L g2413 ( 
.A(n_2032),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2202),
.B(n_717),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1893),
.Y(n_2415)
);

OAI21x1_ASAP7_75t_SL g2416 ( 
.A1(n_2087),
.A2(n_719),
.B(n_721),
.Y(n_2416)
);

BUFx3_ASAP7_75t_L g2417 ( 
.A(n_2046),
.Y(n_2417)
);

INVxp33_ASAP7_75t_L g2418 ( 
.A(n_1979),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_1957),
.A2(n_722),
.B(n_723),
.Y(n_2419)
);

INVx6_ASAP7_75t_L g2420 ( 
.A(n_2078),
.Y(n_2420)
);

INVx2_ASAP7_75t_SL g2421 ( 
.A(n_2116),
.Y(n_2421)
);

INVx1_ASAP7_75t_SL g2422 ( 
.A(n_1967),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_1905),
.Y(n_2423)
);

AO21x1_ASAP7_75t_L g2424 ( 
.A1(n_2098),
.A2(n_724),
.B(n_726),
.Y(n_2424)
);

AO31x2_ASAP7_75t_L g2425 ( 
.A1(n_1867),
.A2(n_727),
.A3(n_730),
.B(n_731),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2057),
.B(n_730),
.Y(n_2426)
);

AO31x2_ASAP7_75t_L g2427 ( 
.A1(n_2097),
.A2(n_731),
.A3(n_733),
.B(n_734),
.Y(n_2427)
);

INVx6_ASAP7_75t_SL g2428 ( 
.A(n_2163),
.Y(n_2428)
);

BUFx3_ASAP7_75t_L g2429 ( 
.A(n_2143),
.Y(n_2429)
);

BUFx8_ASAP7_75t_L g2430 ( 
.A(n_2012),
.Y(n_2430)
);

AO21x2_ASAP7_75t_L g2431 ( 
.A1(n_2025),
.A2(n_736),
.B(n_737),
.Y(n_2431)
);

OA21x2_ASAP7_75t_L g2432 ( 
.A1(n_1915),
.A2(n_738),
.B(n_739),
.Y(n_2432)
);

AOI21xp33_ASAP7_75t_L g2433 ( 
.A1(n_1870),
.A2(n_738),
.B(n_740),
.Y(n_2433)
);

NOR2xp67_ASAP7_75t_SL g2434 ( 
.A(n_2123),
.B(n_741),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_1905),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2162),
.Y(n_2436)
);

OAI22xp33_ASAP7_75t_L g2437 ( 
.A1(n_2137),
.A2(n_741),
.B1(n_743),
.B2(n_744),
.Y(n_2437)
);

INVx2_ASAP7_75t_SL g2438 ( 
.A(n_2199),
.Y(n_2438)
);

NOR2x1p5_ASAP7_75t_L g2439 ( 
.A(n_2199),
.B(n_745),
.Y(n_2439)
);

BUFx2_ASAP7_75t_L g2440 ( 
.A(n_1931),
.Y(n_2440)
);

BUFx3_ASAP7_75t_L g2441 ( 
.A(n_2216),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_1976),
.B(n_747),
.Y(n_2442)
);

CKINVDCx8_ASAP7_75t_R g2443 ( 
.A(n_2201),
.Y(n_2443)
);

OR2x6_ASAP7_75t_L g2444 ( 
.A(n_2201),
.B(n_748),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_2216),
.Y(n_2445)
);

OAI21x1_ASAP7_75t_SL g2446 ( 
.A1(n_1983),
.A2(n_749),
.B(n_751),
.Y(n_2446)
);

NAND3xp33_ASAP7_75t_L g2447 ( 
.A(n_1965),
.B(n_751),
.C(n_752),
.Y(n_2447)
);

BUFx3_ASAP7_75t_L g2448 ( 
.A(n_2232),
.Y(n_2448)
);

AND2x4_ASAP7_75t_L g2449 ( 
.A(n_2227),
.B(n_752),
.Y(n_2449)
);

INVx4_ASAP7_75t_L g2450 ( 
.A(n_1966),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2234),
.B(n_753),
.Y(n_2451)
);

AO21x2_ASAP7_75t_L g2452 ( 
.A1(n_2025),
.A2(n_755),
.B(n_756),
.Y(n_2452)
);

BUFx12f_ASAP7_75t_L g2453 ( 
.A(n_1952),
.Y(n_2453)
);

OAI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_2010),
.A2(n_755),
.B(n_756),
.Y(n_2454)
);

CKINVDCx14_ASAP7_75t_R g2455 ( 
.A(n_2219),
.Y(n_2455)
);

INVx4_ASAP7_75t_L g2456 ( 
.A(n_1966),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2219),
.B(n_759),
.Y(n_2457)
);

AOI21xp5_ASAP7_75t_L g2458 ( 
.A1(n_2061),
.A2(n_760),
.B(n_761),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_1913),
.B(n_760),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2011),
.B(n_761),
.Y(n_2460)
);

OAI21x1_ASAP7_75t_SL g2461 ( 
.A1(n_1983),
.A2(n_763),
.B(n_765),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_1967),
.Y(n_2462)
);

OR2x6_ASAP7_75t_L g2463 ( 
.A(n_2093),
.B(n_2013),
.Y(n_2463)
);

BUFx2_ASAP7_75t_L g2464 ( 
.A(n_1891),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2013),
.Y(n_2465)
);

CKINVDCx20_ASAP7_75t_R g2466 ( 
.A(n_1953),
.Y(n_2466)
);

BUFx12f_ASAP7_75t_L g2467 ( 
.A(n_2093),
.Y(n_2467)
);

INVx6_ASAP7_75t_L g2468 ( 
.A(n_2080),
.Y(n_2468)
);

BUFx6f_ASAP7_75t_L g2469 ( 
.A(n_2054),
.Y(n_2469)
);

OAI21x1_ASAP7_75t_L g2470 ( 
.A1(n_2054),
.A2(n_770),
.B(n_771),
.Y(n_2470)
);

OA21x2_ASAP7_75t_L g2471 ( 
.A1(n_2029),
.A2(n_772),
.B(n_773),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2020),
.Y(n_2472)
);

INVx6_ASAP7_75t_L g2473 ( 
.A(n_2080),
.Y(n_2473)
);

CKINVDCx20_ASAP7_75t_R g2474 ( 
.A(n_1980),
.Y(n_2474)
);

OAI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2014),
.A2(n_777),
.B1(n_779),
.B2(n_2015),
.Y(n_2475)
);

BUFx3_ASAP7_75t_L g2476 ( 
.A(n_1913),
.Y(n_2476)
);

BUFx12f_ASAP7_75t_L g2477 ( 
.A(n_1954),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_1908),
.Y(n_2478)
);

BUFx3_ASAP7_75t_L g2479 ( 
.A(n_1941),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2028),
.Y(n_2480)
);

BUFx10_ASAP7_75t_L g2481 ( 
.A(n_2022),
.Y(n_2481)
);

NOR2xp67_ASAP7_75t_L g2482 ( 
.A(n_2194),
.B(n_2039),
.Y(n_2482)
);

CKINVDCx20_ASAP7_75t_R g2483 ( 
.A(n_2052),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_1871),
.Y(n_2484)
);

AO21x2_ASAP7_75t_L g2485 ( 
.A1(n_2029),
.A2(n_2050),
.B(n_2223),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_1941),
.Y(n_2486)
);

INVx3_ASAP7_75t_L g2487 ( 
.A(n_1946),
.Y(n_2487)
);

OAI21x1_ASAP7_75t_L g2488 ( 
.A1(n_2033),
.A2(n_2132),
.B(n_2050),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_1935),
.Y(n_2489)
);

BUFx2_ASAP7_75t_SL g2490 ( 
.A(n_2043),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2223),
.Y(n_2491)
);

INVx8_ASAP7_75t_L g2492 ( 
.A(n_1946),
.Y(n_2492)
);

INVx3_ASAP7_75t_SL g2493 ( 
.A(n_1892),
.Y(n_2493)
);

AOI21x1_ASAP7_75t_L g2494 ( 
.A1(n_1930),
.A2(n_1984),
.B(n_2011),
.Y(n_2494)
);

INVx1_ASAP7_75t_SL g2495 ( 
.A(n_2040),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2088),
.Y(n_2496)
);

BUFx2_ASAP7_75t_L g2497 ( 
.A(n_2007),
.Y(n_2497)
);

INVx3_ASAP7_75t_L g2498 ( 
.A(n_1969),
.Y(n_2498)
);

INVx3_ASAP7_75t_L g2499 ( 
.A(n_1969),
.Y(n_2499)
);

INVxp67_ASAP7_75t_L g2500 ( 
.A(n_1869),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2088),
.Y(n_2501)
);

AND2x4_ASAP7_75t_L g2502 ( 
.A(n_2138),
.B(n_2161),
.Y(n_2502)
);

AOI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2064),
.A2(n_2004),
.B(n_2067),
.Y(n_2503)
);

NAND2x1p5_ASAP7_75t_L g2504 ( 
.A(n_2138),
.B(n_2161),
.Y(n_2504)
);

OAI21x1_ASAP7_75t_L g2505 ( 
.A1(n_1950),
.A2(n_1960),
.B(n_1956),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2026),
.Y(n_2506)
);

OAI21x1_ASAP7_75t_L g2507 ( 
.A1(n_1971),
.A2(n_1985),
.B(n_1972),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2026),
.Y(n_2508)
);

OAI21x1_ASAP7_75t_L g2509 ( 
.A1(n_1896),
.A2(n_1940),
.B(n_1936),
.Y(n_2509)
);

OAI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2147),
.A2(n_2164),
.B(n_2154),
.Y(n_2510)
);

OA21x2_ASAP7_75t_L g2511 ( 
.A1(n_2110),
.A2(n_2198),
.B(n_2172),
.Y(n_2511)
);

BUFx2_ASAP7_75t_SL g2512 ( 
.A(n_2085),
.Y(n_2512)
);

AOI22xp33_ASAP7_75t_L g2513 ( 
.A1(n_2068),
.A2(n_2044),
.B1(n_2038),
.B2(n_1975),
.Y(n_2513)
);

INVx4_ASAP7_75t_L g2514 ( 
.A(n_2051),
.Y(n_2514)
);

BUFx3_ASAP7_75t_L g2515 ( 
.A(n_2014),
.Y(n_2515)
);

BUFx3_ASAP7_75t_L g2516 ( 
.A(n_2015),
.Y(n_2516)
);

BUFx3_ASAP7_75t_L g2517 ( 
.A(n_2092),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_1986),
.B(n_2101),
.Y(n_2518)
);

BUFx2_ASAP7_75t_L g2519 ( 
.A(n_1922),
.Y(n_2519)
);

HB1xp67_ASAP7_75t_L g2520 ( 
.A(n_2072),
.Y(n_2520)
);

OAI21xp5_ASAP7_75t_L g2521 ( 
.A1(n_1880),
.A2(n_1949),
.B(n_1939),
.Y(n_2521)
);

OR2x6_ASAP7_75t_L g2522 ( 
.A(n_2006),
.B(n_1897),
.Y(n_2522)
);

NOR2xp33_ASAP7_75t_L g2523 ( 
.A(n_2112),
.B(n_2120),
.Y(n_2523)
);

OAI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_1961),
.A2(n_1886),
.B(n_1973),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2042),
.B(n_2149),
.Y(n_2525)
);

INVx5_ASAP7_75t_SL g2526 ( 
.A(n_2086),
.Y(n_2526)
);

BUFx8_ASAP7_75t_SL g2527 ( 
.A(n_2068),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_1878),
.Y(n_2528)
);

CKINVDCx20_ASAP7_75t_R g2529 ( 
.A(n_1876),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_1878),
.Y(n_2530)
);

AOI22x1_ASAP7_75t_L g2531 ( 
.A1(n_2065),
.A2(n_2056),
.B1(n_2036),
.B2(n_2023),
.Y(n_2531)
);

INVx2_ASAP7_75t_SL g2532 ( 
.A(n_2189),
.Y(n_2532)
);

AOI21x1_ASAP7_75t_L g2533 ( 
.A1(n_1974),
.A2(n_2076),
.B(n_1925),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_1878),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2150),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2151),
.B(n_2153),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2158),
.B(n_2160),
.Y(n_2537)
);

OAI22xp5_ASAP7_75t_L g2538 ( 
.A1(n_1965),
.A2(n_1981),
.B1(n_1883),
.B2(n_2044),
.Y(n_2538)
);

OAI21x1_ASAP7_75t_SL g2539 ( 
.A1(n_2059),
.A2(n_2072),
.B(n_2190),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_2176),
.Y(n_2540)
);

AND2x4_ASAP7_75t_L g2541 ( 
.A(n_1964),
.B(n_2173),
.Y(n_2541)
);

INVx1_ASAP7_75t_SL g2542 ( 
.A(n_2040),
.Y(n_2542)
);

INVx1_ASAP7_75t_SL g2543 ( 
.A(n_2181),
.Y(n_2543)
);

OA21x2_ASAP7_75t_L g2544 ( 
.A1(n_1917),
.A2(n_1912),
.B(n_1921),
.Y(n_2544)
);

AOI21xp33_ASAP7_75t_L g2545 ( 
.A1(n_2071),
.A2(n_2124),
.B(n_2086),
.Y(n_2545)
);

AOI21x1_ASAP7_75t_L g2546 ( 
.A1(n_2076),
.A2(n_2071),
.B(n_2084),
.Y(n_2546)
);

HB1xp67_ASAP7_75t_L g2547 ( 
.A(n_1917),
.Y(n_2547)
);

OR2x6_ASAP7_75t_L g2548 ( 
.A(n_2047),
.B(n_1865),
.Y(n_2548)
);

AO21x2_ASAP7_75t_L g2549 ( 
.A1(n_1884),
.A2(n_2105),
.B(n_2155),
.Y(n_2549)
);

OR2x6_ASAP7_75t_L g2550 ( 
.A(n_2099),
.B(n_2108),
.Y(n_2550)
);

INVx2_ASAP7_75t_SL g2551 ( 
.A(n_2182),
.Y(n_2551)
);

BUFx6f_ASAP7_75t_L g2552 ( 
.A(n_1968),
.Y(n_2552)
);

NAND3xp33_ASAP7_75t_L g2553 ( 
.A(n_1907),
.B(n_2002),
.C(n_2055),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2184),
.Y(n_2554)
);

OAI21xp5_ASAP7_75t_L g2555 ( 
.A1(n_1970),
.A2(n_2180),
.B(n_2165),
.Y(n_2555)
);

AO21x2_ASAP7_75t_L g2556 ( 
.A1(n_1884),
.A2(n_2105),
.B(n_2155),
.Y(n_2556)
);

OAI21x1_ASAP7_75t_L g2557 ( 
.A1(n_2128),
.A2(n_2191),
.B(n_2141),
.Y(n_2557)
);

AO21x2_ASAP7_75t_L g2558 ( 
.A1(n_2146),
.A2(n_1994),
.B(n_2035),
.Y(n_2558)
);

HB1xp67_ASAP7_75t_L g2559 ( 
.A(n_1883),
.Y(n_2559)
);

BUFx6f_ASAP7_75t_L g2560 ( 
.A(n_1988),
.Y(n_2560)
);

BUFx6f_ASAP7_75t_L g2561 ( 
.A(n_2187),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2255),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2258),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2245),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2284),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2261),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2344),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2264),
.Y(n_2568)
);

BUFx3_ASAP7_75t_L g2569 ( 
.A(n_2324),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2265),
.Y(n_2570)
);

OAI21x1_ASAP7_75t_SL g2571 ( 
.A1(n_2252),
.A2(n_1981),
.B(n_2168),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2267),
.Y(n_2572)
);

AOI22xp33_ASAP7_75t_L g2573 ( 
.A1(n_2482),
.A2(n_2135),
.B1(n_1999),
.B2(n_2069),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2283),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2294),
.Y(n_2575)
);

NAND2x1p5_ASAP7_75t_L g2576 ( 
.A(n_2314),
.B(n_1866),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2324),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2369),
.Y(n_2578)
);

AO21x2_ASAP7_75t_L g2579 ( 
.A1(n_2494),
.A2(n_1990),
.B(n_1947),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2308),
.Y(n_2580)
);

CKINVDCx5p33_ASAP7_75t_R g2581 ( 
.A(n_2268),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2249),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2249),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2246),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2394),
.Y(n_2585)
);

BUFx12f_ASAP7_75t_L g2586 ( 
.A(n_2270),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2394),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_2529),
.A2(n_2069),
.B1(n_1947),
.B2(n_2075),
.Y(n_2588)
);

OAI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2271),
.A2(n_2081),
.B1(n_2102),
.B2(n_2152),
.Y(n_2589)
);

CKINVDCx20_ASAP7_75t_R g2590 ( 
.A(n_2272),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2271),
.B(n_1874),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2397),
.Y(n_2592)
);

AOI22xp33_ASAP7_75t_L g2593 ( 
.A1(n_2529),
.A2(n_1903),
.B1(n_2148),
.B2(n_2063),
.Y(n_2593)
);

BUFx2_ASAP7_75t_L g2594 ( 
.A(n_2483),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2397),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2373),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2373),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2375),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2375),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2322),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2369),
.Y(n_2601)
);

AO21x2_ASAP7_75t_L g2602 ( 
.A1(n_2345),
.A2(n_1990),
.B(n_2063),
.Y(n_2602)
);

INVx4_ASAP7_75t_L g2603 ( 
.A(n_2324),
.Y(n_2603)
);

OAI22xp33_ASAP7_75t_L g2604 ( 
.A1(n_2271),
.A2(n_2019),
.B1(n_1982),
.B2(n_1977),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2322),
.Y(n_2605)
);

OR2x6_ASAP7_75t_L g2606 ( 
.A(n_2369),
.B(n_2192),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2257),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2257),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2279),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2279),
.Y(n_2610)
);

BUFx2_ASAP7_75t_L g2611 ( 
.A(n_2483),
.Y(n_2611)
);

HB1xp67_ASAP7_75t_L g2612 ( 
.A(n_2462),
.Y(n_2612)
);

INVx4_ASAP7_75t_L g2613 ( 
.A(n_2361),
.Y(n_2613)
);

HB1xp67_ASAP7_75t_L g2614 ( 
.A(n_2462),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2385),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2385),
.Y(n_2616)
);

BUFx10_ASAP7_75t_L g2617 ( 
.A(n_2268),
.Y(n_2617)
);

OAI22xp33_ASAP7_75t_L g2618 ( 
.A1(n_2444),
.A2(n_2229),
.B1(n_2228),
.B2(n_1928),
.Y(n_2618)
);

CKINVDCx20_ASAP7_75t_R g2619 ( 
.A(n_2272),
.Y(n_2619)
);

AOI21x1_ASAP7_75t_L g2620 ( 
.A1(n_2546),
.A2(n_2533),
.B(n_2491),
.Y(n_2620)
);

OAI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_2538),
.A2(n_2203),
.B(n_2175),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2298),
.Y(n_2622)
);

INVx8_ASAP7_75t_L g2623 ( 
.A(n_2274),
.Y(n_2623)
);

INVx2_ASAP7_75t_SL g2624 ( 
.A(n_2384),
.Y(n_2624)
);

HB1xp67_ASAP7_75t_L g2625 ( 
.A(n_2332),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2455),
.B(n_2210),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2455),
.B(n_2024),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2298),
.Y(n_2628)
);

BUFx2_ASAP7_75t_R g2629 ( 
.A(n_2307),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2444),
.B(n_1927),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2450),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2356),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2467),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2356),
.Y(n_2634)
);

CKINVDCx14_ASAP7_75t_R g2635 ( 
.A(n_2307),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2366),
.Y(n_2636)
);

OAI22xp33_ASAP7_75t_L g2637 ( 
.A1(n_2444),
.A2(n_2206),
.B1(n_2186),
.B2(n_2109),
.Y(n_2637)
);

AO21x2_ASAP7_75t_L g2638 ( 
.A1(n_2345),
.A2(n_2545),
.B(n_2247),
.Y(n_2638)
);

BUFx3_ASAP7_75t_L g2639 ( 
.A(n_2384),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2366),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2514),
.B(n_2457),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2274),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2514),
.B(n_2031),
.Y(n_2643)
);

HB1xp67_ASAP7_75t_L g2644 ( 
.A(n_2332),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2274),
.Y(n_2645)
);

INVx3_ASAP7_75t_SL g2646 ( 
.A(n_2248),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2450),
.Y(n_2647)
);

OAI22xp5_ASAP7_75t_L g2648 ( 
.A1(n_2381),
.A2(n_2129),
.B1(n_2073),
.B2(n_2090),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2381),
.A2(n_1879),
.B1(n_2082),
.B2(n_1919),
.Y(n_2649)
);

BUFx2_ASAP7_75t_L g2650 ( 
.A(n_2430),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2238),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2253),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2253),
.Y(n_2653)
);

BUFx2_ASAP7_75t_L g2654 ( 
.A(n_2430),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2459),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2559),
.A2(n_2292),
.B1(n_2513),
.B2(n_2374),
.Y(n_2656)
);

CKINVDCx6p67_ASAP7_75t_R g2657 ( 
.A(n_2277),
.Y(n_2657)
);

INVx3_ASAP7_75t_L g2658 ( 
.A(n_2456),
.Y(n_2658)
);

OAI22xp33_ASAP7_75t_L g2659 ( 
.A1(n_2269),
.A2(n_2074),
.B1(n_2166),
.B2(n_2017),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2370),
.B(n_2166),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2459),
.Y(n_2661)
);

HB1xp67_ASAP7_75t_L g2662 ( 
.A(n_2338),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2273),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2273),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2409),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_2338),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2409),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2276),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2276),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2439),
.B(n_2166),
.Y(n_2670)
);

BUFx3_ASAP7_75t_L g2671 ( 
.A(n_2384),
.Y(n_2671)
);

HB1xp67_ASAP7_75t_L g2672 ( 
.A(n_2362),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_2270),
.Y(n_2673)
);

INVx2_ASAP7_75t_SL g2674 ( 
.A(n_2420),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2263),
.B(n_2074),
.Y(n_2675)
);

INVx3_ASAP7_75t_L g2676 ( 
.A(n_2456),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2295),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2301),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2286),
.Y(n_2679)
);

OAI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_2538),
.A2(n_1997),
.B(n_2083),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2377),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2377),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2380),
.Y(n_2683)
);

NAND2x1p5_ASAP7_75t_L g2684 ( 
.A(n_2244),
.B(n_2343),
.Y(n_2684)
);

INVx2_ASAP7_75t_SL g2685 ( 
.A(n_2420),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2263),
.B(n_2074),
.Y(n_2686)
);

INVxp67_ASAP7_75t_SL g2687 ( 
.A(n_2362),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2380),
.Y(n_2688)
);

OAI222xp33_ASAP7_75t_L g2689 ( 
.A1(n_2269),
.A2(n_1909),
.B1(n_2017),
.B2(n_1993),
.C1(n_1900),
.C2(n_1948),
.Y(n_2689)
);

BUFx2_ASAP7_75t_L g2690 ( 
.A(n_2269),
.Y(n_2690)
);

AOI22xp33_ASAP7_75t_L g2691 ( 
.A1(n_2559),
.A2(n_2079),
.B1(n_2017),
.B2(n_1993),
.Y(n_2691)
);

INVx2_ASAP7_75t_SL g2692 ( 
.A(n_2420),
.Y(n_2692)
);

OAI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2443),
.A2(n_1948),
.B1(n_1959),
.B2(n_1934),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2463),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2463),
.Y(n_2695)
);

AO21x2_ASAP7_75t_L g2696 ( 
.A1(n_2545),
.A2(n_1920),
.B(n_1900),
.Y(n_2696)
);

AND2x4_ASAP7_75t_L g2697 ( 
.A(n_2463),
.B(n_1920),
.Y(n_2697)
);

BUFx2_ASAP7_75t_L g2698 ( 
.A(n_2474),
.Y(n_2698)
);

OR2x2_ASAP7_75t_L g2699 ( 
.A(n_2289),
.B(n_1959),
.Y(n_2699)
);

NAND3xp33_ASAP7_75t_L g2700 ( 
.A(n_2352),
.B(n_1900),
.C(n_1934),
.Y(n_2700)
);

INVx2_ASAP7_75t_SL g2701 ( 
.A(n_2453),
.Y(n_2701)
);

BUFx2_ASAP7_75t_SL g2702 ( 
.A(n_2235),
.Y(n_2702)
);

BUFx2_ASAP7_75t_L g2703 ( 
.A(n_2474),
.Y(n_2703)
);

INVx2_ASAP7_75t_SL g2704 ( 
.A(n_2339),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2496),
.Y(n_2705)
);

HB1xp67_ASAP7_75t_L g2706 ( 
.A(n_2422),
.Y(n_2706)
);

BUFx12f_ASAP7_75t_SL g2707 ( 
.A(n_2277),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2501),
.Y(n_2708)
);

OAI21xp5_ASAP7_75t_L g2709 ( 
.A1(n_2352),
.A2(n_1938),
.B(n_2355),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2251),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_2319),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2289),
.B(n_1938),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2251),
.Y(n_2713)
);

BUFx6f_ASAP7_75t_L g2714 ( 
.A(n_2290),
.Y(n_2714)
);

INVx3_ASAP7_75t_L g2715 ( 
.A(n_2286),
.Y(n_2715)
);

INVx6_ASAP7_75t_L g2716 ( 
.A(n_2259),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2368),
.Y(n_2717)
);

INVx2_ASAP7_75t_SL g2718 ( 
.A(n_2339),
.Y(n_2718)
);

HB1xp67_ASAP7_75t_L g2719 ( 
.A(n_2328),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2395),
.B(n_2293),
.Y(n_2720)
);

INVx3_ASAP7_75t_L g2721 ( 
.A(n_2302),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2408),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2293),
.B(n_2363),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2241),
.B(n_2408),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2311),
.B(n_2312),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2315),
.B(n_2316),
.Y(n_2726)
);

INVx6_ASAP7_75t_L g2727 ( 
.A(n_2259),
.Y(n_2727)
);

HB1xp67_ASAP7_75t_L g2728 ( 
.A(n_2328),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2424),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2470),
.Y(n_2730)
);

HB1xp67_ASAP7_75t_L g2731 ( 
.A(n_2547),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_L g2732 ( 
.A1(n_2513),
.A2(n_2406),
.B1(n_2480),
.B2(n_2527),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2414),
.Y(n_2733)
);

BUFx3_ASAP7_75t_L g2734 ( 
.A(n_2343),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2437),
.Y(n_2735)
);

NAND2x1p5_ASAP7_75t_L g2736 ( 
.A(n_2244),
.B(n_2343),
.Y(n_2736)
);

BUFx2_ASAP7_75t_L g2737 ( 
.A(n_2428),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2436),
.Y(n_2738)
);

BUFx2_ASAP7_75t_L g2739 ( 
.A(n_2428),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2389),
.B(n_2393),
.Y(n_2740)
);

BUFx3_ASAP7_75t_L g2741 ( 
.A(n_2343),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_L g2742 ( 
.A1(n_2406),
.A2(n_2480),
.B1(n_2527),
.B2(n_2248),
.Y(n_2742)
);

AO21x2_ASAP7_75t_L g2743 ( 
.A1(n_2247),
.A2(n_2530),
.B(n_2528),
.Y(n_2743)
);

NAND2x1_ASAP7_75t_L g2744 ( 
.A(n_2440),
.B(n_2254),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_L g2745 ( 
.A1(n_2248),
.A2(n_2278),
.B1(n_2519),
.B2(n_2518),
.Y(n_2745)
);

AO21x2_ASAP7_75t_L g2746 ( 
.A1(n_2534),
.A2(n_2478),
.B(n_2488),
.Y(n_2746)
);

HB1xp67_ASAP7_75t_L g2747 ( 
.A(n_2547),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2285),
.Y(n_2748)
);

AOI22xp33_ASAP7_75t_L g2749 ( 
.A1(n_2278),
.A2(n_2518),
.B1(n_2313),
.B2(n_2523),
.Y(n_2749)
);

INVx3_ASAP7_75t_L g2750 ( 
.A(n_2302),
.Y(n_2750)
);

OR2x6_ASAP7_75t_L g2751 ( 
.A(n_2388),
.B(n_2390),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_2319),
.Y(n_2752)
);

BUFx12f_ASAP7_75t_L g2753 ( 
.A(n_2243),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2389),
.B(n_2393),
.Y(n_2754)
);

BUFx2_ASAP7_75t_L g2755 ( 
.A(n_2466),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_2492),
.Y(n_2756)
);

AOI21x1_ASAP7_75t_L g2757 ( 
.A1(n_2503),
.A2(n_2250),
.B(n_2520),
.Y(n_2757)
);

INVx2_ASAP7_75t_SL g2758 ( 
.A(n_2346),
.Y(n_2758)
);

INVxp67_ASAP7_75t_L g2759 ( 
.A(n_2398),
.Y(n_2759)
);

BUFx3_ASAP7_75t_L g2760 ( 
.A(n_2349),
.Y(n_2760)
);

CKINVDCx6p67_ASAP7_75t_R g2761 ( 
.A(n_2277),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2475),
.Y(n_2762)
);

AOI21x1_ASAP7_75t_L g2763 ( 
.A1(n_2503),
.A2(n_2250),
.B(n_2520),
.Y(n_2763)
);

NAND3xp33_ASAP7_75t_L g2764 ( 
.A(n_2355),
.B(n_2447),
.C(n_2531),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2485),
.Y(n_2765)
);

AND2x2_ASAP7_75t_L g2766 ( 
.A(n_2449),
.B(n_2451),
.Y(n_2766)
);

OAI221xp5_ASAP7_75t_L g2767 ( 
.A1(n_2313),
.A2(n_2410),
.B1(n_2353),
.B2(n_2500),
.C(n_2288),
.Y(n_2767)
);

INVx3_ASAP7_75t_L g2768 ( 
.A(n_2492),
.Y(n_2768)
);

OR2x6_ASAP7_75t_L g2769 ( 
.A(n_2468),
.B(n_2473),
.Y(n_2769)
);

OAI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2304),
.A2(n_2473),
.B1(n_2468),
.B2(n_2475),
.Y(n_2770)
);

BUFx3_ASAP7_75t_L g2771 ( 
.A(n_2492),
.Y(n_2771)
);

AOI22xp33_ASAP7_75t_L g2772 ( 
.A1(n_2523),
.A2(n_2541),
.B1(n_2548),
.B2(n_2473),
.Y(n_2772)
);

NAND2x1p5_ASAP7_75t_L g2773 ( 
.A(n_2403),
.B(n_2495),
.Y(n_2773)
);

INVx3_ASAP7_75t_L g2774 ( 
.A(n_2242),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2449),
.Y(n_2775)
);

BUFx3_ASAP7_75t_L g2776 ( 
.A(n_2242),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2325),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2541),
.A2(n_2548),
.B1(n_2468),
.B2(n_2321),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2296),
.Y(n_2779)
);

BUFx2_ASAP7_75t_SL g2780 ( 
.A(n_2235),
.Y(n_2780)
);

BUFx3_ASAP7_75t_L g2781 ( 
.A(n_2325),
.Y(n_2781)
);

OAI21xp5_ASAP7_75t_L g2782 ( 
.A1(n_2553),
.A2(n_2510),
.B(n_2521),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2296),
.Y(n_2783)
);

INVx3_ASAP7_75t_L g2784 ( 
.A(n_2354),
.Y(n_2784)
);

NOR2xp33_ASAP7_75t_L g2785 ( 
.A(n_2304),
.B(n_2418),
.Y(n_2785)
);

CKINVDCx11_ASAP7_75t_R g2786 ( 
.A(n_2300),
.Y(n_2786)
);

AO21x2_ASAP7_75t_L g2787 ( 
.A1(n_2266),
.A2(n_2335),
.B(n_2280),
.Y(n_2787)
);

NAND2x1p5_ASAP7_75t_L g2788 ( 
.A(n_2403),
.B(n_2495),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2329),
.B(n_2421),
.Y(n_2789)
);

CKINVDCx11_ASAP7_75t_R g2790 ( 
.A(n_2305),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2460),
.Y(n_2791)
);

AO21x1_ASAP7_75t_L g2792 ( 
.A1(n_2310),
.A2(n_2402),
.B(n_2334),
.Y(n_2792)
);

AND2x4_ASAP7_75t_L g2793 ( 
.A(n_2465),
.B(n_2472),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_2354),
.Y(n_2794)
);

CKINVDCx11_ASAP7_75t_R g2795 ( 
.A(n_2243),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2460),
.Y(n_2796)
);

BUFx3_ASAP7_75t_L g2797 ( 
.A(n_2429),
.Y(n_2797)
);

BUFx8_ASAP7_75t_L g2798 ( 
.A(n_2297),
.Y(n_2798)
);

OR2x2_ASAP7_75t_L g2799 ( 
.A(n_2438),
.B(n_2309),
.Y(n_2799)
);

INVx6_ASAP7_75t_L g2800 ( 
.A(n_2413),
.Y(n_2800)
);

BUFx12f_ASAP7_75t_L g2801 ( 
.A(n_2464),
.Y(n_2801)
);

OR2x6_ASAP7_75t_L g2802 ( 
.A(n_2512),
.B(n_2326),
.Y(n_2802)
);

INVx3_ASAP7_75t_L g2803 ( 
.A(n_2504),
.Y(n_2803)
);

AOI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_2548),
.A2(n_2327),
.B1(n_2330),
.B2(n_2320),
.Y(n_2804)
);

INVx3_ASAP7_75t_L g2805 ( 
.A(n_2504),
.Y(n_2805)
);

INVx3_ASAP7_75t_L g2806 ( 
.A(n_2382),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2485),
.Y(n_2807)
);

OAI22xp33_ASAP7_75t_L g2808 ( 
.A1(n_2418),
.A2(n_2402),
.B1(n_2493),
.B2(n_2454),
.Y(n_2808)
);

CKINVDCx5p33_ASAP7_75t_R g2809 ( 
.A(n_2303),
.Y(n_2809)
);

INVx3_ASAP7_75t_L g2810 ( 
.A(n_2382),
.Y(n_2810)
);

BUFx2_ASAP7_75t_L g2811 ( 
.A(n_2466),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2282),
.Y(n_2812)
);

AO21x1_ASAP7_75t_L g2813 ( 
.A1(n_2310),
.A2(n_2334),
.B(n_2256),
.Y(n_2813)
);

HB1xp67_ASAP7_75t_L g2814 ( 
.A(n_2317),
.Y(n_2814)
);

INVx3_ASAP7_75t_L g2815 ( 
.A(n_2417),
.Y(n_2815)
);

AOI22xp33_ASAP7_75t_L g2816 ( 
.A1(n_2331),
.A2(n_2336),
.B1(n_2435),
.B2(n_2342),
.Y(n_2816)
);

OAI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2410),
.A2(n_2542),
.B1(n_2515),
.B2(n_2516),
.Y(n_2817)
);

OAI22xp5_ASAP7_75t_SL g2818 ( 
.A1(n_2350),
.A2(n_2329),
.B1(n_2477),
.B2(n_2493),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2497),
.Y(n_2819)
);

BUFx2_ASAP7_75t_L g2820 ( 
.A(n_2350),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2358),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2360),
.Y(n_2822)
);

HB1xp67_ASAP7_75t_L g2823 ( 
.A(n_2317),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2386),
.Y(n_2824)
);

BUFx3_ASAP7_75t_L g2825 ( 
.A(n_2429),
.Y(n_2825)
);

AOI22xp33_ASAP7_75t_SL g2826 ( 
.A1(n_2416),
.A2(n_2461),
.B1(n_2446),
.B2(n_2333),
.Y(n_2826)
);

AO21x1_ASAP7_75t_SL g2827 ( 
.A1(n_2376),
.A2(n_2288),
.B(n_2353),
.Y(n_2827)
);

HB1xp67_ASAP7_75t_L g2828 ( 
.A(n_2515),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2392),
.Y(n_2829)
);

CKINVDCx5p33_ASAP7_75t_R g2830 ( 
.A(n_2303),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2399),
.Y(n_2831)
);

AOI22xp33_ASAP7_75t_L g2832 ( 
.A1(n_2400),
.A2(n_2415),
.B1(n_2404),
.B2(n_2423),
.Y(n_2832)
);

AOI22xp33_ASAP7_75t_SL g2833 ( 
.A1(n_2260),
.A2(n_2340),
.B1(n_2337),
.B2(n_2333),
.Y(n_2833)
);

BUFx2_ASAP7_75t_L g2834 ( 
.A(n_2413),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2506),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2508),
.Y(n_2836)
);

INVx1_ASAP7_75t_SL g2837 ( 
.A(n_2417),
.Y(n_2837)
);

BUFx2_ASAP7_75t_L g2838 ( 
.A(n_2413),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2396),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_2262),
.Y(n_2840)
);

AOI22xp33_ASAP7_75t_SL g2841 ( 
.A1(n_2260),
.A2(n_2340),
.B1(n_2337),
.B2(n_2287),
.Y(n_2841)
);

OAI21x1_ASAP7_75t_L g2842 ( 
.A1(n_2505),
.A2(n_2507),
.B(n_2509),
.Y(n_2842)
);

CKINVDCx6p67_ASAP7_75t_R g2843 ( 
.A(n_2387),
.Y(n_2843)
);

AOI22xp33_ASAP7_75t_L g2844 ( 
.A1(n_2364),
.A2(n_2378),
.B1(n_2371),
.B2(n_2365),
.Y(n_2844)
);

BUFx6f_ASAP7_75t_SL g2845 ( 
.A(n_2387),
.Y(n_2845)
);

BUFx2_ASAP7_75t_L g2846 ( 
.A(n_2623),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2562),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2766),
.B(n_2426),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2566),
.Y(n_2849)
);

OR2x2_ASAP7_75t_L g2850 ( 
.A(n_2594),
.B(n_2516),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2568),
.Y(n_2851)
);

BUFx2_ASAP7_75t_L g2852 ( 
.A(n_2623),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2563),
.Y(n_2853)
);

HB1xp67_ASAP7_75t_L g2854 ( 
.A(n_2625),
.Y(n_2854)
);

INVx3_ASAP7_75t_L g2855 ( 
.A(n_2751),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2740),
.B(n_2754),
.Y(n_2856)
);

AND2x4_ASAP7_75t_L g2857 ( 
.A(n_2751),
.B(n_2540),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2717),
.B(n_2426),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2570),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2564),
.Y(n_2860)
);

INVx3_ASAP7_75t_L g2861 ( 
.A(n_2751),
.Y(n_2861)
);

HB1xp67_ASAP7_75t_L g2862 ( 
.A(n_2625),
.Y(n_2862)
);

BUFx2_ASAP7_75t_L g2863 ( 
.A(n_2623),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2565),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2567),
.Y(n_2865)
);

BUFx2_ASAP7_75t_L g2866 ( 
.A(n_2840),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2641),
.B(n_2500),
.Y(n_2867)
);

OR2x2_ASAP7_75t_L g2868 ( 
.A(n_2611),
.B(n_2543),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2572),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2733),
.B(n_2535),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2720),
.B(n_2554),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2574),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2789),
.B(n_2442),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2677),
.B(n_2442),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2678),
.B(n_2532),
.Y(n_2875)
);

INVx3_ASAP7_75t_L g2876 ( 
.A(n_2734),
.Y(n_2876)
);

BUFx3_ASAP7_75t_L g2877 ( 
.A(n_2577),
.Y(n_2877)
);

BUFx8_ASAP7_75t_L g2878 ( 
.A(n_2633),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2843),
.B(n_2543),
.Y(n_2879)
);

CKINVDCx5p33_ASAP7_75t_R g2880 ( 
.A(n_2707),
.Y(n_2880)
);

BUFx3_ASAP7_75t_L g2881 ( 
.A(n_2577),
.Y(n_2881)
);

INVx3_ASAP7_75t_L g2882 ( 
.A(n_2734),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2651),
.B(n_2379),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2575),
.Y(n_2884)
);

INVxp67_ASAP7_75t_L g2885 ( 
.A(n_2644),
.Y(n_2885)
);

AOI22xp33_ASAP7_75t_L g2886 ( 
.A1(n_2656),
.A2(n_2553),
.B1(n_2484),
.B2(n_2489),
.Y(n_2886)
);

BUFx2_ASAP7_75t_SL g2887 ( 
.A(n_2603),
.Y(n_2887)
);

INVx1_ASAP7_75t_SL g2888 ( 
.A(n_2837),
.Y(n_2888)
);

AND2x4_ASAP7_75t_L g2889 ( 
.A(n_2697),
.B(n_2540),
.Y(n_2889)
);

AOI22xp5_ASAP7_75t_L g2890 ( 
.A1(n_2656),
.A2(n_2434),
.B1(n_2551),
.B2(n_2481),
.Y(n_2890)
);

AOI22xp33_ASAP7_75t_L g2891 ( 
.A1(n_2732),
.A2(n_2827),
.B1(n_2749),
.B2(n_2742),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2741),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2580),
.Y(n_2893)
);

INVx3_ASAP7_75t_L g2894 ( 
.A(n_2741),
.Y(n_2894)
);

INVx3_ASAP7_75t_L g2895 ( 
.A(n_2578),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2724),
.B(n_2458),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2578),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2821),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2760),
.B(n_2458),
.Y(n_2899)
);

BUFx3_ASAP7_75t_L g2900 ( 
.A(n_2577),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2582),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2760),
.B(n_2476),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2697),
.B(n_2517),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2822),
.Y(n_2904)
);

INVx1_ASAP7_75t_SL g2905 ( 
.A(n_2837),
.Y(n_2905)
);

HB1xp67_ASAP7_75t_L g2906 ( 
.A(n_2662),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2626),
.B(n_2476),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2627),
.B(n_2479),
.Y(n_2908)
);

BUFx2_ASAP7_75t_L g2909 ( 
.A(n_2840),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2698),
.B(n_2479),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2824),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2703),
.B(n_2357),
.Y(n_2912)
);

AND2x4_ASAP7_75t_L g2913 ( 
.A(n_2694),
.B(n_2517),
.Y(n_2913)
);

BUFx3_ASAP7_75t_L g2914 ( 
.A(n_2569),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2759),
.B(n_2357),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2583),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2829),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2831),
.Y(n_2918)
);

CKINVDCx5p33_ASAP7_75t_R g2919 ( 
.A(n_2657),
.Y(n_2919)
);

CKINVDCx14_ASAP7_75t_R g2920 ( 
.A(n_2635),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2835),
.Y(n_2921)
);

AND2x4_ASAP7_75t_L g2922 ( 
.A(n_2695),
.B(n_2441),
.Y(n_2922)
);

BUFx2_ASAP7_75t_L g2923 ( 
.A(n_2631),
.Y(n_2923)
);

HB1xp67_ASAP7_75t_L g2924 ( 
.A(n_2662),
.Y(n_2924)
);

HB1xp67_ASAP7_75t_L g2925 ( 
.A(n_2666),
.Y(n_2925)
);

INVx2_ASAP7_75t_SL g2926 ( 
.A(n_2716),
.Y(n_2926)
);

AOI22xp33_ASAP7_75t_SL g2927 ( 
.A1(n_2723),
.A2(n_2526),
.B1(n_2287),
.B2(n_2239),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2759),
.B(n_2502),
.Y(n_2928)
);

HB1xp67_ASAP7_75t_L g2929 ( 
.A(n_2666),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2722),
.B(n_2502),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2755),
.B(n_2383),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2836),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2705),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2811),
.B(n_2383),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2639),
.B(n_2419),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2708),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2639),
.B(n_2419),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2725),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2762),
.B(n_2558),
.Y(n_2939)
);

HB1xp67_ASAP7_75t_L g2940 ( 
.A(n_2672),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2725),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2726),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2726),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2671),
.B(n_2433),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2671),
.B(n_2433),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2738),
.Y(n_2946)
);

INVx3_ASAP7_75t_SL g2947 ( 
.A(n_2603),
.Y(n_2947)
);

BUFx6f_ASAP7_75t_L g2948 ( 
.A(n_2569),
.Y(n_2948)
);

NOR2x1p5_ASAP7_75t_L g2949 ( 
.A(n_2761),
.B(n_2809),
.Y(n_2949)
);

AOI22xp33_ASAP7_75t_L g2950 ( 
.A1(n_2732),
.A2(n_2525),
.B1(n_2537),
.B2(n_2536),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2612),
.Y(n_2951)
);

BUFx3_ASAP7_75t_L g2952 ( 
.A(n_2771),
.Y(n_2952)
);

HB1xp67_ASAP7_75t_L g2953 ( 
.A(n_2672),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2748),
.B(n_2490),
.Y(n_2954)
);

BUFx3_ASAP7_75t_L g2955 ( 
.A(n_2771),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2612),
.Y(n_2956)
);

OAI22xp5_ASAP7_75t_L g2957 ( 
.A1(n_2749),
.A2(n_2542),
.B1(n_2447),
.B2(n_2471),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2785),
.B(n_2372),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2785),
.B(n_2372),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_L g2960 ( 
.A1(n_2742),
.A2(n_2525),
.B1(n_2537),
.B2(n_2536),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2614),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2614),
.Y(n_2962)
);

BUFx3_ASAP7_75t_L g2963 ( 
.A(n_2756),
.Y(n_2963)
);

BUFx8_ASAP7_75t_SL g2964 ( 
.A(n_2650),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2642),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2645),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2681),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2682),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2683),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2688),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2706),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2706),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2622),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2775),
.B(n_2425),
.Y(n_2974)
);

INVx4_ASAP7_75t_R g2975 ( 
.A(n_2701),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2791),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2628),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2819),
.Y(n_2978)
);

OR2x2_ASAP7_75t_L g2979 ( 
.A(n_2820),
.B(n_2425),
.Y(n_2979)
);

HB1xp67_ASAP7_75t_L g2980 ( 
.A(n_2687),
.Y(n_2980)
);

AND2x2_ASAP7_75t_L g2981 ( 
.A(n_2793),
.B(n_2427),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2596),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2597),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2735),
.B(n_2558),
.Y(n_2984)
);

AND2x4_ASAP7_75t_L g2985 ( 
.A(n_2601),
.B(n_2441),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2598),
.Y(n_2986)
);

AND2x4_ASAP7_75t_L g2987 ( 
.A(n_2601),
.B(n_2445),
.Y(n_2987)
);

HB1xp67_ASAP7_75t_L g2988 ( 
.A(n_2687),
.Y(n_2988)
);

BUFx2_ASAP7_75t_SL g2989 ( 
.A(n_2613),
.Y(n_2989)
);

HB1xp67_ASAP7_75t_L g2990 ( 
.A(n_2719),
.Y(n_2990)
);

BUFx3_ASAP7_75t_L g2991 ( 
.A(n_2756),
.Y(n_2991)
);

AOI22xp33_ASAP7_75t_L g2992 ( 
.A1(n_2767),
.A2(n_2549),
.B1(n_2556),
.B2(n_2544),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2599),
.Y(n_2993)
);

OAI21xp33_ASAP7_75t_L g2994 ( 
.A1(n_2588),
.A2(n_2510),
.B(n_2256),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2793),
.B(n_2624),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2600),
.Y(n_2996)
);

NAND2x1_ASAP7_75t_L g2997 ( 
.A(n_2802),
.B(n_2539),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2605),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2674),
.B(n_2427),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2699),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2632),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2796),
.Y(n_3002)
);

BUFx2_ASAP7_75t_L g3003 ( 
.A(n_2631),
.Y(n_3003)
);

AND2x2_ASAP7_75t_L g3004 ( 
.A(n_2685),
.B(n_2427),
.Y(n_3004)
);

BUFx12f_ASAP7_75t_L g3005 ( 
.A(n_2786),
.Y(n_3005)
);

BUFx2_ASAP7_75t_L g3006 ( 
.A(n_2647),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2692),
.B(n_2427),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2647),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2710),
.B(n_2367),
.Y(n_3009)
);

INVx3_ASAP7_75t_L g3010 ( 
.A(n_2658),
.Y(n_3010)
);

BUFx2_ASAP7_75t_L g3011 ( 
.A(n_2658),
.Y(n_3011)
);

OR2x2_ASAP7_75t_L g3012 ( 
.A(n_2799),
.B(n_2411),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2634),
.Y(n_3013)
);

INVx2_ASAP7_75t_SL g3014 ( 
.A(n_2716),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_L g3015 ( 
.A1(n_2767),
.A2(n_2556),
.B1(n_2549),
.B2(n_2544),
.Y(n_3015)
);

BUFx3_ASAP7_75t_L g3016 ( 
.A(n_2768),
.Y(n_3016)
);

AND2x4_ASAP7_75t_L g3017 ( 
.A(n_2676),
.B(n_2445),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_2713),
.B(n_2367),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2636),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2640),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2676),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2615),
.Y(n_3022)
);

AND2x4_ASAP7_75t_L g3023 ( 
.A(n_2828),
.B(n_2448),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2609),
.B(n_2407),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2610),
.B(n_2407),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2616),
.Y(n_3026)
);

AND2x2_ASAP7_75t_L g3027 ( 
.A(n_2690),
.B(n_2412),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2745),
.B(n_2412),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_L g3029 ( 
.A1(n_2808),
.A2(n_2275),
.B1(n_2291),
.B2(n_2239),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2745),
.B(n_2431),
.Y(n_3030)
);

BUFx2_ASAP7_75t_L g3031 ( 
.A(n_2646),
.Y(n_3031)
);

AND2x4_ASAP7_75t_L g3032 ( 
.A(n_2828),
.B(n_2448),
.Y(n_3032)
);

HB1xp67_ASAP7_75t_L g3033 ( 
.A(n_2728),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2679),
.Y(n_3034)
);

INVx3_ASAP7_75t_L g3035 ( 
.A(n_2684),
.Y(n_3035)
);

BUFx2_ASAP7_75t_L g3036 ( 
.A(n_2646),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2675),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2679),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2591),
.B(n_2431),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2686),
.Y(n_3040)
);

AND2x2_ASAP7_75t_L g3041 ( 
.A(n_2834),
.B(n_2452),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2715),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2652),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2653),
.Y(n_3044)
);

HB1xp67_ASAP7_75t_L g3045 ( 
.A(n_2728),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2715),
.Y(n_3046)
);

OR2x2_ASAP7_75t_L g3047 ( 
.A(n_2772),
.B(n_2452),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2712),
.Y(n_3048)
);

HB1xp67_ASAP7_75t_L g3049 ( 
.A(n_2731),
.Y(n_3049)
);

HB1xp67_ASAP7_75t_L g3050 ( 
.A(n_2731),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2838),
.B(n_2481),
.Y(n_3051)
);

BUFx2_ASAP7_75t_L g3052 ( 
.A(n_2801),
.Y(n_3052)
);

INVx3_ASAP7_75t_L g3053 ( 
.A(n_2684),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2643),
.B(n_2486),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2670),
.B(n_2486),
.Y(n_3055)
);

AND2x4_ASAP7_75t_L g3056 ( 
.A(n_2802),
.B(n_2778),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2721),
.Y(n_3057)
);

CKINVDCx5p33_ASAP7_75t_R g3058 ( 
.A(n_2590),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2721),
.Y(n_3059)
);

INVx2_ASAP7_75t_SL g3060 ( 
.A(n_2716),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2655),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2630),
.B(n_2486),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2816),
.B(n_2560),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2661),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_2772),
.B(n_2240),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2585),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_2832),
.B(n_2306),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_2844),
.B(n_2306),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2750),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2587),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2844),
.B(n_2487),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2592),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2595),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2704),
.B(n_2487),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_2718),
.B(n_2498),
.Y(n_3075)
);

HB1xp67_ASAP7_75t_L g3076 ( 
.A(n_2747),
.Y(n_3076)
);

BUFx3_ASAP7_75t_L g3077 ( 
.A(n_2768),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2750),
.Y(n_3078)
);

AND2x2_ASAP7_75t_L g3079 ( 
.A(n_2588),
.B(n_2498),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2607),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2608),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_2800),
.B(n_2499),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2668),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2669),
.Y(n_3084)
);

AOI22xp33_ASAP7_75t_SL g3085 ( 
.A1(n_2817),
.A2(n_2275),
.B1(n_2291),
.B2(n_2323),
.Y(n_3085)
);

INVxp67_ASAP7_75t_L g3086 ( 
.A(n_2660),
.Y(n_3086)
);

AND2x2_ASAP7_75t_L g3087 ( 
.A(n_2800),
.B(n_2499),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2584),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2800),
.B(n_2391),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2663),
.Y(n_3090)
);

AND2x4_ASAP7_75t_L g3091 ( 
.A(n_2802),
.B(n_2560),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2664),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2729),
.Y(n_3093)
);

INVx2_ASAP7_75t_SL g3094 ( 
.A(n_2727),
.Y(n_3094)
);

BUFx5_ASAP7_75t_L g3095 ( 
.A(n_2665),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2667),
.Y(n_3096)
);

BUFx2_ASAP7_75t_L g3097 ( 
.A(n_2776),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2693),
.Y(n_3098)
);

INVx2_ASAP7_75t_SL g3099 ( 
.A(n_2727),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2693),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2737),
.B(n_2391),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2739),
.B(n_2341),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2773),
.Y(n_3103)
);

AOI22xp33_ASAP7_75t_L g3104 ( 
.A1(n_2808),
.A2(n_2323),
.B1(n_2550),
.B2(n_2555),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2773),
.Y(n_3105)
);

AND2x4_ASAP7_75t_L g3106 ( 
.A(n_2778),
.B(n_2552),
.Y(n_3106)
);

HB1xp67_ASAP7_75t_L g3107 ( 
.A(n_2620),
.Y(n_3107)
);

OR2x2_ASAP7_75t_L g3108 ( 
.A(n_2654),
.B(n_2318),
.Y(n_3108)
);

HB1xp67_ASAP7_75t_L g3109 ( 
.A(n_2812),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2788),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2788),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2659),
.Y(n_3112)
);

BUFx2_ASAP7_75t_L g3113 ( 
.A(n_2776),
.Y(n_3113)
);

CKINVDCx6p67_ASAP7_75t_R g3114 ( 
.A(n_2786),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2659),
.Y(n_3115)
);

OAI221xp5_ASAP7_75t_L g3116 ( 
.A1(n_2593),
.A2(n_2555),
.B1(n_2524),
.B2(n_2521),
.C(n_2550),
.Y(n_3116)
);

A2O1A1Ixp33_ASAP7_75t_L g3117 ( 
.A1(n_2817),
.A2(n_2351),
.B(n_2326),
.C(n_2557),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2804),
.B(n_2359),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_2736),
.Y(n_3119)
);

BUFx2_ASAP7_75t_L g3120 ( 
.A(n_2781),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2845),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_2856),
.B(n_2804),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2867),
.B(n_2782),
.Y(n_3123)
);

OAI22xp5_ASAP7_75t_L g3124 ( 
.A1(n_2891),
.A2(n_2886),
.B1(n_2950),
.B2(n_2770),
.Y(n_3124)
);

OR2x2_ASAP7_75t_L g3125 ( 
.A(n_2980),
.B(n_2806),
.Y(n_3125)
);

AND2x4_ASAP7_75t_L g3126 ( 
.A(n_2889),
.B(n_2781),
.Y(n_3126)
);

BUFx2_ASAP7_75t_L g3127 ( 
.A(n_3097),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_3054),
.B(n_2782),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_2871),
.B(n_2794),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_3062),
.B(n_2794),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2853),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2860),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2907),
.B(n_2797),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2847),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2849),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2923),
.B(n_2770),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2851),
.Y(n_3137)
);

AOI22xp33_ASAP7_75t_L g3138 ( 
.A1(n_2891),
.A2(n_2589),
.B1(n_2604),
.B2(n_2648),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_2908),
.B(n_2797),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2864),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2928),
.B(n_2825),
.Y(n_3141)
);

AND2x2_ASAP7_75t_L g3142 ( 
.A(n_2848),
.B(n_2825),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_2875),
.B(n_2806),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2859),
.Y(n_3144)
);

BUFx8_ASAP7_75t_SL g3145 ( 
.A(n_3005),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2869),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2865),
.Y(n_3147)
);

OR2x2_ASAP7_75t_L g3148 ( 
.A(n_2980),
.B(n_2810),
.Y(n_3148)
);

AND2x4_ASAP7_75t_L g3149 ( 
.A(n_2889),
.B(n_2810),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2873),
.B(n_2815),
.Y(n_3150)
);

OR2x2_ASAP7_75t_L g3151 ( 
.A(n_2988),
.B(n_2815),
.Y(n_3151)
);

HB1xp67_ASAP7_75t_L g3152 ( 
.A(n_2988),
.Y(n_3152)
);

AND2x4_ASAP7_75t_L g3153 ( 
.A(n_3056),
.B(n_2774),
.Y(n_3153)
);

AND2x4_ASAP7_75t_L g3154 ( 
.A(n_3056),
.B(n_2774),
.Y(n_3154)
);

AND2x2_ASAP7_75t_L g3155 ( 
.A(n_2930),
.B(n_2777),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2872),
.Y(n_3156)
);

AND2x4_ASAP7_75t_L g3157 ( 
.A(n_2903),
.B(n_2777),
.Y(n_3157)
);

OAI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_2886),
.A2(n_2593),
.B1(n_2573),
.B2(n_2589),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_SL g3159 ( 
.A(n_3003),
.B(n_2809),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_2912),
.B(n_2870),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2884),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2893),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2910),
.B(n_2784),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_3113),
.B(n_2784),
.Y(n_3164)
);

INVxp67_ASAP7_75t_L g3165 ( 
.A(n_2854),
.Y(n_3165)
);

AOI22xp33_ASAP7_75t_L g3166 ( 
.A1(n_2896),
.A2(n_2604),
.B1(n_2648),
.B2(n_2649),
.Y(n_3166)
);

AOI22xp33_ASAP7_75t_L g3167 ( 
.A1(n_2950),
.A2(n_2649),
.B1(n_2618),
.B2(n_2573),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2898),
.Y(n_3168)
);

OR2x2_ASAP7_75t_L g3169 ( 
.A(n_2938),
.B(n_2696),
.Y(n_3169)
);

BUFx2_ASAP7_75t_L g3170 ( 
.A(n_3120),
.Y(n_3170)
);

NAND2x1_ASAP7_75t_L g3171 ( 
.A(n_2857),
.B(n_2727),
.Y(n_3171)
);

HB1xp67_ASAP7_75t_L g3172 ( 
.A(n_2854),
.Y(n_3172)
);

AND2x2_ASAP7_75t_L g3173 ( 
.A(n_2883),
.B(n_2787),
.Y(n_3173)
);

AND2x4_ASAP7_75t_L g3174 ( 
.A(n_2903),
.B(n_2606),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2904),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_3024),
.B(n_2779),
.Y(n_3176)
);

INVxp67_ASAP7_75t_L g3177 ( 
.A(n_2862),
.Y(n_3177)
);

AOI22xp33_ASAP7_75t_SL g3178 ( 
.A1(n_3116),
.A2(n_2845),
.B1(n_2818),
.B2(n_2830),
.Y(n_3178)
);

INVx3_ASAP7_75t_L g3179 ( 
.A(n_2857),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2931),
.B(n_2787),
.Y(n_3180)
);

INVx3_ASAP7_75t_L g3181 ( 
.A(n_3010),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_3025),
.B(n_2783),
.Y(n_3182)
);

AND2x2_ASAP7_75t_SL g3183 ( 
.A(n_2846),
.B(n_2613),
.Y(n_3183)
);

AND2x2_ASAP7_75t_L g3184 ( 
.A(n_2934),
.B(n_2769),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2911),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_2978),
.B(n_2879),
.Y(n_3186)
);

INVxp67_ASAP7_75t_SL g3187 ( 
.A(n_3107),
.Y(n_3187)
);

AND2x2_ASAP7_75t_L g3188 ( 
.A(n_2915),
.B(n_2769),
.Y(n_3188)
);

AO22x1_ASAP7_75t_L g3189 ( 
.A1(n_2947),
.A2(n_2830),
.B1(n_2798),
.B2(n_2673),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2918),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_2995),
.B(n_2769),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2941),
.B(n_2814),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2965),
.B(n_2691),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_2966),
.B(n_3079),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2921),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2932),
.Y(n_3196)
);

BUFx2_ASAP7_75t_L g3197 ( 
.A(n_3006),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2936),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2946),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2917),
.Y(n_3200)
);

AOI22xp33_ASAP7_75t_L g3201 ( 
.A1(n_2960),
.A2(n_2618),
.B1(n_2637),
.B2(n_2550),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_3039),
.B(n_2691),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_3055),
.B(n_2826),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2933),
.Y(n_3204)
);

AND2x2_ASAP7_75t_L g3205 ( 
.A(n_3011),
.B(n_2826),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3066),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_2868),
.B(n_2823),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_3043),
.B(n_2621),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3070),
.Y(n_3209)
);

BUFx2_ASAP7_75t_L g3210 ( 
.A(n_2947),
.Y(n_3210)
);

AND2x4_ASAP7_75t_L g3211 ( 
.A(n_2913),
.B(n_2606),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3072),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3073),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2967),
.Y(n_3214)
);

OR2x2_ASAP7_75t_L g3215 ( 
.A(n_2906),
.B(n_2638),
.Y(n_3215)
);

HB1xp67_ASAP7_75t_L g3216 ( 
.A(n_2906),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2942),
.B(n_2638),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_3044),
.B(n_2621),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2968),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2969),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2901),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_2970),
.Y(n_3222)
);

INVx2_ASAP7_75t_L g3223 ( 
.A(n_2916),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_2888),
.B(n_2803),
.Y(n_3224)
);

HB1xp67_ASAP7_75t_L g3225 ( 
.A(n_2924),
.Y(n_3225)
);

BUFx2_ASAP7_75t_L g3226 ( 
.A(n_2852),
.Y(n_3226)
);

NOR2x1_ASAP7_75t_SL g3227 ( 
.A(n_2887),
.B(n_2702),
.Y(n_3227)
);

BUFx2_ASAP7_75t_L g3228 ( 
.A(n_2863),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3088),
.Y(n_3229)
);

AND2x4_ASAP7_75t_L g3230 ( 
.A(n_2913),
.B(n_2606),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3080),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3081),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2976),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2943),
.B(n_2602),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_2888),
.B(n_2803),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3002),
.Y(n_3236)
);

BUFx2_ASAP7_75t_L g3237 ( 
.A(n_2878),
.Y(n_3237)
);

BUFx3_ASAP7_75t_L g3238 ( 
.A(n_2878),
.Y(n_3238)
);

BUFx3_ASAP7_75t_L g3239 ( 
.A(n_2964),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_2905),
.B(n_2805),
.Y(n_3240)
);

CKINVDCx6p67_ASAP7_75t_R g3241 ( 
.A(n_2989),
.Y(n_3241)
);

AND2x4_ASAP7_75t_L g3242 ( 
.A(n_3106),
.B(n_2842),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2971),
.Y(n_3243)
);

NOR2xp67_ASAP7_75t_L g3244 ( 
.A(n_3107),
.B(n_2700),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_3009),
.B(n_2602),
.Y(n_3245)
);

CKINVDCx20_ASAP7_75t_R g3246 ( 
.A(n_2964),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3018),
.B(n_2765),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_2958),
.B(n_2765),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_2905),
.B(n_2805),
.Y(n_3249)
);

INVxp67_ASAP7_75t_SL g3250 ( 
.A(n_2925),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2959),
.B(n_2807),
.Y(n_3251)
);

AND2x4_ASAP7_75t_L g3252 ( 
.A(n_3106),
.B(n_2743),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_2972),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2951),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2956),
.Y(n_3255)
);

INVx4_ASAP7_75t_L g3256 ( 
.A(n_2948),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2961),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_3090),
.B(n_2709),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2962),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3092),
.B(n_2709),
.Y(n_3260)
);

AND2x2_ASAP7_75t_L g3261 ( 
.A(n_3001),
.B(n_2839),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2973),
.Y(n_3262)
);

BUFx2_ASAP7_75t_L g3263 ( 
.A(n_2914),
.Y(n_3263)
);

NOR2xp33_ASAP7_75t_L g3264 ( 
.A(n_3058),
.B(n_2590),
.Y(n_3264)
);

INVxp67_ASAP7_75t_SL g3265 ( 
.A(n_2925),
.Y(n_3265)
);

AND2x4_ASAP7_75t_L g3266 ( 
.A(n_3086),
.B(n_2746),
.Y(n_3266)
);

AOI22xp33_ASAP7_75t_L g3267 ( 
.A1(n_2960),
.A2(n_2637),
.B1(n_2561),
.B2(n_2680),
.Y(n_3267)
);

BUFx2_ASAP7_75t_L g3268 ( 
.A(n_2914),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_3013),
.B(n_2680),
.Y(n_3269)
);

INVxp67_ASAP7_75t_SL g3270 ( 
.A(n_2929),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_2858),
.A2(n_2792),
.B1(n_2524),
.B2(n_2351),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2977),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2982),
.Y(n_3273)
);

NOR2x1_ASAP7_75t_L g3274 ( 
.A(n_3010),
.B(n_2997),
.Y(n_3274)
);

INVxp67_ASAP7_75t_SL g3275 ( 
.A(n_2940),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_3019),
.B(n_2341),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_3061),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3020),
.B(n_2359),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3064),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2983),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2986),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_3086),
.B(n_2579),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2993),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3096),
.B(n_2579),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_2996),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2998),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3083),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3084),
.Y(n_3288)
);

AND2x4_ASAP7_75t_L g3289 ( 
.A(n_3091),
.B(n_2746),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_3101),
.B(n_2730),
.Y(n_3290)
);

HB1xp67_ASAP7_75t_L g3291 ( 
.A(n_2940),
.Y(n_3291)
);

INVx3_ASAP7_75t_L g3292 ( 
.A(n_2855),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3022),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3026),
.Y(n_3294)
);

INVxp67_ASAP7_75t_L g3295 ( 
.A(n_2953),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2953),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_2885),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2990),
.Y(n_3298)
);

OAI22xp5_ASAP7_75t_L g3299 ( 
.A1(n_3116),
.A2(n_2841),
.B1(n_2833),
.B2(n_2471),
.Y(n_3299)
);

AOI22xp33_ASAP7_75t_L g3300 ( 
.A1(n_2899),
.A2(n_2561),
.B1(n_2571),
.B2(n_2236),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3102),
.B(n_2736),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3000),
.B(n_2700),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_2885),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2990),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_2902),
.B(n_2757),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_2850),
.B(n_2763),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3033),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_2948),
.B(n_2798),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_2874),
.B(n_2714),
.Y(n_3309)
);

OAI222xp33_ASAP7_75t_L g3310 ( 
.A1(n_2927),
.A2(n_2744),
.B1(n_2841),
.B2(n_2833),
.C1(n_2619),
.C2(n_2711),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3180),
.B(n_3037),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3160),
.B(n_3040),
.Y(n_3312)
);

AND2x4_ASAP7_75t_L g3313 ( 
.A(n_3179),
.B(n_3112),
.Y(n_3313)
);

AND2x2_ASAP7_75t_L g3314 ( 
.A(n_3186),
.B(n_3048),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3134),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3135),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3137),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3144),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_3184),
.B(n_2981),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3146),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3150),
.B(n_3108),
.Y(n_3321)
);

OR2x6_ASAP7_75t_L g3322 ( 
.A(n_3274),
.B(n_2855),
.Y(n_3322)
);

AND2x2_ASAP7_75t_L g3323 ( 
.A(n_3202),
.B(n_3115),
.Y(n_3323)
);

OA211x2_ASAP7_75t_L g3324 ( 
.A1(n_3171),
.A2(n_3104),
.B(n_2994),
.C(n_3029),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3156),
.Y(n_3325)
);

OR2x2_ASAP7_75t_L g3326 ( 
.A(n_3152),
.B(n_3248),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3161),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3162),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3290),
.B(n_3194),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3123),
.B(n_2979),
.Y(n_3330)
);

NAND3xp33_ASAP7_75t_L g3331 ( 
.A(n_3158),
.B(n_3015),
.C(n_2992),
.Y(n_3331)
);

OR2x2_ASAP7_75t_L g3332 ( 
.A(n_3248),
.B(n_3251),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3282),
.B(n_3098),
.Y(n_3333)
);

AND2x2_ASAP7_75t_L g3334 ( 
.A(n_3128),
.B(n_3100),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3168),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_3258),
.B(n_2999),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_L g3337 ( 
.A(n_3158),
.B(n_3124),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3269),
.B(n_3207),
.Y(n_3338)
);

INVx3_ASAP7_75t_L g3339 ( 
.A(n_3181),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3166),
.B(n_2974),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_3260),
.B(n_3004),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3175),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3127),
.B(n_3033),
.Y(n_3343)
);

INVx2_ASAP7_75t_SL g3344 ( 
.A(n_3263),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3170),
.B(n_3045),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3301),
.B(n_3045),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3185),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3142),
.B(n_3007),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3190),
.Y(n_3349)
);

AND2x4_ASAP7_75t_SL g3350 ( 
.A(n_3241),
.B(n_2861),
.Y(n_3350)
);

OR2x2_ASAP7_75t_L g3351 ( 
.A(n_3251),
.B(n_3049),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3195),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_3203),
.B(n_3103),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3196),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_3129),
.B(n_3105),
.Y(n_3355)
);

HB1xp67_ASAP7_75t_L g3356 ( 
.A(n_3172),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3198),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3197),
.B(n_3110),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_3173),
.B(n_3111),
.Y(n_3359)
);

INVxp67_ASAP7_75t_SL g3360 ( 
.A(n_3187),
.Y(n_3360)
);

OR2x2_ASAP7_75t_L g3361 ( 
.A(n_3291),
.B(n_3049),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3169),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3163),
.B(n_3027),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3309),
.B(n_3041),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_3133),
.B(n_3050),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3208),
.B(n_3093),
.Y(n_3366)
);

NOR2xp67_ASAP7_75t_L g3367 ( 
.A(n_3238),
.B(n_2880),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3199),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_3139),
.B(n_3050),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_3131),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3132),
.Y(n_3371)
);

INVxp67_ASAP7_75t_L g3372 ( 
.A(n_3187),
.Y(n_3372)
);

INVx1_ASAP7_75t_SL g3373 ( 
.A(n_3210),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3214),
.Y(n_3374)
);

OR2x2_ASAP7_75t_L g3375 ( 
.A(n_3125),
.B(n_3076),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_3140),
.Y(n_3376)
);

OR2x2_ASAP7_75t_L g3377 ( 
.A(n_3148),
.B(n_3076),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3218),
.B(n_3028),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3147),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3219),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3193),
.B(n_3030),
.Y(n_3381)
);

HB1xp67_ASAP7_75t_L g3382 ( 
.A(n_3172),
.Y(n_3382)
);

NAND2x1_ASAP7_75t_SL g3383 ( 
.A(n_3274),
.B(n_2861),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3220),
.Y(n_3384)
);

NOR2x1_ASAP7_75t_L g3385 ( 
.A(n_3239),
.B(n_2949),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_3179),
.B(n_3109),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3222),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3284),
.B(n_3305),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_3306),
.B(n_3118),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_SL g3390 ( 
.A(n_3178),
.B(n_2927),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3206),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3209),
.Y(n_3392)
);

AND2x2_ASAP7_75t_L g3393 ( 
.A(n_3122),
.B(n_3071),
.Y(n_3393)
);

INVxp67_ASAP7_75t_L g3394 ( 
.A(n_3216),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3212),
.Y(n_3395)
);

HB1xp67_ASAP7_75t_L g3396 ( 
.A(n_3216),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3143),
.B(n_3089),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3155),
.B(n_3023),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3213),
.Y(n_3399)
);

OR2x2_ASAP7_75t_L g3400 ( 
.A(n_3151),
.B(n_3012),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3141),
.B(n_3023),
.Y(n_3401)
);

OR2x2_ASAP7_75t_L g3402 ( 
.A(n_3298),
.B(n_3063),
.Y(n_3402)
);

OR2x2_ASAP7_75t_L g3403 ( 
.A(n_3332),
.B(n_3247),
.Y(n_3403)
);

AND2x2_ASAP7_75t_L g3404 ( 
.A(n_3329),
.B(n_3153),
.Y(n_3404)
);

OR2x2_ASAP7_75t_L g3405 ( 
.A(n_3326),
.B(n_3247),
.Y(n_3405)
);

INVx1_ASAP7_75t_SL g3406 ( 
.A(n_3373),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3372),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_3329),
.B(n_3153),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_3372),
.Y(n_3409)
);

OR2x2_ASAP7_75t_L g3410 ( 
.A(n_3338),
.B(n_3225),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3388),
.B(n_3154),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3365),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3315),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3316),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3317),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3318),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3320),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3369),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3325),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_3327),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3328),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3335),
.Y(n_3422)
);

HB1xp67_ASAP7_75t_L g3423 ( 
.A(n_3360),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3370),
.Y(n_3424)
);

OR2x2_ASAP7_75t_L g3425 ( 
.A(n_3351),
.B(n_3225),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3342),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3333),
.B(n_3234),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3347),
.Y(n_3428)
);

OR2x2_ASAP7_75t_L g3429 ( 
.A(n_3388),
.B(n_3250),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3333),
.B(n_3234),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3349),
.Y(n_3431)
);

INVxp67_ASAP7_75t_SL g3432 ( 
.A(n_3360),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_3350),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_3381),
.B(n_3245),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3381),
.B(n_3245),
.Y(n_3435)
);

NOR2xp67_ASAP7_75t_R g3436 ( 
.A(n_3339),
.B(n_3268),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3370),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3352),
.Y(n_3438)
);

OR2x2_ASAP7_75t_L g3439 ( 
.A(n_3330),
.B(n_3250),
.Y(n_3439)
);

INVx2_ASAP7_75t_SL g3440 ( 
.A(n_3350),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3354),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3357),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3321),
.B(n_3154),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3378),
.B(n_3217),
.Y(n_3444)
);

INVx2_ASAP7_75t_SL g3445 ( 
.A(n_3401),
.Y(n_3445)
);

OR2x2_ASAP7_75t_L g3446 ( 
.A(n_3400),
.B(n_3265),
.Y(n_3446)
);

AND2x2_ASAP7_75t_L g3447 ( 
.A(n_3363),
.B(n_3205),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3368),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3371),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3374),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3378),
.B(n_3217),
.Y(n_3451)
);

INVx2_ASAP7_75t_L g3452 ( 
.A(n_3371),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3380),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3384),
.Y(n_3454)
);

OR2x2_ASAP7_75t_L g3455 ( 
.A(n_3311),
.B(n_3265),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3364),
.B(n_3130),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3387),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3391),
.Y(n_3458)
);

NAND2xp67_ASAP7_75t_L g3459 ( 
.A(n_3343),
.B(n_2954),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3392),
.Y(n_3460)
);

OR2x2_ASAP7_75t_L g3461 ( 
.A(n_3311),
.B(n_3270),
.Y(n_3461)
);

OR2x6_ASAP7_75t_L g3462 ( 
.A(n_3322),
.B(n_3174),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3395),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3399),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3376),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3398),
.B(n_3188),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3361),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3397),
.B(n_3224),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_L g3469 ( 
.A(n_3385),
.B(n_3237),
.Y(n_3469)
);

NAND2x1p5_ASAP7_75t_L g3470 ( 
.A(n_3367),
.B(n_3183),
.Y(n_3470)
);

OR2x2_ASAP7_75t_L g3471 ( 
.A(n_3334),
.B(n_3270),
.Y(n_3471)
);

OR2x2_ASAP7_75t_L g3472 ( 
.A(n_3334),
.B(n_3275),
.Y(n_3472)
);

OR2x2_ASAP7_75t_L g3473 ( 
.A(n_3402),
.B(n_3275),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3376),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3356),
.Y(n_3475)
);

NOR2xp33_ASAP7_75t_L g3476 ( 
.A(n_3337),
.B(n_3246),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3379),
.Y(n_3477)
);

INVxp67_ASAP7_75t_SL g3478 ( 
.A(n_3356),
.Y(n_3478)
);

HB1xp67_ASAP7_75t_L g3479 ( 
.A(n_3382),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3425),
.Y(n_3480)
);

OR2x2_ASAP7_75t_L g3481 ( 
.A(n_3444),
.B(n_3389),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3411),
.B(n_3313),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3413),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3414),
.Y(n_3484)
);

HB1xp67_ASAP7_75t_L g3485 ( 
.A(n_3423),
.Y(n_3485)
);

OAI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3470),
.A2(n_3390),
.B(n_2920),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3415),
.Y(n_3487)
);

NAND4xp25_ASAP7_75t_L g3488 ( 
.A(n_3469),
.B(n_3337),
.C(n_3324),
.D(n_3167),
.Y(n_3488)
);

OR2x2_ASAP7_75t_L g3489 ( 
.A(n_3444),
.B(n_3389),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3416),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3417),
.Y(n_3491)
);

AOI22xp5_ASAP7_75t_L g3492 ( 
.A1(n_3476),
.A2(n_3390),
.B1(n_3124),
.B2(n_3178),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3427),
.B(n_3430),
.Y(n_3493)
);

AOI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_3436),
.A2(n_3310),
.B(n_3227),
.Y(n_3494)
);

OAI21xp33_ASAP7_75t_SL g3495 ( 
.A1(n_3462),
.A2(n_3344),
.B(n_3383),
.Y(n_3495)
);

OAI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3470),
.A2(n_2920),
.B(n_3310),
.Y(n_3496)
);

INVx2_ASAP7_75t_L g3497 ( 
.A(n_3423),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3419),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3420),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3421),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3422),
.Y(n_3501)
);

INVxp67_ASAP7_75t_SL g3502 ( 
.A(n_3432),
.Y(n_3502)
);

NOR4xp75_ASAP7_75t_L g3503 ( 
.A(n_3433),
.B(n_3308),
.C(n_3159),
.D(n_3014),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3429),
.Y(n_3504)
);

AND2x4_ASAP7_75t_L g3505 ( 
.A(n_3462),
.B(n_3313),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3426),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3479),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3428),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3431),
.Y(n_3509)
);

HB1xp67_ASAP7_75t_SL g3510 ( 
.A(n_3440),
.Y(n_3510)
);

NOR2xp33_ASAP7_75t_L g3511 ( 
.A(n_3433),
.B(n_3114),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3438),
.Y(n_3512)
);

INVx1_ASAP7_75t_SL g3513 ( 
.A(n_3406),
.Y(n_3513)
);

INVxp33_ASAP7_75t_SL g3514 ( 
.A(n_3406),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3441),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3442),
.Y(n_3516)
);

AND2x2_ASAP7_75t_L g3517 ( 
.A(n_3443),
.B(n_3313),
.Y(n_3517)
);

INVx1_ASAP7_75t_SL g3518 ( 
.A(n_3446),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3427),
.B(n_3323),
.Y(n_3519)
);

INVx1_ASAP7_75t_SL g3520 ( 
.A(n_3456),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3404),
.B(n_3312),
.Y(n_3521)
);

AOI22xp5_ASAP7_75t_L g3522 ( 
.A1(n_3467),
.A2(n_3138),
.B1(n_3331),
.B2(n_3323),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3424),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3448),
.Y(n_3524)
);

NAND2x1_ASAP7_75t_L g3525 ( 
.A(n_3462),
.B(n_3322),
.Y(n_3525)
);

OAI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3445),
.A2(n_3201),
.B1(n_3344),
.B2(n_3432),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_SL g3527 ( 
.A(n_3436),
.B(n_3478),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3450),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3408),
.B(n_3348),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3437),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3453),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_3468),
.B(n_3447),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3454),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3449),
.Y(n_3534)
);

AOI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_3478),
.A2(n_3136),
.B(n_3322),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3457),
.Y(n_3536)
);

NOR2xp33_ASAP7_75t_L g3537 ( 
.A(n_3405),
.B(n_3145),
.Y(n_3537)
);

AOI211x1_ASAP7_75t_SL g3538 ( 
.A1(n_3407),
.A2(n_3299),
.B(n_3244),
.C(n_3366),
.Y(n_3538)
);

OAI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_3475),
.A2(n_3228),
.B(n_3226),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3466),
.B(n_3319),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3458),
.Y(n_3541)
);

NAND4xp25_ASAP7_75t_L g3542 ( 
.A(n_3430),
.B(n_3267),
.C(n_2890),
.D(n_3264),
.Y(n_3542)
);

INVx1_ASAP7_75t_SL g3543 ( 
.A(n_3455),
.Y(n_3543)
);

HB1xp67_ASAP7_75t_L g3544 ( 
.A(n_3461),
.Y(n_3544)
);

OAI31xp33_ASAP7_75t_L g3545 ( 
.A1(n_3471),
.A2(n_3036),
.A3(n_3031),
.B(n_2955),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3460),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3434),
.B(n_3393),
.Y(n_3547)
);

INVxp67_ASAP7_75t_L g3548 ( 
.A(n_3510),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3544),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3494),
.A2(n_3189),
.B(n_3451),
.Y(n_3550)
);

OAI21xp33_ASAP7_75t_SL g3551 ( 
.A1(n_3527),
.A2(n_3472),
.B(n_3435),
.Y(n_3551)
);

OAI22xp5_ASAP7_75t_L g3552 ( 
.A1(n_3486),
.A2(n_3410),
.B1(n_3403),
.B2(n_3451),
.Y(n_3552)
);

NAND3xp33_ASAP7_75t_L g3553 ( 
.A(n_3492),
.B(n_2880),
.C(n_2919),
.Y(n_3553)
);

OAI21xp33_ASAP7_75t_L g3554 ( 
.A1(n_3488),
.A2(n_3459),
.B(n_3435),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3483),
.Y(n_3555)
);

OAI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3495),
.A2(n_3394),
.B(n_3271),
.Y(n_3556)
);

NAND2x1p5_ASAP7_75t_L g3557 ( 
.A(n_3513),
.B(n_2952),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3513),
.B(n_3434),
.Y(n_3558)
);

OAI221xp5_ASAP7_75t_L g3559 ( 
.A1(n_3488),
.A2(n_3439),
.B1(n_3473),
.B2(n_3104),
.C(n_3340),
.Y(n_3559)
);

AOI21xp33_ASAP7_75t_L g3560 ( 
.A1(n_3511),
.A2(n_3060),
.B(n_2926),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3484),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3487),
.Y(n_3562)
);

AOI31xp33_ASAP7_75t_L g3563 ( 
.A1(n_3496),
.A2(n_3537),
.A3(n_2919),
.B(n_2635),
.Y(n_3563)
);

AOI22xp5_ASAP7_75t_L g3564 ( 
.A1(n_3526),
.A2(n_3345),
.B1(n_3353),
.B2(n_3358),
.Y(n_3564)
);

AOI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_3542),
.A2(n_3174),
.B1(n_3230),
.B2(n_3211),
.Y(n_3565)
);

NOR2xp33_ASAP7_75t_L g3566 ( 
.A(n_3514),
.B(n_2586),
.Y(n_3566)
);

AOI22xp5_ASAP7_75t_L g3567 ( 
.A1(n_3522),
.A2(n_3314),
.B1(n_3346),
.B2(n_3359),
.Y(n_3567)
);

O2A1O1Ixp33_ASAP7_75t_L g3568 ( 
.A1(n_3502),
.A2(n_3099),
.B(n_3094),
.C(n_3052),
.Y(n_3568)
);

NOR2x1_ASAP7_75t_L g3569 ( 
.A(n_3525),
.B(n_2619),
.Y(n_3569)
);

OAI21xp5_ASAP7_75t_SL g3570 ( 
.A1(n_3538),
.A2(n_2909),
.B(n_2866),
.Y(n_3570)
);

OR2x2_ASAP7_75t_L g3571 ( 
.A(n_3493),
.B(n_3409),
.Y(n_3571)
);

OAI22xp5_ASAP7_75t_L g3572 ( 
.A1(n_3520),
.A2(n_3505),
.B1(n_3543),
.B2(n_3518),
.Y(n_3572)
);

A2O1A1Ixp33_ASAP7_75t_L g3573 ( 
.A1(n_3545),
.A2(n_2955),
.B(n_2952),
.C(n_3058),
.Y(n_3573)
);

AOI32xp33_ASAP7_75t_L g3574 ( 
.A1(n_3518),
.A2(n_3412),
.A3(n_3418),
.B1(n_3386),
.B2(n_3355),
.Y(n_3574)
);

INVxp67_ASAP7_75t_L g3575 ( 
.A(n_3485),
.Y(n_3575)
);

BUFx3_ASAP7_75t_L g3576 ( 
.A(n_3507),
.Y(n_3576)
);

OAI22xp5_ASAP7_75t_L g3577 ( 
.A1(n_3505),
.A2(n_3375),
.B1(n_3377),
.B2(n_3126),
.Y(n_3577)
);

OAI221xp5_ASAP7_75t_SL g3578 ( 
.A1(n_3545),
.A2(n_3300),
.B1(n_3271),
.B2(n_3121),
.C(n_2992),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3543),
.B(n_3382),
.Y(n_3579)
);

AOI21xp33_ASAP7_75t_SL g3580 ( 
.A1(n_3539),
.A2(n_2673),
.B(n_2711),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3480),
.B(n_3396),
.Y(n_3581)
);

A2O1A1Ixp33_ASAP7_75t_L g3582 ( 
.A1(n_3535),
.A2(n_2780),
.B(n_3126),
.C(n_3463),
.Y(n_3582)
);

OAI32xp33_ASAP7_75t_L g3583 ( 
.A1(n_3538),
.A2(n_3396),
.A3(n_3256),
.B1(n_3339),
.B2(n_3394),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3519),
.B(n_3464),
.Y(n_3584)
);

AOI22xp5_ASAP7_75t_L g3585 ( 
.A1(n_3542),
.A2(n_3504),
.B1(n_3491),
.B2(n_3498),
.Y(n_3585)
);

INVxp33_ASAP7_75t_L g3586 ( 
.A(n_3517),
.Y(n_3586)
);

AOI221xp5_ASAP7_75t_L g3587 ( 
.A1(n_3490),
.A2(n_3299),
.B1(n_3255),
.B2(n_3259),
.C(n_3257),
.Y(n_3587)
);

AOI22xp5_ASAP7_75t_L g3588 ( 
.A1(n_3499),
.A2(n_3341),
.B1(n_3336),
.B2(n_3386),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3500),
.Y(n_3589)
);

AOI22xp5_ASAP7_75t_L g3590 ( 
.A1(n_3501),
.A2(n_3341),
.B1(n_3336),
.B2(n_3386),
.Y(n_3590)
);

AOI22xp5_ASAP7_75t_L g3591 ( 
.A1(n_3506),
.A2(n_3164),
.B1(n_3051),
.B2(n_3211),
.Y(n_3591)
);

INVxp67_ASAP7_75t_SL g3592 ( 
.A(n_3497),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3571),
.Y(n_3593)
);

AOI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_3553),
.A2(n_3509),
.B1(n_3512),
.B2(n_3508),
.Y(n_3594)
);

A2O1A1Ixp33_ASAP7_75t_L g3595 ( 
.A1(n_3548),
.A2(n_3521),
.B(n_3489),
.C(n_3481),
.Y(n_3595)
);

AOI221xp5_ASAP7_75t_L g3596 ( 
.A1(n_3553),
.A2(n_3515),
.B1(n_3528),
.B2(n_3524),
.C(n_3516),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3569),
.A2(n_3533),
.B(n_3531),
.Y(n_3597)
);

AOI21xp33_ASAP7_75t_L g3598 ( 
.A1(n_3568),
.A2(n_2752),
.B(n_3536),
.Y(n_3598)
);

AOI211xp5_ASAP7_75t_L g3599 ( 
.A1(n_3578),
.A2(n_2752),
.B(n_3503),
.C(n_2376),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3549),
.Y(n_3600)
);

AOI221xp5_ASAP7_75t_L g3601 ( 
.A1(n_3554),
.A2(n_3546),
.B1(n_3541),
.B2(n_3547),
.C(n_3532),
.Y(n_3601)
);

OAI221xp5_ASAP7_75t_L g3602 ( 
.A1(n_3551),
.A2(n_3015),
.B1(n_3029),
.B2(n_3085),
.C(n_3523),
.Y(n_3602)
);

AOI221xp5_ASAP7_75t_L g3603 ( 
.A1(n_3559),
.A2(n_3534),
.B1(n_3530),
.B2(n_3229),
.C(n_3254),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3585),
.B(n_3540),
.Y(n_3604)
);

NAND4xp25_ASAP7_75t_SL g3605 ( 
.A(n_3550),
.B(n_3482),
.C(n_3529),
.D(n_2975),
.Y(n_3605)
);

AOI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_3563),
.A2(n_2758),
.B(n_3165),
.Y(n_3606)
);

AOI221xp5_ASAP7_75t_L g3607 ( 
.A1(n_3572),
.A2(n_3273),
.B1(n_3280),
.B2(n_3272),
.C(n_3262),
.Y(n_3607)
);

HB1xp67_ASAP7_75t_L g3608 ( 
.A(n_3575),
.Y(n_3608)
);

AOI32xp33_ASAP7_75t_L g3609 ( 
.A1(n_3565),
.A2(n_3256),
.A3(n_3339),
.B1(n_3149),
.B2(n_2963),
.Y(n_3609)
);

INVx2_ASAP7_75t_SL g3610 ( 
.A(n_3557),
.Y(n_3610)
);

NAND3xp33_ASAP7_75t_L g3611 ( 
.A(n_3556),
.B(n_2795),
.C(n_2790),
.Y(n_3611)
);

AOI32xp33_ASAP7_75t_L g3612 ( 
.A1(n_3552),
.A2(n_3149),
.A3(n_2963),
.B1(n_3077),
.B2(n_3016),
.Y(n_3612)
);

O2A1O1Ixp33_ASAP7_75t_L g3613 ( 
.A1(n_3583),
.A2(n_2689),
.B(n_3117),
.C(n_2957),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3581),
.Y(n_3614)
);

AOI222xp33_ASAP7_75t_L g3615 ( 
.A1(n_3570),
.A2(n_2795),
.B1(n_3281),
.B2(n_3286),
.C1(n_3287),
.C2(n_3288),
.Y(n_3615)
);

AOI221xp5_ASAP7_75t_L g3616 ( 
.A1(n_3580),
.A2(n_3294),
.B1(n_3293),
.B2(n_3283),
.C(n_3243),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_L g3617 ( 
.A(n_3587),
.B(n_3304),
.Y(n_3617)
);

OA22x2_ASAP7_75t_L g3618 ( 
.A1(n_3564),
.A2(n_3567),
.B1(n_3590),
.B2(n_3588),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3555),
.Y(n_3619)
);

XNOR2xp5_ASAP7_75t_L g3620 ( 
.A(n_3591),
.B(n_2581),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3558),
.B(n_3307),
.Y(n_3621)
);

AOI322xp5_ASAP7_75t_L g3622 ( 
.A1(n_3566),
.A2(n_2753),
.A3(n_3177),
.B1(n_3295),
.B2(n_3165),
.C1(n_3067),
.C2(n_3068),
.Y(n_3622)
);

AO22x1_ASAP7_75t_L g3623 ( 
.A1(n_3586),
.A2(n_2581),
.B1(n_3157),
.B2(n_2948),
.Y(n_3623)
);

NOR2xp33_ASAP7_75t_L g3624 ( 
.A(n_3584),
.B(n_2790),
.Y(n_3624)
);

OAI221xp5_ASAP7_75t_SL g3625 ( 
.A1(n_3574),
.A2(n_3065),
.B1(n_3047),
.B2(n_3191),
.C(n_3117),
.Y(n_3625)
);

BUFx2_ASAP7_75t_L g3626 ( 
.A(n_3576),
.Y(n_3626)
);

AOI21x1_ASAP7_75t_L g3627 ( 
.A1(n_3579),
.A2(n_3244),
.B(n_3021),
.Y(n_3627)
);

AOI211xp5_ASAP7_75t_L g3628 ( 
.A1(n_3573),
.A2(n_2957),
.B(n_3230),
.C(n_2689),
.Y(n_3628)
);

NAND3x1_ASAP7_75t_L g3629 ( 
.A(n_3561),
.B(n_2882),
.C(n_2876),
.Y(n_3629)
);

OAI21xp33_ASAP7_75t_L g3630 ( 
.A1(n_3582),
.A2(n_3577),
.B(n_3592),
.Y(n_3630)
);

OAI21xp33_ASAP7_75t_SL g3631 ( 
.A1(n_3589),
.A2(n_3295),
.B(n_3177),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3562),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3560),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_SL g3634 ( 
.A(n_3569),
.B(n_3452),
.Y(n_3634)
);

AOI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_3548),
.A2(n_3474),
.B(n_3465),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3571),
.Y(n_3636)
);

AOI222xp33_ASAP7_75t_L g3637 ( 
.A1(n_3548),
.A2(n_3253),
.B1(n_3200),
.B2(n_3204),
.C1(n_2945),
.C2(n_2944),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3585),
.B(n_3477),
.Y(n_3638)
);

AOI221xp5_ASAP7_75t_L g3639 ( 
.A1(n_3553),
.A2(n_3296),
.B1(n_3362),
.B2(n_3236),
.C(n_3233),
.Y(n_3639)
);

AOI221xp5_ASAP7_75t_L g3640 ( 
.A1(n_3553),
.A2(n_3362),
.B1(n_3232),
.B2(n_3266),
.C(n_3302),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3608),
.Y(n_3641)
);

AOI221xp5_ASAP7_75t_L g3642 ( 
.A1(n_3602),
.A2(n_3266),
.B1(n_3302),
.B2(n_3252),
.C(n_3279),
.Y(n_3642)
);

NAND4xp25_ASAP7_75t_L g3643 ( 
.A(n_3611),
.B(n_2877),
.C(n_2900),
.D(n_2881),
.Y(n_3643)
);

NOR4xp25_ASAP7_75t_L g3644 ( 
.A(n_3633),
.B(n_3074),
.C(n_3075),
.D(n_2764),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3637),
.B(n_3593),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3626),
.Y(n_3646)
);

NOR2xp33_ASAP7_75t_SL g3647 ( 
.A(n_3605),
.B(n_2629),
.Y(n_3647)
);

NOR2x1_ASAP7_75t_L g3648 ( 
.A(n_3634),
.B(n_2877),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_SL g3649 ( 
.A(n_3631),
.B(n_2617),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3636),
.Y(n_3650)
);

NAND3xp33_ASAP7_75t_SL g3651 ( 
.A(n_3599),
.B(n_2813),
.C(n_2629),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3600),
.Y(n_3652)
);

OAI21xp5_ASAP7_75t_L g3653 ( 
.A1(n_3618),
.A2(n_3085),
.B(n_2764),
.Y(n_3653)
);

INVx1_ASAP7_75t_SL g3654 ( 
.A(n_3606),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3603),
.B(n_3277),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3614),
.B(n_3285),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_SL g3657 ( 
.A(n_3630),
.B(n_2617),
.Y(n_3657)
);

NAND2xp33_ASAP7_75t_L g3658 ( 
.A(n_3612),
.B(n_3095),
.Y(n_3658)
);

NOR2x1_ASAP7_75t_L g3659 ( 
.A(n_3635),
.B(n_2881),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3607),
.B(n_3261),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3621),
.Y(n_3661)
);

A2O1A1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3609),
.A2(n_2900),
.B(n_3016),
.C(n_2991),
.Y(n_3662)
);

NAND3xp33_ASAP7_75t_L g3663 ( 
.A(n_3601),
.B(n_3008),
.C(n_2561),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_L g3664 ( 
.A(n_3624),
.B(n_3157),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_SL g3665 ( 
.A(n_3615),
.B(n_3181),
.Y(n_3665)
);

AOI21xp5_ASAP7_75t_L g3666 ( 
.A1(n_3623),
.A2(n_2984),
.B(n_2939),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3619),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_SL g3668 ( 
.A(n_3639),
.B(n_3379),
.Y(n_3668)
);

AOI221xp5_ASAP7_75t_L g3669 ( 
.A1(n_3625),
.A2(n_3252),
.B1(n_3182),
.B2(n_3176),
.C(n_3192),
.Y(n_3669)
);

OA22x2_ASAP7_75t_L g3670 ( 
.A1(n_3594),
.A2(n_3091),
.B1(n_3292),
.B2(n_3053),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3617),
.B(n_3596),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3595),
.B(n_3297),
.Y(n_3672)
);

NOR2x1p5_ASAP7_75t_SL g3673 ( 
.A(n_3646),
.B(n_3627),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3641),
.Y(n_3674)
);

OAI211xp5_ASAP7_75t_L g3675 ( 
.A1(n_3657),
.A2(n_3622),
.B(n_3598),
.C(n_3628),
.Y(n_3675)
);

NAND4xp25_ASAP7_75t_L g3676 ( 
.A(n_3651),
.B(n_3622),
.C(n_3613),
.D(n_3640),
.Y(n_3676)
);

NAND3xp33_ASAP7_75t_SL g3677 ( 
.A(n_3654),
.B(n_3597),
.C(n_3604),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3656),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3650),
.Y(n_3679)
);

XNOR2xp5_ASAP7_75t_L g3680 ( 
.A(n_3643),
.B(n_3620),
.Y(n_3680)
);

NAND2x1_ASAP7_75t_SL g3681 ( 
.A(n_3648),
.B(n_3659),
.Y(n_3681)
);

NAND2x1_ASAP7_75t_SL g3682 ( 
.A(n_3652),
.B(n_3632),
.Y(n_3682)
);

NOR2xp33_ASAP7_75t_L g3683 ( 
.A(n_3647),
.B(n_3610),
.Y(n_3683)
);

AO22x2_ASAP7_75t_L g3684 ( 
.A1(n_3671),
.A2(n_3638),
.B1(n_3629),
.B2(n_2876),
.Y(n_3684)
);

AOI22x1_ASAP7_75t_SL g3685 ( 
.A1(n_3667),
.A2(n_2897),
.B1(n_2895),
.B2(n_2882),
.Y(n_3685)
);

NOR2x1_ASAP7_75t_L g3686 ( 
.A(n_3649),
.B(n_2991),
.Y(n_3686)
);

NOR2xp67_ASAP7_75t_L g3687 ( 
.A(n_3663),
.B(n_3292),
.Y(n_3687)
);

AOI22xp5_ASAP7_75t_L g3688 ( 
.A1(n_3653),
.A2(n_3616),
.B1(n_3240),
.B2(n_3249),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_3645),
.B(n_3077),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3661),
.Y(n_3690)
);

INVx2_ASAP7_75t_SL g3691 ( 
.A(n_3664),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_L g3692 ( 
.A(n_3660),
.B(n_2895),
.Y(n_3692)
);

NOR2xp33_ASAP7_75t_L g3693 ( 
.A(n_3655),
.B(n_2897),
.Y(n_3693)
);

NOR2xp33_ASAP7_75t_L g3694 ( 
.A(n_3672),
.B(n_2892),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3644),
.B(n_3303),
.Y(n_3695)
);

NOR2x1_ASAP7_75t_L g3696 ( 
.A(n_3665),
.B(n_3035),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3668),
.B(n_2892),
.Y(n_3697)
);

NAND3xp33_ASAP7_75t_L g3698 ( 
.A(n_3642),
.B(n_2401),
.C(n_2522),
.Y(n_3698)
);

NAND3xp33_ASAP7_75t_L g3699 ( 
.A(n_3674),
.B(n_3669),
.C(n_3658),
.Y(n_3699)
);

NOR2x1p5_ASAP7_75t_L g3700 ( 
.A(n_3677),
.B(n_3670),
.Y(n_3700)
);

NOR2x1_ASAP7_75t_L g3701 ( 
.A(n_3675),
.B(n_3662),
.Y(n_3701)
);

NOR3xp33_ASAP7_75t_L g3702 ( 
.A(n_3676),
.B(n_3666),
.C(n_3670),
.Y(n_3702)
);

NAND2x1p5_ASAP7_75t_L g3703 ( 
.A(n_3686),
.B(n_3035),
.Y(n_3703)
);

NOR2x1_ASAP7_75t_L g3704 ( 
.A(n_3680),
.B(n_3053),
.Y(n_3704)
);

NOR4xp75_ASAP7_75t_L g3705 ( 
.A(n_3682),
.B(n_2894),
.C(n_3119),
.D(n_2281),
.Y(n_3705)
);

NOR2x1_ASAP7_75t_L g3706 ( 
.A(n_3696),
.B(n_3679),
.Y(n_3706)
);

NAND3xp33_ASAP7_75t_L g3707 ( 
.A(n_3689),
.B(n_2522),
.C(n_3082),
.Y(n_3707)
);

NAND2x1p5_ASAP7_75t_SL g3708 ( 
.A(n_3691),
.B(n_3087),
.Y(n_3708)
);

AOI22xp5_ASAP7_75t_L g3709 ( 
.A1(n_3683),
.A2(n_3693),
.B1(n_3692),
.B2(n_3694),
.Y(n_3709)
);

NAND3xp33_ASAP7_75t_L g3710 ( 
.A(n_3690),
.B(n_2522),
.C(n_2469),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3678),
.B(n_3221),
.Y(n_3711)
);

OA22x2_ASAP7_75t_SL g3712 ( 
.A1(n_3681),
.A2(n_3231),
.B1(n_3223),
.B2(n_3038),
.Y(n_3712)
);

AND3x1_ASAP7_75t_L g3713 ( 
.A(n_3697),
.B(n_2894),
.C(n_3119),
.Y(n_3713)
);

OAI22x1_ASAP7_75t_L g3714 ( 
.A1(n_3688),
.A2(n_2576),
.B1(n_3017),
.B2(n_2987),
.Y(n_3714)
);

NOR3xp33_ASAP7_75t_L g3715 ( 
.A(n_3695),
.B(n_2299),
.C(n_2348),
.Y(n_3715)
);

NAND4xp75_ASAP7_75t_L g3716 ( 
.A(n_3673),
.B(n_2347),
.C(n_2237),
.D(n_2935),
.Y(n_3716)
);

INVxp33_ASAP7_75t_L g3717 ( 
.A(n_3698),
.Y(n_3717)
);

NAND4xp75_ASAP7_75t_L g3718 ( 
.A(n_3687),
.B(n_2347),
.C(n_2237),
.D(n_2937),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3702),
.B(n_3684),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3711),
.Y(n_3720)
);

NOR2x1_ASAP7_75t_L g3721 ( 
.A(n_3701),
.B(n_3684),
.Y(n_3721)
);

NOR2x1_ASAP7_75t_L g3722 ( 
.A(n_3700),
.B(n_3685),
.Y(n_3722)
);

AOI22xp5_ASAP7_75t_L g3723 ( 
.A1(n_3717),
.A2(n_3235),
.B1(n_2922),
.B2(n_3095),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3704),
.B(n_3242),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3708),
.B(n_3276),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3706),
.Y(n_3726)
);

NOR2x1_ASAP7_75t_L g3727 ( 
.A(n_3699),
.B(n_2405),
.Y(n_3727)
);

NAND4xp75_ASAP7_75t_L g3728 ( 
.A(n_3713),
.B(n_2432),
.C(n_2405),
.D(n_2511),
.Y(n_3728)
);

NOR2xp33_ASAP7_75t_L g3729 ( 
.A(n_3709),
.B(n_2576),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3712),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3714),
.Y(n_3731)
);

INVxp33_ASAP7_75t_SL g3732 ( 
.A(n_3705),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3720),
.Y(n_3733)
);

AND3x4_ASAP7_75t_L g3734 ( 
.A(n_3722),
.B(n_3715),
.C(n_3707),
.Y(n_3734)
);

NAND3x1_ASAP7_75t_L g3735 ( 
.A(n_3721),
.B(n_3703),
.C(n_3710),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3731),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3719),
.B(n_3716),
.Y(n_3737)
);

BUFx2_ASAP7_75t_L g3738 ( 
.A(n_3730),
.Y(n_3738)
);

AOI22xp33_ASAP7_75t_L g3739 ( 
.A1(n_3732),
.A2(n_3718),
.B1(n_3242),
.B2(n_3278),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3726),
.Y(n_3740)
);

OR2x2_ASAP7_75t_L g3741 ( 
.A(n_3725),
.B(n_3215),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3729),
.B(n_3289),
.Y(n_3742)
);

INVx2_ASAP7_75t_SL g3743 ( 
.A(n_3724),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3723),
.B(n_3017),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3736),
.Y(n_3745)
);

NOR2xp33_ASAP7_75t_L g3746 ( 
.A(n_3738),
.B(n_3727),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3740),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_3743),
.B(n_3728),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3744),
.B(n_2985),
.Y(n_3749)
);

AO22x2_ASAP7_75t_L g3750 ( 
.A1(n_3733),
.A2(n_2987),
.B1(n_2985),
.B2(n_3034),
.Y(n_3750)
);

AOI22xp5_ASAP7_75t_L g3751 ( 
.A1(n_3734),
.A2(n_3095),
.B1(n_2922),
.B2(n_3057),
.Y(n_3751)
);

AOI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_3735),
.A2(n_3095),
.B1(n_3046),
.B2(n_3042),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3750),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3750),
.Y(n_3754)
);

AOI22xp5_ASAP7_75t_SL g3755 ( 
.A1(n_3748),
.A2(n_3737),
.B1(n_3733),
.B2(n_3742),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3753),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3755),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3754),
.Y(n_3758)
);

AOI22xp5_ASAP7_75t_L g3759 ( 
.A1(n_3757),
.A2(n_3746),
.B1(n_3745),
.B2(n_3747),
.Y(n_3759)
);

OAI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_3759),
.A2(n_3756),
.B1(n_3758),
.B2(n_3749),
.Y(n_3760)
);

AOI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_3760),
.A2(n_3741),
.B(n_3751),
.Y(n_3761)
);

AOI221xp5_ASAP7_75t_L g3762 ( 
.A1(n_3761),
.A2(n_3739),
.B1(n_3752),
.B2(n_3059),
.C(n_3069),
.Y(n_3762)
);

AOI22xp33_ASAP7_75t_L g3763 ( 
.A1(n_3762),
.A2(n_3095),
.B1(n_3078),
.B2(n_3032),
.Y(n_3763)
);


endmodule