module fake_jpeg_20484_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_4),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_8),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_8),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_48),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_28),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_30),
.B1(n_31),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_62),
.B1(n_23),
.B2(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_30),
.B1(n_31),
.B2(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_28),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_26),
.B(n_0),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_42),
.B1(n_30),
.B2(n_39),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_76),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_42),
.B1(n_30),
.B2(n_39),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_41),
.B1(n_39),
.B2(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_78),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_41),
.B1(n_33),
.B2(n_34),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_41),
.B1(n_34),
.B2(n_33),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_46),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_19),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_60),
.B1(n_58),
.B2(n_65),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_95),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_21),
.C(n_26),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_104),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_60),
.B1(n_58),
.B2(n_53),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_71),
.B1(n_68),
.B2(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g124 ( 
.A(n_97),
.Y(n_124)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_64),
.C(n_33),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_110),
.C(n_64),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_84),
.B1(n_78),
.B2(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_102),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_105),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_20),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_52),
.Y(n_105)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_73),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_17),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_113),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_72),
.B(n_87),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_95),
.B(n_22),
.Y(n_149)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_91),
.B1(n_109),
.B2(n_90),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_129),
.B1(n_134),
.B2(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_104),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_70),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_76),
.B1(n_80),
.B2(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_19),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_61),
.B1(n_57),
.B2(n_65),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_89),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_54),
.B1(n_63),
.B2(n_32),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_25),
.B1(n_63),
.B2(n_24),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_109),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_149),
.B(n_134),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_99),
.C(n_110),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_147),
.C(n_26),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g143 ( 
.A(n_124),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_132),
.B1(n_128),
.B2(n_117),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_26),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_92),
.C(n_98),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_115),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_153),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_118),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_133),
.B1(n_116),
.B2(n_123),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_16),
.Y(n_155)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_22),
.B(n_23),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_106),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_126),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_32),
.B1(n_31),
.B2(n_20),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_16),
.B(n_24),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_119),
.B(n_123),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_163),
.B(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_166),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_168),
.B1(n_169),
.B2(n_176),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_129),
.B1(n_113),
.B2(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_135),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_179),
.C(n_173),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_117),
.B1(n_16),
.B2(n_24),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_142),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_19),
.B1(n_26),
.B2(n_59),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_180),
.B1(n_144),
.B2(n_143),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_59),
.C(n_26),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_147),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_189),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_192),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_146),
.C(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_183),
.B(n_186),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_149),
.B(n_136),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_157),
.Y(n_189)
);

XNOR2x2_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_155),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_166),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_151),
.C(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_196),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_197),
.B1(n_164),
.B2(n_161),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_144),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_207),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_175),
.B(n_167),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_166),
.C(n_165),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_168),
.B1(n_180),
.B2(n_172),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_210),
.A2(n_211),
.B1(n_191),
.B2(n_197),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_178),
.B1(n_170),
.B2(n_164),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_184),
.B1(n_182),
.B2(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_189),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_181),
.C(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_222),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_140),
.C(n_165),
.Y(n_222)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_224),
.CI(n_201),
.CON(n_229),
.SN(n_229)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_206),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_152),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_210),
.B1(n_211),
.B2(n_3),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_215),
.A2(n_199),
.B(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_229),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_224),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_237),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_219),
.B(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_234),
.B(n_216),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_214),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_240),
.A2(n_233),
.B(n_229),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_240),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_218),
.A3(n_223),
.B1(n_221),
.B2(n_7),
.C1(n_10),
.C2(n_11),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_14),
.B1(n_5),
.B2(n_6),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g247 ( 
.A1(n_239),
.A2(n_5),
.A3(n_7),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_0),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_5),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_250),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_235),
.C(n_7),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_246),
.B(n_243),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_248),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_253),
.B1(n_250),
.B2(n_13),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_12),
.B(n_13),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_0),
.Y(n_257)
);


endmodule