module fake_jpeg_27563_n_227 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_36),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_0),
.CON(n_37),
.SN(n_37)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_0),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_20),
.B(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_58),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_18),
.B1(n_33),
.B2(n_32),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_32),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_40),
.B1(n_38),
.B2(n_29),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_57),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_26),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_17),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_43),
.C(n_34),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_67),
.Y(n_100)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_78),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_29),
.A3(n_26),
.B1(n_19),
.B2(n_28),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_57),
.A3(n_62),
.B1(n_46),
.B2(n_59),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_72),
.B(n_89),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_77),
.B1(n_90),
.B2(n_48),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_40),
.B1(n_38),
.B2(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_50),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_31),
.C(n_34),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_84),
.C(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_87),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_29),
.B1(n_22),
.B2(n_31),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_88),
.B1(n_42),
.B2(n_30),
.Y(n_103)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_34),
.B1(n_31),
.B2(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_30),
.B1(n_34),
.B2(n_17),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_101),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_98),
.B1(n_99),
.B2(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_46),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_97),
.B(n_108),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_65),
.B1(n_48),
.B2(n_23),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_30),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_78),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_21),
.B(n_55),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_80),
.B(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_61),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_81),
.B1(n_87),
.B2(n_67),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_1),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_1),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_96),
.B(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_124),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_80),
.C(n_74),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_127),
.C(n_98),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_74),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_83),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_123),
.B1(n_132),
.B2(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_114),
.A2(n_85),
.B1(n_2),
.B2(n_4),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_1),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_85),
.C(n_4),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_134),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_5),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_8),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_145),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_141),
.B(n_144),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_101),
.B(n_110),
.C(n_112),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_108),
.B1(n_103),
.B2(n_94),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_117),
.B1(n_119),
.B2(n_132),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_112),
.B(n_110),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_159),
.Y(n_160)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_94),
.C(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_92),
.C(n_6),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_5),
.C(n_7),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_131),
.B1(n_123),
.B2(n_132),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_115),
.B1(n_127),
.B2(n_131),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_169),
.B1(n_141),
.B2(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_155),
.B1(n_141),
.B2(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_173),
.A2(n_171),
.B1(n_177),
.B2(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_135),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_159),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_142),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_178),
.B(n_182),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_153),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_169),
.B(n_167),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_150),
.C(n_146),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_188),
.C(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_190),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_141),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_188),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_179),
.B(n_182),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_178),
.C(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_186),
.B(n_184),
.C(n_187),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_165),
.B1(n_173),
.B2(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_194),
.C(n_193),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_206),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_195),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_189),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_196),
.A2(n_147),
.B(n_11),
.C(n_12),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_209),
.B(n_198),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_192),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_204),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_193),
.C(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_216),
.B(n_217),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_207),
.B1(n_11),
.B2(n_12),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_211),
.B(n_215),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_215),
.B(n_13),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_10),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_220),
.B1(n_224),
.B2(n_13),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_14),
.Y(n_227)
);


endmodule