module fake_jpeg_20501_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_37),
.B2(n_43),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_43),
.B1(n_39),
.B2(n_36),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_25),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_57),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_26),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_33),
.B1(n_32),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_62),
.A2(n_74),
.B1(n_42),
.B2(n_40),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_68),
.Y(n_116)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_66),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_21),
.B(n_23),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_25),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_48),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_71),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_23),
.B1(n_16),
.B2(n_18),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_76),
.B1(n_80),
.B2(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_16),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_79),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_33),
.B1(n_32),
.B2(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_77),
.Y(n_108)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_18),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_32),
.B1(n_33),
.B2(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_85),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_30),
.B1(n_28),
.B2(n_19),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_89),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_30),
.B1(n_28),
.B2(n_19),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_31),
.B1(n_20),
.B2(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_95),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_104),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_69),
.B(n_74),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_99),
.A2(n_120),
.B(n_34),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_66),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_85),
.B1(n_94),
.B2(n_65),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_42),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_42),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_115),
.B1(n_88),
.B2(n_78),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_20),
.B1(n_31),
.B2(n_29),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_40),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_121),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_40),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_38),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_70),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_34),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_102),
.Y(n_157)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_154),
.B1(n_110),
.B2(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_135),
.B1(n_139),
.B2(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_64),
.C(n_38),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_120),
.C(n_100),
.Y(n_161)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_99),
.A2(n_86),
.B1(n_88),
.B2(n_35),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_143),
.Y(n_182)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_34),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_152),
.B(n_97),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_34),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_21),
.B1(n_29),
.B2(n_24),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_150),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_104),
.B(n_125),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_122),
.B(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_153),
.Y(n_158)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_185),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_147),
.A2(n_100),
.B1(n_123),
.B2(n_109),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_175),
.B1(n_134),
.B2(n_154),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_157),
.B(n_159),
.Y(n_212)
);

AO21x2_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_143),
.B(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_164),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_136),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_178),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_168),
.C(n_173),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_165),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_112),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_122),
.C(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_172),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_137),
.B1(n_129),
.B2(n_21),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_119),
.C(n_97),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_146),
.A2(n_102),
.B1(n_29),
.B2(n_24),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_183),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_27),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_140),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_194),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_191),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_149),
.B1(n_138),
.B2(n_141),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_152),
.C(n_153),
.Y(n_195)
);

NOR4xp25_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_200),
.C(n_172),
.D(n_162),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_196),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_0),
.B(n_1),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_198),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_29),
.B1(n_24),
.B2(n_22),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_217),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_27),
.C(n_24),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_181),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_27),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_22),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_219),
.C(n_182),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_208),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_165),
.B(n_22),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_213),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_155),
.A2(n_22),
.B1(n_1),
.B2(n_0),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_217),
.B1(n_175),
.B2(n_201),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_159),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_1),
.B(n_2),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_158),
.A2(n_1),
.B(n_3),
.C(n_5),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_15),
.C(n_5),
.Y(n_219)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_162),
.B(n_163),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_228),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_229),
.B1(n_230),
.B2(n_198),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_167),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_3),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_159),
.C(n_185),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_211),
.C(n_206),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_159),
.Y(n_239)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g240 ( 
.A1(n_187),
.A2(n_185),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_261),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_193),
.B1(n_210),
.B2(n_194),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_248),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_247),
.A2(n_225),
.B(n_220),
.Y(n_283)
);

FAx1_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_206),
.CI(n_188),
.CON(n_248),
.SN(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_193),
.B1(n_196),
.B2(n_199),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_254),
.B1(n_241),
.B2(n_222),
.Y(n_278)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_208),
.Y(n_255)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_207),
.C(n_219),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_264),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_3),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_259),
.Y(n_270)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_260),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_200),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_242),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_15),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_245),
.B(n_239),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_276),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_233),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_248),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_280),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_237),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_282),
.B1(n_248),
.B2(n_224),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_222),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_243),
.B1(n_220),
.B2(n_231),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_243),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_265),
.B1(n_246),
.B2(n_256),
.Y(n_287)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_247),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_292),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_265),
.C(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_296),
.C(n_6),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_231),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_253),
.C(n_240),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_268),
.B1(n_224),
.B2(n_274),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_223),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_227),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_297),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_257),
.C(n_244),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_223),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_296),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_7),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_285),
.A2(n_273),
.B1(n_280),
.B2(n_267),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_308),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_276),
.B(n_275),
.Y(n_304)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_291),
.C(n_284),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_312),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_298),
.C(n_284),
.Y(n_312)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_7),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_305),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_315),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_8),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_317),
.B(n_307),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_303),
.A2(n_8),
.B(n_9),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_300),
.B(n_306),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_325),
.A3(n_319),
.B1(n_313),
.B2(n_314),
.C1(n_316),
.C2(n_308),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_309),
.C(n_304),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_312),
.Y(n_327)
);

AOI21xp33_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_328),
.B(n_323),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_326),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_321),
.C(n_10),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_11),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_14),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_14),
.Y(n_335)
);


endmodule