module fake_jpeg_4412_n_208 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_24),
.B1(n_30),
.B2(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_58),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_24),
.B1(n_32),
.B2(n_39),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_59),
.B1(n_60),
.B2(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_35),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_53),
.B1(n_55),
.B2(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_20),
.B1(n_28),
.B2(n_23),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_28),
.B1(n_23),
.B2(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_16),
.B1(n_15),
.B2(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_32),
.A2(n_16),
.B1(n_19),
.B2(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_38),
.C(n_36),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_75),
.C(n_73),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx4f_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_38),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_78),
.B1(n_46),
.B2(n_40),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_45),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_0),
.C(n_1),
.Y(n_113)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_59),
.B1(n_44),
.B2(n_57),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_94),
.B1(n_71),
.B2(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_48),
.B1(n_51),
.B2(n_21),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_45),
.C(n_51),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_65),
.B1(n_62),
.B2(n_48),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_101),
.B1(n_107),
.B2(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_63),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_113),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_98),
.A2(n_70),
.B1(n_68),
.B2(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_68),
.B1(n_72),
.B2(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_120),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_124),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_80),
.B1(n_84),
.B2(n_81),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_134),
.B1(n_136),
.B2(n_100),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_126),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_80),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_132),
.C(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_100),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_95),
.B(n_81),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_106),
.B(n_105),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_87),
.C(n_86),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_87),
.C(n_86),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_68),
.B1(n_82),
.B2(n_96),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_86),
.B1(n_97),
.B2(n_66),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_130),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_138),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_147),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_112),
.C(n_103),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_152),
.B1(n_133),
.B2(n_135),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_118),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_138),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_121),
.B1(n_125),
.B2(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_164),
.B1(n_166),
.B2(n_148),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_127),
.B1(n_18),
.B2(n_26),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_163),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_117),
.B1(n_97),
.B2(n_19),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_29),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_145),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_177),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_148),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_161),
.B(n_160),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_29),
.C(n_25),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_173),
.A2(n_176),
.B1(n_18),
.B2(n_29),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVxp33_ASAP7_75t_SL g184 ( 
.A(n_174),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_162),
.A2(n_151),
.B1(n_147),
.B2(n_145),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_154),
.B1(n_158),
.B2(n_155),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_22),
.B1(n_18),
.B2(n_26),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_155),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_182),
.C(n_29),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_180),
.B(n_174),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_14),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_186),
.B1(n_11),
.B2(n_2),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_185),
.B(n_1),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_175),
.A2(n_13),
.B1(n_11),
.B2(n_3),
.Y(n_186)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_189),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_167),
.B(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_190),
.B1(n_191),
.B2(n_4),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_182),
.B(n_13),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_183),
.C(n_25),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_193),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_183),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_194),
.A2(n_188),
.B(n_192),
.C(n_8),
.D(n_5),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.C(n_198),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_196),
.CI(n_7),
.CON(n_204),
.SN(n_204)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

AOI321xp33_ASAP7_75t_SL g206 ( 
.A1(n_205),
.A2(n_203),
.A3(n_204),
.B1(n_199),
.B2(n_5),
.C(n_7),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_25),
.C(n_29),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_25),
.Y(n_208)
);


endmodule