module fake_jpeg_16232_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_74),
.Y(n_88)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_57),
.B1(n_60),
.B2(n_2),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_87),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_61),
.B1(n_48),
.B2(n_62),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_49),
.B1(n_52),
.B2(n_51),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_51),
.B1(n_52),
.B2(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_80),
.B1(n_92),
.B2(n_84),
.Y(n_102)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_56),
.C(n_63),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_65),
.CON(n_106),
.SN(n_106)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_0),
.Y(n_108)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_99),
.Y(n_119)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_113),
.B1(n_56),
.B2(n_47),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_103),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_111),
.B1(n_4),
.B2(n_5),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g118 ( 
.A(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_64),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_55),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_24),
.B1(n_46),
.B2(n_44),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_116),
.B1(n_123),
.B2(n_124),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_106),
.B(n_7),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_6),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_102),
.B1(n_96),
.B2(n_95),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_23),
.B1(n_42),
.B2(n_41),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_126),
.A2(n_129),
.B(n_130),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_103),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_128),
.A2(n_123),
.B1(n_115),
.B2(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

AO22x1_ASAP7_75t_SL g136 ( 
.A1(n_128),
.A2(n_117),
.B1(n_114),
.B2(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_117),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_29),
.B(n_43),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_139),
.B(n_25),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_138),
.B(n_136),
.Y(n_142)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_134),
.C(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_150),
.A2(n_151),
.B1(n_144),
.B2(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_144),
.C(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_118),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_22),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_31),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_21),
.C(n_39),
.Y(n_157)
);

OAI21x1_ASAP7_75t_SL g158 ( 
.A1(n_157),
.A2(n_20),
.B(n_37),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_13),
.B(n_36),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_12),
.B(n_34),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_33),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_118),
.C(n_32),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_107),
.C(n_9),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_8),
.Y(n_164)
);


endmodule