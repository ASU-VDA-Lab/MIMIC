module fake_jpeg_8629_n_335 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_SL g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_16),
.Y(n_71)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_76),
.Y(n_91)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_58),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_38),
.B1(n_37),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_55),
.A2(n_37),
.B1(n_31),
.B2(n_25),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_56),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_46),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_59),
.B(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_20),
.B1(n_36),
.B2(n_30),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_77),
.B1(n_17),
.B2(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_69),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_24),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_23),
.C(n_27),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_18),
.B1(n_36),
.B2(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_37),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_35),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_39),
.B(n_18),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_88),
.Y(n_129)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_17),
.B1(n_36),
.B2(n_30),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_89),
.A2(n_90),
.B(n_99),
.Y(n_137)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_17),
.B1(n_20),
.B2(n_29),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_94),
.A2(n_106),
.B1(n_109),
.B2(n_117),
.Y(n_126)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_28),
.A3(n_33),
.B1(n_32),
.B2(n_21),
.Y(n_95)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_21),
.B(n_74),
.C(n_54),
.D(n_56),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_29),
.B1(n_22),
.B2(n_24),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_103),
.Y(n_135)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_55),
.A2(n_21),
.B1(n_32),
.B2(n_26),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_113),
.B1(n_122),
.B2(n_62),
.Y(n_134)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_29),
.B1(n_33),
.B2(n_28),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_79),
.A2(n_22),
.B1(n_31),
.B2(n_25),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_120),
.B(n_13),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_123),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_22),
.B1(n_32),
.B2(n_33),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_56),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_33),
.B1(n_28),
.B2(n_31),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_60),
.A2(n_28),
.B1(n_21),
.B2(n_15),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_119),
.B1(n_83),
.B2(n_67),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_21),
.B1(n_15),
.B2(n_14),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_61),
.A2(n_15),
.B1(n_13),
.B2(n_10),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_59),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_122),
.Y(n_160)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_125),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_187)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_149),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_117),
.B(n_109),
.C(n_118),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_143),
.B1(n_145),
.B2(n_103),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_131),
.A2(n_134),
.B1(n_142),
.B2(n_3),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_56),
.C(n_61),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_138),
.C(n_110),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_83),
.B1(n_66),
.B2(n_63),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_155),
.B1(n_116),
.B2(n_114),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_80),
.B(n_1),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_151),
.B(n_156),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_74),
.B(n_62),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_88),
.B(n_122),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_95),
.A2(n_72),
.B1(n_70),
.B2(n_74),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_106),
.A2(n_72),
.B1(n_70),
.B2(n_74),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_0),
.Y(n_146)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_97),
.B(n_72),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_0),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_152),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_91),
.A2(n_70),
.B(n_2),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_105),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_108),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_154),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_91),
.A2(n_113),
.B1(n_121),
.B2(n_101),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_122),
.A2(n_0),
.B(n_2),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_86),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_158),
.Y(n_183)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_160),
.B(n_134),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_161),
.A2(n_171),
.B(n_137),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_101),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_162),
.A2(n_144),
.B(n_146),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_SL g214 ( 
.A1(n_165),
.A2(n_156),
.B(n_124),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_182),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_92),
.B1(n_116),
.B2(n_112),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_170),
.B1(n_181),
.B2(n_187),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_104),
.B(n_114),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_174),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_186),
.C(n_141),
.Y(n_203)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_128),
.A2(n_143),
.B1(n_126),
.B2(n_131),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_185),
.Y(n_217)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_105),
.C(n_104),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_126),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_142),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_9),
.B1(n_5),
.B2(n_6),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_8),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_162),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_195),
.C(n_203),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_196),
.B(n_199),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_156),
.B(n_137),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_197),
.A2(n_200),
.B(n_216),
.Y(n_227)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_177),
.B1(n_163),
.B2(n_180),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_153),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_206),
.B(n_209),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_167),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_219),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_132),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_190),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_223),
.B1(n_188),
.B2(n_184),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_163),
.B(n_139),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_221),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_147),
.B(n_157),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_161),
.A2(n_124),
.B1(n_154),
.B2(n_149),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_218),
.A2(n_222),
.B1(n_164),
.B2(n_125),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_172),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_144),
.B(n_148),
.Y(n_222)
);

XOR2x2_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_140),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_224),
.B(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_181),
.B1(n_165),
.B2(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_238),
.C(n_203),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_228),
.B(n_232),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_179),
.B1(n_178),
.B2(n_177),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_229),
.B1(n_218),
.B2(n_241),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_164),
.B1(n_174),
.B2(n_158),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_234),
.B(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_169),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_164),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_247),
.B(n_219),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_201),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_175),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_244),
.Y(n_264)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_201),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_248),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_125),
.B1(n_6),
.B2(n_7),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_199),
.B(n_205),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_223),
.C(n_216),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_249),
.B(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_215),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_256),
.B(n_263),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_229),
.A2(n_197),
.B(n_200),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_258),
.B(n_268),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_240),
.C(n_193),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_195),
.C(n_206),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_205),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_266),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_230),
.B(n_208),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_221),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_269),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_230),
.A2(n_208),
.B(n_204),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_231),
.B(n_196),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_279),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_245),
.CI(n_227),
.CON(n_272),
.SN(n_272)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_240),
.C(n_238),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_280),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_248),
.B(n_227),
.C(n_246),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_282),
.B(n_259),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_224),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_226),
.C(n_239),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_253),
.A2(n_225),
.B(n_244),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_243),
.C(n_211),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_258),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_250),
.A2(n_234),
.B1(n_198),
.B2(n_204),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_287),
.B1(n_262),
.B2(n_198),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_250),
.A2(n_198),
.B1(n_212),
.B2(n_247),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_276),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_294),
.C(n_299),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_259),
.B1(n_283),
.B2(n_278),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_292),
.B(n_293),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_268),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_277),
.B1(n_254),
.B2(n_282),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_256),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_266),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_300),
.A2(n_273),
.B(n_277),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_273),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_305),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_310),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_274),
.C(n_270),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_288),
.C(n_294),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_308),
.A2(n_301),
.B1(n_254),
.B2(n_298),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_251),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_276),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_319),
.B(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_311),
.Y(n_320)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_309),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_295),
.B(n_277),
.C(n_249),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_306),
.B(n_251),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_249),
.B1(n_272),
.B2(n_212),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_288),
.C(n_299),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_321),
.B(n_322),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_317),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_236),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_315),
.B(n_316),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_316),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_304),
.C(n_312),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

NAND3xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_331),
.C(n_329),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_319),
.B1(n_327),
.B2(n_290),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_314),
.Y(n_335)
);


endmodule