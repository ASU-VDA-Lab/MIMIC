module real_jpeg_6329_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g128 ( 
.A(n_0),
.Y(n_128)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_56),
.B1(n_60),
.B2(n_64),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_64),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_3),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_3),
.Y(n_162)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_3),
.Y(n_167)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_5),
.Y(n_267)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_5),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_5),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_6),
.A2(n_44),
.B1(n_79),
.B2(n_83),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_6),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_6),
.A2(n_83),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_6),
.A2(n_83),
.B1(n_311),
.B2(n_313),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_6),
.A2(n_83),
.B1(n_265),
.B2(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_7),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_7),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_8),
.A2(n_43),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_8),
.B(n_162),
.C(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_8),
.B(n_124),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_8),
.B(n_49),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_8),
.B(n_239),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_8),
.B(n_147),
.Y(n_362)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_9),
.Y(n_87)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_11),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_12),
.A2(n_170),
.B1(n_173),
.B2(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_12),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_12),
.A2(n_175),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_12),
.A2(n_175),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_13),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_13),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_14),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_14),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_14),
.A2(n_31),
.B1(n_82),
.B2(n_138),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_14),
.A2(n_138),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_14),
.A2(n_138),
.B1(n_352),
.B2(n_354),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_15),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_15),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_15),
.A2(n_95),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_15),
.A2(n_95),
.B1(n_129),
.B2(n_198),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_15),
.A2(n_95),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_16),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_16),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_16),
.A2(n_72),
.B1(n_170),
.B2(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_248),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_247),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_215),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_21),
.B(n_215),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_149),
.C(n_194),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_22),
.B(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_75),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_23),
.B(n_76),
.C(n_109),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_24),
.A2(n_45),
.B1(n_46),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_24),
.Y(n_257)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.A3(n_33),
.B1(n_35),
.B2(n_42),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_29),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_30),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_30),
.Y(n_147)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_30),
.Y(n_211)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_30),
.Y(n_229)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_SL g203 ( 
.A1(n_42),
.A2(n_43),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_43),
.B(n_84),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_43),
.A2(n_47),
.B(n_297),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_SL g357 ( 
.A1(n_43),
.A2(n_358),
.B(n_361),
.Y(n_357)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_54),
.B1(n_65),
.B2(n_68),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_47),
.A2(n_183),
.B1(n_193),
.B2(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_47),
.A2(n_292),
.B(n_297),
.Y(n_291)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_48),
.A2(n_69),
.B1(n_182),
.B2(n_192),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_48),
.A2(n_55),
.B1(n_262),
.B2(n_266),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_48),
.B(n_301),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_48),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_53),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_57),
.Y(n_302)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_59),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_60),
.B(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_63),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_63),
.Y(n_264)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22x1_ASAP7_75t_L g164 ( 
.A1(n_70),
.A2(n_161),
.B1(n_165),
.B2(n_168),
.Y(n_164)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_73),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_74),
.Y(n_243)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_74),
.Y(n_289)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_74),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_108),
.B2(n_109),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_84),
.B(n_93),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_78),
.A2(n_84),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_85),
.B(n_94),
.Y(n_207)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_86)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_103)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_102),
.A2(n_203),
.B(n_206),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_102),
.Y(n_231)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_133),
.B(n_143),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_110),
.A2(n_124),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_110),
.B(n_222),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_110),
.A2(n_143),
.B(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_111),
.A2(n_134),
.B1(n_148),
.B2(n_209),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_124),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B1(n_119),
.B2(n_122),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_115),
.Y(n_369)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_121),
.Y(n_374)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_124),
.Y(n_148)
);

AO22x2_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_131),
.Y(n_124)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_126),
.Y(n_286)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_126),
.Y(n_312)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_127),
.Y(n_353)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_128),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_130),
.Y(n_315)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g366 ( 
.A1(n_139),
.A2(n_352),
.A3(n_362),
.B1(n_367),
.B2(n_370),
.Y(n_366)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_142),
.Y(n_226)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_142),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_148),
.A2(n_209),
.B(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_149),
.A2(n_150),
.B1(n_194),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_181),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_151),
.B(n_181),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_164),
.B1(n_169),
.B2(n_176),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_152),
.A2(n_279),
.B(n_283),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_152),
.A2(n_164),
.B1(n_310),
.B2(n_351),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_152),
.A2(n_283),
.B(n_351),
.Y(n_381)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_153),
.A2(n_177),
.B1(n_237),
.B2(n_239),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_164),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_158),
.B1(n_161),
.B2(n_163),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_157),
.Y(n_354)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_169),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_164),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_164),
.A2(n_196),
.B(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g370 ( 
.A(n_178),
.B(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_187),
.Y(n_296)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_189),
.Y(n_265)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_193),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_193),
.A2(n_332),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_194),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.C(n_208),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_195),
.B(n_208),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_197),
.B(n_239),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_201),
.A2(n_202),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_235),
.B1(n_245),
.B2(n_246),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_230),
.B1(n_233),
.B2(n_234),
.Y(n_220)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_238),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_272),
.B(n_393),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_269),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_251),
.B(n_269),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_258),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_252),
.B(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_253),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_258),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.C(n_268),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_259),
.B(n_384),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_261),
.B(n_268),
.Y(n_384)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_262),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_263),
.Y(n_293)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI21x1_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_387),
.B(n_392),
.Y(n_272)
);

AO21x1_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_376),
.B(n_386),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_345),
.B(n_375),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_318),
.B(n_344),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_290),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_290),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_278),
.A2(n_284),
.B1(n_285),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_307),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_308),
.C(n_317),
.Y(n_346)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_316),
.B2(n_317),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_335),
.B(n_343),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_324),
.B(n_334),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_333),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_333),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_329),
.B(n_332),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_326),
.Y(n_337)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_336),
.B(n_341),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_347),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_363),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_355),
.B2(n_356),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_355),
.C(n_363),
.Y(n_377)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_366),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx8_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_377),
.B(n_378),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_380),
.B1(n_383),
.B2(n_385),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_382),
.C(n_385),
.Y(n_388)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_383),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_388),
.B(n_389),
.Y(n_392)
);


endmodule