module fake_jpeg_3620_n_681 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_681);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_681;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_64),
.B(n_71),
.Y(n_150)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_9),
.C(n_1),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_67),
.B(n_0),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_68),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_69),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_70),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_72),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_26),
.B(n_9),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_74),
.B(n_82),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_10),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_77),
.B(n_81),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_78),
.Y(n_174)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_10),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_26),
.B(n_10),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_87),
.B(n_93),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_10),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_96),
.Y(n_144)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_90),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_92),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_23),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_94),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_23),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_95),
.B(n_97),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_47),
.B(n_8),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_98),
.B(n_101),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_54),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_99),
.B(n_103),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_100),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_8),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_106),
.Y(n_218)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_54),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_111),
.B(n_122),
.Y(n_184)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_11),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_130),
.Y(n_167)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_115),
.Y(n_221)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_30),
.Y(n_116)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_20),
.Y(n_118)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_34),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_20),
.Y(n_121)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_34),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_34),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_125),
.B(n_126),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_57),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_20),
.Y(n_127)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_38),
.Y(n_129)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_51),
.B(n_7),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_20),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_131),
.B(n_132),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_40),
.B(n_0),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_75),
.A2(n_35),
.B1(n_36),
.B2(n_44),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_133),
.A2(n_151),
.B1(n_160),
.B2(n_178),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_134),
.B(n_180),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_67),
.A2(n_56),
.B1(n_40),
.B2(n_48),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_141),
.A2(n_182),
.B1(n_183),
.B2(n_192),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_75),
.A2(n_35),
.B1(n_36),
.B2(n_44),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_44),
.B1(n_36),
.B2(n_52),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_155),
.A2(n_157),
.B1(n_163),
.B2(n_133),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_52),
.B1(n_56),
.B2(n_48),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_79),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_64),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_168),
.B(n_15),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_71),
.A2(n_41),
.B1(n_33),
.B2(n_24),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_119),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_62),
.Y(n_181)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_90),
.A2(n_41),
.B1(n_33),
.B2(n_38),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_106),
.A2(n_33),
.B1(n_24),
.B2(n_32),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_99),
.A2(n_33),
.B1(n_24),
.B2(n_32),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_185),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_83),
.Y(n_189)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_69),
.A2(n_33),
.B1(n_32),
.B2(n_22),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_103),
.A2(n_33),
.B1(n_32),
.B2(n_22),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_66),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_200),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_124),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_68),
.Y(n_238)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_102),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_80),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_85),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_102),
.Y(n_209)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_113),
.A2(n_32),
.B1(n_22),
.B2(n_4),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_210),
.A2(n_212),
.B1(n_219),
.B2(n_224),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_120),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g213 ( 
.A1(n_60),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_213),
.A2(n_215),
.B1(n_220),
.B2(n_222),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_59),
.B(n_86),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_214),
.A2(n_226),
.B(n_219),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_70),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_112),
.Y(n_217)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_217),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_126),
.A2(n_5),
.B1(n_6),
.B2(n_12),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_72),
.A2(n_6),
.B1(n_12),
.B2(n_14),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g222 ( 
.A1(n_73),
.A2(n_6),
.B1(n_12),
.B2(n_14),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_115),
.Y(n_223)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_223),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_84),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_131),
.A2(n_89),
.B1(n_65),
.B2(n_78),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_226),
.A2(n_185),
.B1(n_197),
.B2(n_151),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_116),
.B(n_15),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_144),
.C(n_138),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_178),
.A2(n_83),
.B(n_110),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_232),
.A2(n_228),
.B(n_188),
.Y(n_331)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_238),
.Y(n_349)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_146),
.Y(n_239)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_239),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_135),
.B(n_123),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_240),
.B(n_245),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_241),
.B(n_280),
.Y(n_371)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_242),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_172),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_243),
.B(n_248),
.Y(n_352)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_244),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_152),
.B(n_107),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_190),
.A2(n_100),
.B1(n_108),
.B2(n_105),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_247),
.A2(n_263),
.B1(n_269),
.B2(n_140),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_143),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_171),
.Y(n_249)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_249),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_168),
.A2(n_76),
.B(n_127),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_250),
.A2(n_316),
.B(n_145),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_158),
.B(n_117),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_251),
.B(n_259),
.Y(n_339)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_177),
.Y(n_252)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_252),
.Y(n_362)
);

AO22x1_ASAP7_75t_SL g253 ( 
.A1(n_214),
.A2(n_121),
.B1(n_118),
.B2(n_61),
.Y(n_253)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_253),
.Y(n_328)
);

AND2x2_ASAP7_75t_SL g255 ( 
.A(n_176),
.B(n_63),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_255),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_92),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_256),
.B(n_257),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_137),
.B(n_94),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_167),
.B(n_128),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_260),
.B(n_273),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_261),
.A2(n_294),
.B1(n_140),
.B2(n_164),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_157),
.A2(n_16),
.B1(n_19),
.B2(n_129),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_143),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_264),
.B(n_265),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_150),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_139),
.B(n_19),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_266),
.B(n_267),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_184),
.B(n_19),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_268),
.Y(n_354)
);

AOI22x1_ASAP7_75t_L g269 ( 
.A1(n_186),
.A2(n_218),
.B1(n_187),
.B2(n_222),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_154),
.B(n_198),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_270),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_166),
.B(n_203),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_271),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_147),
.B(n_221),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_272),
.B(n_274),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_166),
.B(n_173),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_213),
.B(n_179),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_186),
.Y(n_276)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_276),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_193),
.B(n_225),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_277),
.B(n_278),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_169),
.B(n_199),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_218),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_SL g281 ( 
.A(n_155),
.B(n_206),
.C(n_217),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_281),
.B(n_285),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_205),
.Y(n_282)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_159),
.Y(n_283)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_283),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_161),
.B(n_211),
.Y(n_285)
);

OR2x2_ASAP7_75t_SL g287 ( 
.A(n_202),
.B(n_148),
.Y(n_287)
);

AOI21xp33_ASAP7_75t_L g350 ( 
.A1(n_287),
.A2(n_307),
.B(n_309),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_153),
.B(n_174),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_288),
.B(n_291),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_136),
.B(n_160),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_290),
.B(n_292),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_153),
.B(n_174),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_136),
.B(n_187),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_159),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_293),
.Y(n_366)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_165),
.Y(n_295)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_148),
.B(n_202),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_165),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_SL g318 ( 
.A(n_297),
.B(n_298),
.C(n_304),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_191),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_142),
.Y(n_301)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_142),
.B(n_156),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_302),
.Y(n_374)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_191),
.Y(n_303)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_303),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_194),
.Y(n_304)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_208),
.Y(n_305)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_156),
.Y(n_306)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_194),
.B(n_229),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_313),
.Y(n_348)
);

OR2x2_ASAP7_75t_SL g309 ( 
.A(n_170),
.B(n_212),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_170),
.Y(n_310)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_310),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_229),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_208),
.Y(n_314)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_314),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_162),
.B(n_188),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_315),
.B(n_296),
.Y(n_369)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_210),
.A2(n_175),
.B(n_145),
.C(n_228),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_175),
.B(n_230),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_302),
.C(n_296),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_322),
.A2(n_330),
.B(n_368),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_311),
.A2(n_230),
.B1(n_164),
.B2(n_195),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_325),
.A2(n_332),
.B1(n_337),
.B2(n_343),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_290),
.A2(n_279),
.B(n_275),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_331),
.A2(n_351),
.B(n_235),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_256),
.B(n_258),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_336),
.B(n_273),
.C(n_254),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_294),
.A2(n_195),
.B1(n_311),
.B2(n_286),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_338),
.A2(n_353),
.B1(n_253),
.B2(n_317),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_286),
.A2(n_300),
.B1(n_274),
.B2(n_279),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_275),
.A2(n_232),
.B(n_250),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_257),
.A2(n_308),
.B1(n_269),
.B2(n_266),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_L g426 ( 
.A1(n_357),
.A2(n_365),
.B(n_323),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_269),
.A2(n_300),
.B1(n_267),
.B2(n_260),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_361),
.A2(n_364),
.B1(n_377),
.B2(n_355),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_255),
.A2(n_292),
.B1(n_233),
.B2(n_270),
.Y(n_364)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_235),
.Y(n_367)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_367),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_278),
.A2(n_260),
.B(n_277),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_289),
.Y(n_370)
);

INVx6_ASAP7_75t_L g418 ( 
.A(n_370),
.Y(n_418)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_272),
.Y(n_375)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_375),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_255),
.A2(n_233),
.B1(n_270),
.B2(n_309),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_326),
.B(n_234),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_380),
.B(n_385),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_352),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_382),
.B(n_399),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_383),
.A2(n_390),
.B1(n_391),
.B2(n_401),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_377),
.A2(n_343),
.B1(n_374),
.B2(n_233),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_384),
.A2(n_389),
.B(n_403),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_326),
.B(n_246),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_335),
.B(n_253),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_386),
.B(n_388),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_379),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_387),
.B(n_411),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_335),
.B(n_347),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_351),
.A2(n_316),
.B(n_233),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_338),
.A2(n_317),
.B1(n_283),
.B2(n_303),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_337),
.A2(n_295),
.B1(n_314),
.B2(n_302),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_330),
.A2(n_287),
.B(n_285),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_392),
.A2(n_428),
.B(n_324),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_299),
.Y(n_393)
);

OAI21xp33_ASAP7_75t_L g465 ( 
.A1(n_393),
.A2(n_394),
.B(n_413),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_339),
.B(n_271),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_375),
.B(n_268),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_396),
.B(n_421),
.Y(n_463)
);

MAJx2_ASAP7_75t_L g398 ( 
.A(n_327),
.B(n_271),
.C(n_285),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_426),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_356),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_400),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_328),
.A2(n_305),
.B1(n_282),
.B2(n_262),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_348),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_402),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_350),
.A2(n_347),
.B(n_322),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_336),
.B(n_252),
.C(n_249),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_407),
.C(n_357),
.Y(n_431)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_327),
.B(n_273),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_405),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_328),
.A2(n_276),
.B1(n_306),
.B2(n_301),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_406),
.A2(n_420),
.B1(n_429),
.B2(n_321),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_244),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_331),
.A2(n_242),
.B(n_239),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_409),
.A2(n_410),
.B(n_412),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_333),
.B(n_312),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_364),
.A2(n_236),
.B1(n_284),
.B2(n_237),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_349),
.B(n_312),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_374),
.A2(n_236),
.B1(n_284),
.B2(n_237),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_414),
.Y(n_453)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_354),
.Y(n_416)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

NAND2x1_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_310),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_417),
.A2(n_359),
.B(n_363),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_348),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_419),
.B(n_425),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_333),
.B(n_334),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_334),
.B(n_366),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_422),
.B(n_424),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_323),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_371),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_341),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_427),
.B(n_319),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_355),
.A2(n_324),
.B1(n_342),
.B2(n_325),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_353),
.A2(n_324),
.B1(n_323),
.B2(n_354),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_431),
.B(n_450),
.Y(n_474)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_416),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_432),
.Y(n_477)
);

AO21x1_ASAP7_75t_L g472 ( 
.A1(n_434),
.A2(n_441),
.B(n_454),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_359),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_437),
.B(n_438),
.C(n_444),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_403),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_363),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_446),
.B(n_413),
.Y(n_495)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_406),
.Y(n_447)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_447),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_423),
.B(n_318),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_397),
.Y(n_452)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_423),
.A2(n_372),
.B(n_318),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_397),
.Y(n_455)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_455),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_381),
.A2(n_345),
.B1(n_341),
.B2(n_320),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_456),
.A2(n_464),
.B1(n_467),
.B2(n_428),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_422),
.B(n_372),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_457),
.B(n_400),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_384),
.A2(n_345),
.B1(n_373),
.B2(n_378),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_459),
.A2(n_461),
.B1(n_469),
.B2(n_391),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_404),
.B(n_319),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_466),
.C(n_392),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_420),
.A2(n_373),
.B1(n_360),
.B2(n_358),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_462),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_424),
.B(n_321),
.C(n_346),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_383),
.A2(n_381),
.B1(n_429),
.B2(n_419),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_418),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_402),
.A2(n_320),
.B1(n_367),
.B2(n_376),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_410),
.A2(n_376),
.B(n_344),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_471),
.A2(n_409),
.B(n_389),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_382),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_475),
.B(n_478),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_451),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_483),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g478 ( 
.A(n_465),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_431),
.B(n_399),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_479),
.B(n_490),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_395),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_480),
.B(n_502),
.C(n_504),
.Y(n_512)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_481),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_458),
.B(n_380),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_482),
.B(n_498),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_446),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_484),
.A2(n_485),
.B1(n_494),
.B2(n_501),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_467),
.A2(n_387),
.B1(n_415),
.B2(n_386),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_487),
.A2(n_445),
.B(n_440),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_443),
.A2(n_412),
.B1(n_385),
.B2(n_396),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_488),
.A2(n_470),
.B1(n_464),
.B2(n_463),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_398),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_457),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_497),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_435),
.A2(n_411),
.B1(n_425),
.B2(n_394),
.Y(n_494)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_495),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_449),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_448),
.B(n_393),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_499),
.B(n_362),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_450),
.B(n_408),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_500),
.B(n_417),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_435),
.A2(n_392),
.B1(n_390),
.B2(n_414),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_437),
.B(n_398),
.C(n_405),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_469),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_503),
.B(n_401),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_430),
.B(n_405),
.C(n_417),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_432),
.Y(n_505)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_505),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_506),
.A2(n_427),
.B1(n_408),
.B2(n_418),
.Y(n_545)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_436),
.Y(n_507)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_507),
.Y(n_516)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_508),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_430),
.B(n_405),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_466),
.C(n_434),
.Y(n_519)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_452),
.Y(n_510)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_510),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_519),
.B(n_547),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_521),
.A2(n_531),
.B1(n_536),
.B2(n_545),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_487),
.A2(n_440),
.B(n_445),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_522),
.A2(n_523),
.B(n_525),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_479),
.B(n_442),
.C(n_444),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_524),
.B(n_538),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_472),
.A2(n_454),
.B(n_471),
.Y(n_525)
);

INVxp33_ASAP7_75t_SL g526 ( 
.A(n_481),
.Y(n_526)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_526),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_528),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_473),
.A2(n_443),
.B1(n_470),
.B2(n_447),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_529),
.A2(n_530),
.B1(n_540),
.B2(n_508),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_473),
.A2(n_492),
.B1(n_503),
.B2(n_506),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_483),
.A2(n_459),
.B1(n_456),
.B2(n_463),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_495),
.Y(n_532)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_532),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_497),
.B(n_433),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_533),
.B(n_534),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_482),
.B(n_433),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_488),
.A2(n_461),
.B1(n_453),
.B2(n_441),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_477),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_537),
.B(n_541),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_474),
.B(n_442),
.C(n_462),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_472),
.A2(n_453),
.B1(n_455),
.B2(n_468),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_474),
.B(n_344),
.C(n_346),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_476),
.B(n_408),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_542),
.B(n_520),
.Y(n_573)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_543),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_499),
.A2(n_340),
.B1(n_370),
.B2(n_362),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_546),
.A2(n_504),
.B1(n_502),
.B2(n_509),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_486),
.B(n_418),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_548),
.B(n_490),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_515),
.B(n_486),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_549),
.B(n_548),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_SL g551 ( 
.A(n_539),
.B(n_480),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_551),
.B(n_568),
.Y(n_592)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_554),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_517),
.A2(n_477),
.B1(n_507),
.B2(n_493),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_557),
.A2(n_572),
.B1(n_544),
.B2(n_554),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_511),
.B(n_505),
.Y(n_562)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_562),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_511),
.B(n_489),
.Y(n_563)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_563),
.Y(n_589)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_535),
.Y(n_564)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_564),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_565),
.B(n_571),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_566),
.A2(n_579),
.B1(n_512),
.B2(n_541),
.Y(n_588)
);

XNOR2x1_ASAP7_75t_L g568 ( 
.A(n_538),
.B(n_489),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_SL g569 ( 
.A(n_539),
.B(n_493),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_569),
.B(n_570),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_SL g570 ( 
.A(n_524),
.B(n_491),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_512),
.B(n_491),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_530),
.A2(n_496),
.B1(n_510),
.B2(n_529),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_573),
.B(n_547),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_535),
.B(n_496),
.Y(n_574)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_574),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_521),
.A2(n_531),
.B1(n_527),
.B2(n_513),
.Y(n_575)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_575),
.Y(n_598)
);

NAND4xp25_ASAP7_75t_SL g576 ( 
.A(n_536),
.B(n_546),
.C(n_543),
.D(n_525),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_576),
.B(n_519),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_540),
.B(n_522),
.Y(n_577)
);

BUFx4f_ASAP7_75t_SL g604 ( 
.A(n_577),
.Y(n_604)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_516),
.Y(n_578)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_578),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_513),
.A2(n_523),
.B1(n_514),
.B2(n_516),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_563),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_580),
.B(n_581),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_574),
.Y(n_581)
);

BUFx12f_ASAP7_75t_SL g583 ( 
.A(n_553),
.Y(n_583)
);

CKINVDCx14_ASAP7_75t_R g607 ( 
.A(n_583),
.Y(n_607)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_584),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_586),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_587),
.A2(n_603),
.B(n_558),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_588),
.B(n_568),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_556),
.B(n_514),
.Y(n_590)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_590),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_562),
.B(n_518),
.Y(n_593)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_593),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_552),
.B(n_518),
.Y(n_597)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_597),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_599),
.A2(n_601),
.B1(n_567),
.B2(n_577),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_555),
.A2(n_544),
.B1(n_567),
.B2(n_579),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_559),
.B(n_572),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_602),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_553),
.A2(n_577),
.B(n_576),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_606),
.B(n_621),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_608),
.B(n_615),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_590),
.B(n_593),
.Y(n_609)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_609),
.Y(n_629)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_611),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_595),
.B(n_571),
.C(n_560),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_612),
.B(n_618),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_588),
.B(n_560),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_603),
.A2(n_550),
.B(n_557),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_616),
.A2(n_602),
.B(n_601),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_595),
.B(n_565),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_594),
.B(n_570),
.Y(n_619)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_619),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_585),
.A2(n_569),
.B(n_561),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_594),
.B(n_561),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_622),
.B(n_604),
.Y(n_639)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_592),
.B(n_551),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_624),
.B(n_604),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_584),
.B(n_596),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_625),
.B(n_598),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_612),
.B(n_615),
.C(n_618),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_626),
.B(n_631),
.C(n_636),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_627),
.B(n_634),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_614),
.B(n_598),
.Y(n_628)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_628),
.Y(n_645)
);

AOI21x1_ASAP7_75t_L g650 ( 
.A1(n_630),
.A2(n_617),
.B(n_609),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_608),
.B(n_582),
.C(n_599),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_611),
.A2(n_582),
.B1(n_589),
.B2(n_585),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_606),
.B(n_592),
.C(n_596),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_622),
.B(n_589),
.C(n_591),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_637),
.B(n_614),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_607),
.A2(n_583),
.B(n_591),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_SL g656 ( 
.A(n_638),
.B(n_639),
.C(n_630),
.Y(n_656)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_639),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_SL g642 ( 
.A(n_620),
.B(n_604),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g652 ( 
.A(n_642),
.B(n_643),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_644),
.B(n_648),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_642),
.A2(n_616),
.B(n_610),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_646),
.A2(n_656),
.B(n_625),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_631),
.B(n_623),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_650),
.B(n_651),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_638),
.B(n_605),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_632),
.A2(n_629),
.B1(n_613),
.B2(n_633),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_653),
.B(n_655),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_633),
.B(n_619),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g657 ( 
.A(n_640),
.B(n_621),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_657),
.B(n_626),
.C(n_640),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_659),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_645),
.B(n_641),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_660),
.B(n_654),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_646),
.B(n_637),
.Y(n_661)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_661),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_647),
.B(n_634),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_662),
.B(n_666),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_SL g664 ( 
.A1(n_652),
.A2(n_635),
.B(n_636),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_664),
.B(n_654),
.C(n_650),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_649),
.A2(n_600),
.B1(n_624),
.B2(n_652),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_667),
.B(n_657),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_670),
.B(n_673),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_672),
.Y(n_674)
);

A2O1A1O1Ixp25_ASAP7_75t_L g675 ( 
.A1(n_669),
.A2(n_663),
.B(n_661),
.C(n_665),
.D(n_662),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_675),
.A2(n_668),
.B(n_658),
.Y(n_678)
);

AO21x1_ASAP7_75t_L g677 ( 
.A1(n_674),
.A2(n_671),
.B(n_668),
.Y(n_677)
);

OAI21x1_ASAP7_75t_SL g679 ( 
.A1(n_677),
.A2(n_678),
.B(n_676),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_649),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_680),
.B(n_600),
.Y(n_681)
);


endmodule