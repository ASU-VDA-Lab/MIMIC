module fake_jpeg_4366_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_33),
.B1(n_29),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_28),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_24),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_41),
.B(n_40),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_44),
.Y(n_73)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_85),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_20),
.B1(n_27),
.B2(n_19),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_29),
.B1(n_33),
.B2(n_24),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_70),
.C(n_74),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_88),
.B(n_20),
.Y(n_126)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_91),
.Y(n_123)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_37),
.C(n_42),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_37),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_95),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_33),
.B1(n_29),
.B2(n_47),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_63),
.B1(n_65),
.B2(n_49),
.Y(n_105)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_69),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_24),
.B1(n_18),
.B2(n_30),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_107)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_121),
.Y(n_133)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_49),
.B1(n_63),
.B2(n_65),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_113),
.Y(n_140)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_108),
.B(n_110),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_76),
.C(n_44),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_51),
.B1(n_54),
.B2(n_66),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_68),
.B1(n_23),
.B2(n_42),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_126),
.B1(n_127),
.B2(n_96),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_115),
.B(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_26),
.Y(n_150)
);

XNOR2x2_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_23),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_120),
.B(n_22),
.Y(n_147)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_22),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_22),
.B(n_41),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_41),
.B1(n_42),
.B2(n_20),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_129),
.A2(n_106),
.B1(n_102),
.B2(n_101),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_120),
.B1(n_118),
.B2(n_110),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_131),
.A2(n_81),
.B1(n_21),
.B2(n_35),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_138),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_136),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_146),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_109),
.C(n_111),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_86),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_145),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_46),
.C(n_44),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_148),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_21),
.B(n_35),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_17),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_96),
.B1(n_22),
.B2(n_93),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_156),
.B1(n_121),
.B2(n_116),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_114),
.B1(n_121),
.B2(n_120),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_121),
.B1(n_120),
.B2(n_105),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_159),
.A2(n_148),
.B1(n_142),
.B2(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_168),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_121),
.B1(n_108),
.B2(n_124),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_143),
.B1(n_136),
.B2(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_171),
.B1(n_182),
.B2(n_184),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_17),
.A3(n_103),
.B1(n_46),
.B2(n_45),
.Y(n_170)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_34),
.B(n_46),
.C(n_45),
.D(n_84),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_91),
.B1(n_55),
.B2(n_98),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_34),
.B(n_84),
.Y(n_198)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_137),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_21),
.A3(n_35),
.B1(n_34),
.B2(n_55),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_183),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_141),
.A2(n_69),
.B1(n_56),
.B2(n_21),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_187),
.A2(n_196),
.B1(n_210),
.B2(n_171),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_175),
.A2(n_141),
.B1(n_130),
.B2(n_147),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_188),
.A2(n_205),
.B1(n_174),
.B2(n_167),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_130),
.C(n_151),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_194),
.C(n_209),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_130),
.C(n_149),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_181),
.A2(n_154),
.B(n_142),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_198),
.B(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_45),
.B(n_34),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_163),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_213),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_165),
.B(n_179),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_211),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_186),
.C(n_180),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_0),
.C(n_1),
.Y(n_211)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_16),
.B(n_15),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_182),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_193),
.B(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_224),
.Y(n_262)
);

FAx1_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_172),
.CI(n_170),
.CON(n_222),
.SN(n_222)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_222),
.B(n_232),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_167),
.B1(n_161),
.B2(n_170),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_234),
.B1(n_202),
.B2(n_201),
.Y(n_248)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_230),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_161),
.C(n_173),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_203),
.B(n_166),
.Y(n_229)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_231),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_187),
.B(n_166),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_235),
.Y(n_254)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_190),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_240),
.A2(n_199),
.B1(n_202),
.B2(n_191),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_241),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_194),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_249),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_259),
.B1(n_260),
.B2(n_215),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_225),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_209),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_211),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_255),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_206),
.C(n_208),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_238),
.C(n_236),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_206),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_217),
.B1(n_218),
.B2(n_191),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_263),
.B1(n_230),
.B2(n_224),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_188),
.B1(n_208),
.B2(n_197),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_215),
.A2(n_183),
.B1(n_198),
.B2(n_184),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_234),
.A2(n_158),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_274),
.B(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_233),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_279),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_222),
.B1(n_221),
.B2(n_228),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_272),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_280),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_247),
.A2(n_228),
.B(n_237),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_284),
.C(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_16),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_282),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_249),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_248),
.Y(n_292)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_5),
.C(n_6),
.Y(n_284)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_271),
.B(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_295),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_244),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_298),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_251),
.B(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_245),
.C(n_258),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_265),
.C(n_260),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_272),
.B1(n_267),
.B2(n_284),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_305),
.B1(n_290),
.B2(n_6),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_286),
.A2(n_264),
.B1(n_283),
.B2(n_7),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_293),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_10),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_13),
.C(n_14),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_287),
.A2(n_15),
.B(n_10),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_311),
.B(n_312),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_317),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_285),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_311),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_12),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_294),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_321),
.A2(n_324),
.B(n_5),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_301),
.A2(n_298),
.B(n_294),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_313),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_5),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_326),
.C(n_330),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_307),
.B(n_314),
.Y(n_326)
);

NAND2x1_ASAP7_75t_SL g333 ( 
.A(n_327),
.B(n_323),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_12),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_318),
.A2(n_7),
.B(n_8),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_11),
.C(n_12),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_332),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_333),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_7),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_337),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_336),
.C(n_334),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_335),
.B(n_338),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_8),
.B(n_9),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_14),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_9),
.C(n_340),
.Y(n_344)
);


endmodule