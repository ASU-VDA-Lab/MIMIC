module fake_netlist_5_2250_n_1720 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1720);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1720;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_102),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_62),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_32),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_48),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_67),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_96),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_44),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_82),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_119),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_110),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_70),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_21),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_45),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_3),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_108),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_83),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_14),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_47),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_74),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_28),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_29),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_64),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_60),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_34),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_22),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_107),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_94),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_105),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_73),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_149),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_28),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_22),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_152),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_112),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_99),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_11),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_19),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_116),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_71),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_38),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_68),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_90),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_44),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_115),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_6),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_95),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_25),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_29),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_114),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_131),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_38),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_158),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_150),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_81),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_151),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_160),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_164),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_127),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_42),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_142),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_129),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_147),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_87),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_41),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_132),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_55),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_97),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_34),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_23),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_3),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_9),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_78),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_52),
.Y(n_250)
);

BUFx2_ASAP7_75t_SL g251 ( 
.A(n_72),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_53),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_136),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_126),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_46),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_159),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_42),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_137),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_0),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_79),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_45),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_141),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_69),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_148),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_153),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_123),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_93),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_21),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_20),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_4),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_57),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_49),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_98),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_120),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_56),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_134),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_32),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_24),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_163),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_101),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_2),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_24),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_48),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_47),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_49),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_113),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_156),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_106),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_11),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_46),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_36),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_161),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_50),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_23),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_140),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_63),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_76),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_100),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_51),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_92),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_30),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_89),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_138),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_7),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_66),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_111),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_6),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_19),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_36),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_12),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_37),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_133),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_91),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_86),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_56),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_165),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_15),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_40),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_41),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_57),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_88),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_26),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_50),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_55),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_75),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_118),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_39),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_0),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_80),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_43),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_39),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_31),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_84),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_154),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_85),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_25),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_103),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_18),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_180),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_175),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_175),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_228),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_211),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_228),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_214),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_273),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_177),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_221),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_187),
.B(n_1),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_221),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_228),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_219),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_169),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_296),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_199),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_228),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_248),
.B(n_1),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_224),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_228),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_236),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_250),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_243),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_185),
.B(n_2),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_250),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_250),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_246),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_185),
.B(n_4),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_240),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_257),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_250),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_213),
.B(n_5),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_300),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_194),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_250),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_192),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_225),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_259),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_245),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_247),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_287),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_271),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_255),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_261),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_269),
.B(n_270),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_213),
.B(n_5),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_275),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_277),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_281),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_208),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_282),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_244),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_283),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_209),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_272),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_284),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_285),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_289),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_291),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_210),
.Y(n_401)
);

INVxp33_ASAP7_75t_SL g402 ( 
.A(n_169),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_210),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_301),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_293),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_170),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_248),
.B(n_7),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_301),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_315),
.B(n_8),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_294),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_304),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_307),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_194),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_182),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_191),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_215),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_193),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_195),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_194),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_218),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_201),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_395),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_349),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_419),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_367),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_376),
.B(n_220),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_342),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_369),
.B(n_220),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_367),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_R g435 ( 
.A(n_343),
.B(n_183),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_342),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_375),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_348),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_344),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_376),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_375),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_423),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_343),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_352),
.B(n_232),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_375),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_232),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_376),
.B(n_262),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_R g451 ( 
.A(n_345),
.B(n_226),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_353),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_372),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_353),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_358),
.A2(n_266),
.B(n_265),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_361),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_361),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_345),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_359),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_347),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_418),
.B(n_262),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_363),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_354),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_416),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_339),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_366),
.B(n_265),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_420),
.B(n_266),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_366),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_416),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_354),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_365),
.B(n_207),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_401),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_360),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_360),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_R g478 ( 
.A(n_362),
.B(n_227),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_416),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_404),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_421),
.B(n_166),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_416),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_373),
.B(n_233),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_362),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_422),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_404),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_422),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_364),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_422),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_405),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_424),
.B(n_314),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_422),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_350),
.B(n_287),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_364),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_410),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_411),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_357),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_461),
.B(n_346),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_445),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_474),
.B(n_393),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_440),
.B(n_449),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_474),
.B(n_356),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_451),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_440),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_442),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_453),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_461),
.B(n_368),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_479),
.B(n_368),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_442),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_387),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_442),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_432),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_426),
.B(n_351),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_442),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_432),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_426),
.B(n_382),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_442),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_489),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_485),
.A2(n_391),
.B1(n_350),
.B2(n_414),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_433),
.A2(n_338),
.B1(n_412),
.B2(n_314),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

BUFx4f_ASAP7_75t_L g531 ( 
.A(n_467),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_430),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_433),
.B(n_371),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_428),
.B(n_325),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_489),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_436),
.Y(n_536)
);

AO22x2_ASAP7_75t_L g537 ( 
.A1(n_496),
.A2(n_325),
.B1(n_222),
.B2(n_206),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_434),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_489),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_447),
.A2(n_386),
.B1(n_378),
.B2(n_403),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_459),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_402),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_451),
.Y(n_544)
);

INVxp33_ASAP7_75t_L g545 ( 
.A(n_496),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_428),
.B(n_371),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_478),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_428),
.B(n_379),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_489),
.Y(n_549)
);

INVx4_ASAP7_75t_SL g550 ( 
.A(n_489),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_483),
.B(n_379),
.Y(n_551)
);

NAND2x1p5_ASAP7_75t_L g552 ( 
.A(n_469),
.B(n_333),
.Y(n_552)
);

INVx6_ASAP7_75t_L g553 ( 
.A(n_487),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_443),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_447),
.B(n_383),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_449),
.B(n_377),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_489),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_438),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_495),
.Y(n_559)
);

OAI22xp33_ASAP7_75t_L g560 ( 
.A1(n_435),
.A2(n_299),
.B1(n_407),
.B2(n_386),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_495),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_429),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_447),
.B(n_383),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_452),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_468),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_449),
.B(n_463),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_454),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_483),
.B(n_396),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_463),
.B(n_396),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_462),
.B(n_397),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_478),
.B(n_194),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_462),
.B(n_397),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_495),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_454),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_463),
.B(n_194),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_435),
.A2(n_339),
.B1(n_415),
.B2(n_414),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_456),
.B(n_400),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_468),
.B(n_316),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_456),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_469),
.B(n_380),
.Y(n_580)
);

AO22x2_ASAP7_75t_L g581 ( 
.A1(n_469),
.A2(n_237),
.B1(n_205),
.B2(n_212),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_457),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_494),
.B(n_216),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_494),
.B(n_316),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_494),
.B(n_400),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_495),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_495),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_431),
.B(n_316),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_468),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_468),
.B(n_316),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_467),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_457),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_458),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_458),
.B(n_406),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_467),
.B(n_406),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_468),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_495),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_460),
.B(n_413),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_465),
.B(n_316),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_460),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_464),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_455),
.A2(n_381),
.B1(n_399),
.B2(n_398),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_471),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_431),
.B(n_382),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_444),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_471),
.B(n_413),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_473),
.B(n_415),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_476),
.B(n_340),
.Y(n_611)
);

INVx8_ASAP7_75t_L g612 ( 
.A(n_477),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_441),
.B(n_229),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_486),
.B(n_370),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_450),
.B(n_341),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_455),
.A2(n_384),
.B1(n_394),
.B2(n_392),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_441),
.B(n_230),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_450),
.B(n_223),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_490),
.B(n_385),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_441),
.B(n_231),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_499),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_482),
.Y(n_622)
);

OAI22xp33_ASAP7_75t_L g623 ( 
.A1(n_498),
.A2(n_203),
.B1(n_183),
.B2(n_184),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_437),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_488),
.B(n_251),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_441),
.B(n_234),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_488),
.B(n_235),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_492),
.B(n_388),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_492),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_441),
.B(n_238),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_493),
.B(n_390),
.C(n_389),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_448),
.B(n_239),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_455),
.B(n_425),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_499),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_499),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_437),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_448),
.B(n_249),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_497),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_475),
.B(n_166),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_500),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_500),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_501),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_517),
.B(n_487),
.Y(n_643)
);

INVx8_ASAP7_75t_L g644 ( 
.A(n_612),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_607),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_509),
.B(n_167),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_532),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_555),
.B(n_374),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_565),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_551),
.B(n_568),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_633),
.A2(n_537),
.B1(n_534),
.B2(n_529),
.Y(n_651)
);

OR2x2_ASAP7_75t_SL g652 ( 
.A(n_507),
.B(n_171),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_566),
.A2(n_487),
.B(n_499),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_563),
.B(n_167),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_568),
.A2(n_286),
.B1(n_253),
.B2(n_256),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_545),
.A2(n_242),
.B1(n_267),
.B2(n_264),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_543),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_585),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_508),
.B(n_487),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_546),
.A2(n_258),
.B1(n_260),
.B2(n_263),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_508),
.B(n_448),
.Y(n_662)
);

INVx8_ASAP7_75t_L g663 ( 
.A(n_612),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_545),
.B(n_254),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_SL g665 ( 
.A(n_510),
.B(n_427),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_546),
.A2(n_298),
.B1(n_274),
.B2(n_276),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_544),
.B(n_427),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_508),
.B(n_448),
.Y(n_668)
);

AND2x6_ASAP7_75t_SL g669 ( 
.A(n_572),
.B(n_425),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_565),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g671 ( 
.A(n_533),
.B(n_184),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_548),
.B(n_280),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_612),
.B(n_292),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_548),
.B(n_297),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_569),
.A2(n_313),
.B1(n_305),
.B2(n_302),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_513),
.B(n_472),
.Y(n_676)
);

BUFx5_ASAP7_75t_L g677 ( 
.A(n_633),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_543),
.B(n_168),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_633),
.A2(n_217),
.B1(n_252),
.B2(n_268),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_589),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_589),
.B(n_279),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_572),
.A2(n_306),
.B1(n_288),
.B2(n_295),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_597),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_504),
.B(n_472),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_SL g685 ( 
.A1(n_528),
.A2(n_330),
.B1(n_324),
.B2(n_336),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_539),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_534),
.A2(n_303),
.B1(n_168),
.B2(n_179),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_577),
.B(n_172),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_597),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_613),
.A2(n_499),
.B(n_446),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_622),
.B(n_629),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_552),
.B(n_172),
.Y(n_692)
);

O2A1O1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_627),
.A2(n_502),
.B(n_501),
.C(n_475),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_595),
.B(n_609),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_524),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_638),
.B(n_484),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_537),
.A2(n_309),
.B1(n_290),
.B2(n_190),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_514),
.A2(n_176),
.B1(n_173),
.B2(n_174),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_579),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_640),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_520),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_515),
.A2(n_176),
.B1(n_173),
.B2(n_174),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_641),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_591),
.B(n_188),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_519),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_523),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_529),
.A2(n_502),
.B(n_319),
.C(n_188),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g708 ( 
.A(n_575),
.B(n_178),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_599),
.B(n_178),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_547),
.B(n_438),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_552),
.A2(n_179),
.B1(n_181),
.B2(n_186),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_536),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_538),
.B(n_484),
.Y(n_713)
);

XOR2x2_ASAP7_75t_L g714 ( 
.A(n_576),
.B(n_8),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_558),
.B(n_190),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_570),
.B(n_197),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_599),
.B(n_181),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_554),
.B(n_437),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_619),
.B(n_186),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_611),
.B(n_189),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_564),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_L g722 ( 
.A(n_562),
.B(n_481),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_596),
.B(n_197),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_575),
.B(n_189),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_567),
.B(n_466),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_574),
.B(n_466),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_582),
.B(n_466),
.Y(n_727)
);

AOI22x1_ASAP7_75t_L g728 ( 
.A1(n_537),
.A2(n_480),
.B1(n_470),
.B2(n_491),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_628),
.Y(n_729)
);

NOR3x1_ASAP7_75t_L g730 ( 
.A(n_610),
.B(n_241),
.C(n_197),
.Y(n_730)
);

O2A1O1Ixp5_ASAP7_75t_L g731 ( 
.A1(n_578),
.A2(n_571),
.B(n_606),
.C(n_603),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_560),
.B(n_198),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_579),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_SL g734 ( 
.A1(n_562),
.A2(n_503),
.B1(n_319),
.B2(n_318),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_615),
.B(n_470),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_615),
.B(n_470),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_642),
.B(n_480),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_580),
.B(n_481),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_593),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_593),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_556),
.B(n_480),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_531),
.B(n_241),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_556),
.B(n_491),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_600),
.B(n_198),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_583),
.B(n_491),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_583),
.B(n_200),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_594),
.B(n_200),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_580),
.A2(n_329),
.B1(n_337),
.B2(n_335),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_614),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_594),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_580),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_601),
.B(n_202),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_601),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_602),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_553),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_600),
.B(n_202),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_560),
.B(n_204),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_581),
.A2(n_618),
.B1(n_575),
.B2(n_605),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_610),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_628),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_581),
.A2(n_320),
.B1(n_203),
.B2(n_310),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_628),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_625),
.B(n_321),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_602),
.B(n_326),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_624),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_639),
.B(n_326),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_581),
.A2(n_320),
.B1(n_310),
.B2(n_311),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_624),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_512),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_639),
.B(n_204),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_512),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_571),
.B(n_321),
.Y(n_772)
);

INVxp33_ASAP7_75t_L g773 ( 
.A(n_541),
.Y(n_773)
);

BUFx6f_ASAP7_75t_SL g774 ( 
.A(n_506),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_625),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_636),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_617),
.B(n_337),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_636),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_620),
.B(n_335),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_625),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_623),
.B(n_334),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_626),
.B(n_334),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_630),
.B(n_312),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_627),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_623),
.B(n_329),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_632),
.B(n_312),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_618),
.A2(n_287),
.B1(n_503),
.B2(n_308),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_637),
.B(n_332),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_525),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_755),
.A2(n_561),
.B(n_540),
.Y(n_790)
);

NOR2x1_ASAP7_75t_L g791 ( 
.A(n_657),
.B(n_631),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_731),
.A2(n_643),
.B(n_650),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_680),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_701),
.B(n_608),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_694),
.B(n_605),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_695),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_694),
.B(n_616),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_677),
.B(n_616),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_651),
.A2(n_553),
.B1(n_541),
.B2(n_608),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_709),
.A2(n_588),
.B(n_635),
.C(n_598),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_SL g801 ( 
.A(n_774),
.B(n_506),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_SL g802 ( 
.A(n_774),
.B(n_542),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_699),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_653),
.A2(n_635),
.B(n_598),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_699),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_755),
.A2(n_521),
.B(n_561),
.Y(n_806)
);

AOI21x1_ASAP7_75t_L g807 ( 
.A1(n_660),
.A2(n_553),
.B(n_550),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_644),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_662),
.A2(n_540),
.B(n_621),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_680),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_668),
.A2(n_540),
.B(n_621),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_733),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_741),
.A2(n_521),
.B(n_621),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_707),
.A2(n_634),
.B(n_522),
.C(n_604),
.Y(n_814)
);

OAI21x1_ASAP7_75t_L g815 ( 
.A1(n_690),
.A2(n_789),
.B(n_684),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_733),
.Y(n_816)
);

AOI21x1_ASAP7_75t_L g817 ( 
.A1(n_745),
.A2(n_743),
.B(n_736),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_677),
.B(n_618),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_739),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_680),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_759),
.B(n_542),
.Y(n_821)
);

NAND2x1p5_ASAP7_75t_L g822 ( 
.A(n_680),
.B(n_516),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_657),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_723),
.Y(n_824)
);

AND2x2_ASAP7_75t_SL g825 ( 
.A(n_679),
.B(n_542),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_769),
.A2(n_516),
.B(n_561),
.Y(n_826)
);

AO22x1_ASAP7_75t_L g827 ( 
.A1(n_773),
.A2(n_196),
.B1(n_332),
.B2(n_331),
.Y(n_827)
);

INVx11_ASAP7_75t_L g828 ( 
.A(n_644),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_677),
.B(n_618),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_739),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_659),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_749),
.B(n_526),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_789),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_SL g834 ( 
.A1(n_672),
.A2(n_559),
.B(n_527),
.C(n_557),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_773),
.B(n_512),
.Y(n_835)
);

BUFx8_ASAP7_75t_L g836 ( 
.A(n_648),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_753),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_677),
.B(n_618),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_709),
.B(n_196),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_771),
.A2(n_735),
.B(n_676),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_677),
.B(n_651),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_717),
.A2(n_575),
.B1(n_584),
.B2(n_590),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_771),
.A2(n_592),
.B(n_535),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_771),
.A2(n_535),
.B(n_587),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_740),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_750),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_644),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_717),
.B(n_328),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_677),
.B(n_559),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_754),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_716),
.B(n_241),
.Y(n_851)
);

AND2x6_ASAP7_75t_SL g852 ( 
.A(n_781),
.B(n_311),
.Y(n_852)
);

OR2x6_ASAP7_75t_L g853 ( 
.A(n_663),
.B(n_518),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_718),
.A2(n_550),
.B(n_526),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_738),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_751),
.B(n_535),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_646),
.A2(n_527),
.B(n_557),
.C(n_328),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_691),
.A2(n_518),
.B(n_587),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_649),
.Y(n_859)
);

BUFx8_ASAP7_75t_L g860 ( 
.A(n_742),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_737),
.A2(n_518),
.B(n_587),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_722),
.B(n_518),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_646),
.B(n_575),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_784),
.B(n_587),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_784),
.B(n_535),
.Y(n_865)
);

NAND2x1p5_ASAP7_75t_L g866 ( 
.A(n_670),
.B(n_573),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_645),
.B(n_688),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_728),
.A2(n_674),
.B(n_758),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_765),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_654),
.B(n_700),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_776),
.Y(n_871)
);

AO21x1_ASAP7_75t_L g872 ( 
.A1(n_674),
.A2(n_584),
.B(n_590),
.Y(n_872)
);

OAI21xp33_ASAP7_75t_L g873 ( 
.A1(n_678),
.A2(n_318),
.B(n_327),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_647),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_696),
.A2(n_530),
.B(n_586),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_715),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_766),
.B(n_331),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_703),
.B(n_584),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_732),
.A2(n_584),
.B(n_590),
.C(n_327),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_713),
.A2(n_549),
.B(n_584),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_725),
.A2(n_146),
.B(n_145),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_738),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_726),
.A2(n_727),
.B(n_681),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_678),
.B(n_9),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_681),
.A2(n_139),
.B(n_135),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_758),
.A2(n_128),
.B1(n_125),
.B2(n_124),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_788),
.A2(n_122),
.B(n_117),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_705),
.B(n_61),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_706),
.B(n_58),
.Y(n_889)
);

O2A1O1Ixp5_ASAP7_75t_L g890 ( 
.A1(n_777),
.A2(n_59),
.B(n_12),
.C(n_13),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_659),
.B(n_10),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_720),
.B(n_719),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_744),
.A2(n_10),
.B(n_13),
.C(n_15),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_779),
.A2(n_16),
.B(n_17),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_768),
.A2(n_16),
.B(n_17),
.Y(n_895)
);

AO32x2_ASAP7_75t_L g896 ( 
.A1(n_656),
.A2(n_675),
.A3(n_711),
.B1(n_734),
.B2(n_697),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_778),
.A2(n_18),
.B(n_20),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_782),
.A2(n_26),
.B(n_27),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_744),
.A2(n_756),
.B(n_720),
.C(n_785),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_683),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_729),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_783),
.A2(n_33),
.B(n_35),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_732),
.A2(n_33),
.B(n_35),
.C(n_37),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_712),
.B(n_51),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_671),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_757),
.A2(n_54),
.B(n_664),
.C(n_785),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_689),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_777),
.A2(n_54),
.B(n_786),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_679),
.B(n_719),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_729),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_704),
.B(n_652),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_721),
.B(n_770),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_685),
.B(n_781),
.C(n_697),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_686),
.A2(n_764),
.B(n_752),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_757),
.A2(n_664),
.B(n_772),
.C(n_692),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_747),
.A2(n_746),
.B(n_724),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_756),
.A2(n_692),
.B(n_693),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_761),
.B(n_767),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_761),
.B(n_767),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_763),
.A2(n_748),
.B(n_702),
.C(n_698),
.Y(n_920)
);

NOR2x1_ASAP7_75t_L g921 ( 
.A(n_673),
.B(n_762),
.Y(n_921)
);

BUFx8_ASAP7_75t_SL g922 ( 
.A(n_673),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_663),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_763),
.A2(n_775),
.B1(n_780),
.B2(n_655),
.Y(n_924)
);

AOI21x1_ASAP7_75t_L g925 ( 
.A1(n_760),
.A2(n_673),
.B(n_714),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_760),
.A2(n_661),
.B(n_666),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_708),
.A2(n_762),
.B(n_682),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_665),
.B(n_667),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_687),
.A2(n_787),
.B(n_663),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_730),
.A2(n_669),
.B(n_710),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_680),
.Y(n_931)
);

NOR2x1_ASAP7_75t_L g932 ( 
.A(n_657),
.B(n_510),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_755),
.A2(n_660),
.B(n_662),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_SL g934 ( 
.A(n_650),
.B(n_685),
.C(n_709),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_699),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_755),
.A2(n_660),
.B(n_662),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_755),
.A2(n_660),
.B(n_662),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_755),
.A2(n_660),
.B(n_662),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_650),
.A2(n_694),
.B1(n_717),
.B2(n_709),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_653),
.A2(n_690),
.B(n_789),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_723),
.B(n_505),
.Y(n_941)
);

NOR3xp33_ASAP7_75t_L g942 ( 
.A(n_650),
.B(n_685),
.C(n_528),
.Y(n_942)
);

NOR3xp33_ASAP7_75t_L g943 ( 
.A(n_650),
.B(n_685),
.C(n_528),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_650),
.A2(n_651),
.B1(n_773),
.B2(n_717),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_699),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_650),
.A2(n_651),
.B1(n_773),
.B2(n_717),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_650),
.B(n_658),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_755),
.A2(n_660),
.B(n_662),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_644),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_650),
.B(n_694),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_755),
.A2(n_660),
.B(n_662),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_723),
.B(n_505),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_731),
.A2(n_643),
.B(n_650),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_755),
.A2(n_660),
.B(n_662),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_650),
.B(n_694),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_941),
.B(n_952),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_923),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_910),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_947),
.B(n_950),
.Y(n_959)
);

OAI21x1_ASAP7_75t_SL g960 ( 
.A1(n_841),
.A2(n_868),
.B(n_927),
.Y(n_960)
);

NOR2xp67_ASAP7_75t_L g961 ( 
.A(n_821),
.B(n_824),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_939),
.A2(n_899),
.B(n_892),
.C(n_839),
.Y(n_962)
);

AND2x6_ASAP7_75t_L g963 ( 
.A(n_841),
.B(n_798),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_950),
.B(n_955),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_851),
.B(n_942),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_955),
.B(n_848),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_795),
.B(n_797),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_793),
.Y(n_968)
);

CKINVDCx6p67_ASAP7_75t_R g969 ( 
.A(n_808),
.Y(n_969)
);

AOI21xp33_ASAP7_75t_L g970 ( 
.A1(n_884),
.A2(n_913),
.B(n_944),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_SL g971 ( 
.A1(n_943),
.A2(n_909),
.B(n_934),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_933),
.A2(n_937),
.B(n_936),
.Y(n_972)
);

OAI22x1_ASAP7_75t_L g973 ( 
.A1(n_918),
.A2(n_919),
.B1(n_924),
.B2(n_925),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_795),
.B(n_797),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_946),
.B(n_912),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_938),
.A2(n_948),
.B(n_951),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_803),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_940),
.A2(n_815),
.B(n_854),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_831),
.B(n_876),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_792),
.A2(n_953),
.B(n_834),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_951),
.A2(n_954),
.B(n_790),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_870),
.B(n_912),
.Y(n_982)
);

NAND2x1_ASAP7_75t_L g983 ( 
.A(n_833),
.B(n_793),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_915),
.A2(n_906),
.B(n_920),
.C(n_917),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_954),
.A2(n_790),
.B(n_849),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_804),
.A2(n_811),
.B(n_813),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_901),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_825),
.A2(n_799),
.B1(n_867),
.B2(n_918),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_870),
.B(n_864),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_796),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_823),
.B(n_794),
.Y(n_991)
);

AOI21xp33_ASAP7_75t_L g992 ( 
.A1(n_919),
.A2(n_897),
.B(n_895),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_823),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_891),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_849),
.A2(n_798),
.B(n_806),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_823),
.B(n_855),
.Y(n_996)
);

O2A1O1Ixp5_ASAP7_75t_L g997 ( 
.A1(n_863),
.A2(n_916),
.B(n_857),
.C(n_872),
.Y(n_997)
);

AOI21xp33_ASAP7_75t_L g998 ( 
.A1(n_873),
.A2(n_903),
.B(n_911),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_883),
.A2(n_840),
.B(n_809),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_793),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_818),
.A2(n_838),
.B(n_829),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_886),
.A2(n_904),
.B1(n_893),
.B2(n_908),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_928),
.B(n_882),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_817),
.A2(n_914),
.B(n_818),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_905),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_810),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_904),
.A2(n_865),
.B1(n_864),
.B2(n_889),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_829),
.A2(n_838),
.B(n_826),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_865),
.B(n_832),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_810),
.Y(n_1010)
);

CKINVDCx16_ASAP7_75t_R g1011 ( 
.A(n_801),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_800),
.A2(n_858),
.B(n_843),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_822),
.A2(n_835),
.B(n_862),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_861),
.A2(n_814),
.B(n_875),
.Y(n_1014)
);

AOI221xp5_ASAP7_75t_SL g1015 ( 
.A1(n_894),
.A2(n_898),
.B1(n_902),
.B2(n_887),
.C(n_846),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_810),
.B(n_932),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_877),
.B(n_827),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_907),
.B(n_859),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_805),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_930),
.B(n_921),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_822),
.A2(n_844),
.B(n_878),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_907),
.A2(n_850),
.B1(n_791),
.B2(n_837),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_888),
.A2(n_889),
.B1(n_900),
.B2(n_929),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_896),
.B(n_845),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_896),
.B(n_802),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_812),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_820),
.B(n_931),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_931),
.B(n_945),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_842),
.A2(n_833),
.B1(n_819),
.B2(n_830),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_926),
.A2(n_879),
.B(n_890),
.C(n_878),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_856),
.A2(n_880),
.B(n_853),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_816),
.B(n_935),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_869),
.A2(n_874),
.B(n_871),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_853),
.A2(n_885),
.B(n_866),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_866),
.B(n_847),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_881),
.A2(n_923),
.B(n_828),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_860),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_923),
.A2(n_949),
.B(n_896),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_852),
.A2(n_860),
.B1(n_836),
.B2(n_922),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_836),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_950),
.B(n_955),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_940),
.A2(n_815),
.B(n_807),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_SL g1043 ( 
.A1(n_899),
.A2(n_755),
.B(n_798),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_941),
.B(n_952),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_SL g1045 ( 
.A1(n_913),
.A2(n_943),
.B(n_942),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_950),
.B(n_955),
.Y(n_1046)
);

AO31x2_ASAP7_75t_L g1047 ( 
.A1(n_899),
.A2(n_857),
.A3(n_946),
.B(n_944),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_940),
.A2(n_815),
.B(n_807),
.Y(n_1048)
);

AND3x2_ASAP7_75t_L g1049 ( 
.A(n_801),
.B(n_802),
.C(n_884),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_796),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_950),
.B(n_955),
.Y(n_1051)
);

NOR2x1_ASAP7_75t_SL g1052 ( 
.A(n_853),
.B(n_923),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_934),
.A2(n_939),
.B1(n_943),
.B2(n_942),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_950),
.B(n_955),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_939),
.A2(n_899),
.B(n_944),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_831),
.Y(n_1056)
);

NAND2xp33_ASAP7_75t_L g1057 ( 
.A(n_899),
.B(n_939),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_950),
.B(n_955),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_831),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_939),
.A2(n_899),
.B(n_944),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_939),
.A2(n_899),
.B(n_944),
.Y(n_1061)
);

OAI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_839),
.A2(n_650),
.B(n_848),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_941),
.B(n_952),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_939),
.A2(n_899),
.B(n_944),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_950),
.B(n_955),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_950),
.B(n_955),
.Y(n_1066)
);

XOR2xp5_ASAP7_75t_L g1067 ( 
.A(n_934),
.B(n_438),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_950),
.B(n_955),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_R g1069 ( 
.A(n_934),
.B(n_562),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_823),
.B(n_855),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_939),
.A2(n_899),
.B(n_892),
.C(n_650),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_950),
.B(n_955),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_933),
.A2(n_755),
.B(n_936),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_899),
.A2(n_857),
.A3(n_946),
.B(n_944),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_939),
.A2(n_899),
.B(n_944),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_939),
.A2(n_950),
.B1(n_955),
.B2(n_650),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_950),
.B(n_955),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_950),
.B(n_955),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_950),
.B(n_955),
.Y(n_1079)
);

NAND2x1p5_ASAP7_75t_L g1080 ( 
.A(n_923),
.B(n_847),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_803),
.Y(n_1081)
);

OAI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_839),
.A2(n_650),
.B(n_848),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_941),
.B(n_952),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_933),
.A2(n_755),
.B(n_936),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_939),
.A2(n_899),
.B(n_892),
.C(n_650),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_950),
.B(n_955),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_947),
.B(n_650),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_823),
.B(n_855),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_939),
.A2(n_899),
.B(n_944),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_939),
.A2(n_950),
.B1(n_955),
.B2(n_650),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_962),
.A2(n_1062),
.B(n_1082),
.C(n_966),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_958),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_976),
.A2(n_972),
.B(n_999),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_1087),
.B(n_959),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_956),
.B(n_1044),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_996),
.B(n_1070),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1063),
.B(n_1083),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_957),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_977),
.Y(n_1099)
);

NAND2x1p5_ASAP7_75t_L g1100 ( 
.A(n_957),
.B(n_968),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_965),
.A2(n_1053),
.B1(n_1045),
.B2(n_1057),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1019),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_996),
.B(n_1070),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_968),
.Y(n_1104)
);

BUFx12f_ASAP7_75t_L g1105 ( 
.A(n_1040),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1081),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_968),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_964),
.B(n_1041),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_982),
.B(n_979),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1046),
.B(n_1051),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_990),
.Y(n_1111)
);

INVx3_ASAP7_75t_SL g1112 ( 
.A(n_969),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1088),
.B(n_993),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1054),
.B(n_1058),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1065),
.B(n_1066),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_1059),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1032),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1073),
.A2(n_1084),
.B(n_981),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1068),
.A2(n_1072),
.B1(n_1077),
.B2(n_1079),
.Y(n_1119)
);

CKINVDCx16_ASAP7_75t_R g1120 ( 
.A(n_1040),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_994),
.B(n_1059),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1040),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1088),
.B(n_991),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1020),
.B(n_994),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1050),
.B(n_1003),
.Y(n_1125)
);

OA21x2_ASAP7_75t_L g1126 ( 
.A1(n_980),
.A2(n_986),
.B(n_978),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1078),
.B(n_1086),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1086),
.A2(n_1071),
.B1(n_1085),
.B2(n_1090),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_970),
.A2(n_1060),
.B(n_1055),
.C(n_1089),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1076),
.B(n_1090),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1000),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_985),
.A2(n_1043),
.B(n_984),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1055),
.A2(n_1089),
.B(n_1075),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_961),
.B(n_1005),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1000),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1076),
.B(n_1056),
.Y(n_1136)
);

BUFx4_ASAP7_75t_SL g1137 ( 
.A(n_1037),
.Y(n_1137)
);

BUFx10_ASAP7_75t_L g1138 ( 
.A(n_1049),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1060),
.A2(n_1064),
.B(n_1061),
.Y(n_1139)
);

OR2x6_ASAP7_75t_SL g1140 ( 
.A(n_1039),
.B(n_975),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_989),
.B(n_974),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_971),
.B(n_987),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1037),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_973),
.B(n_1017),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1016),
.B(n_1052),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1061),
.A2(n_1075),
.B1(n_1064),
.B2(n_975),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_988),
.A2(n_974),
.B1(n_967),
.B2(n_1024),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_995),
.A2(n_1012),
.B(n_1023),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1000),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1028),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_963),
.B(n_970),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_998),
.B(n_1023),
.C(n_992),
.Y(n_1152)
);

OR2x6_ASAP7_75t_SL g1153 ( 
.A(n_1039),
.B(n_1035),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1034),
.A2(n_1008),
.B(n_1007),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1080),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_960),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_1006),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_992),
.B(n_1080),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1018),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1025),
.B(n_1069),
.Y(n_1160)
);

AOI222xp33_ASAP7_75t_L g1161 ( 
.A1(n_1002),
.A2(n_963),
.B1(n_1022),
.B2(n_1033),
.C1(n_980),
.C2(n_1009),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_998),
.B(n_1047),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1027),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1002),
.B(n_1010),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1006),
.B(n_1010),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_983),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1036),
.B(n_1038),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1029),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1047),
.B(n_1074),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_963),
.B(n_1074),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_963),
.B(n_1074),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1029),
.B(n_1013),
.Y(n_1172)
);

INVx5_ASAP7_75t_L g1173 ( 
.A(n_997),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1047),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1031),
.B(n_1001),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1015),
.B(n_1030),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1021),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1004),
.Y(n_1178)
);

BUFx4f_ASAP7_75t_SL g1179 ( 
.A(n_1015),
.Y(n_1179)
);

INVx3_ASAP7_75t_SL g1180 ( 
.A(n_1014),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1042),
.B(n_1048),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_956),
.B(n_1044),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_976),
.A2(n_972),
.B(n_999),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_966),
.A2(n_899),
.B(n_939),
.C(n_1062),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_SL g1185 ( 
.A1(n_966),
.A2(n_884),
.B(n_848),
.C(n_839),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_959),
.B(n_950),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_996),
.B(n_1070),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_957),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_968),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_982),
.B(n_558),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_962),
.A2(n_650),
.B(n_899),
.C(n_1062),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_977),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1011),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_982),
.B(n_558),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_959),
.B(n_950),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_958),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_958),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_958),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_976),
.A2(n_972),
.B(n_999),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1059),
.Y(n_1200)
);

INVxp33_ASAP7_75t_L g1201 ( 
.A(n_958),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1062),
.A2(n_943),
.B1(n_942),
.B2(n_913),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_957),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_958),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_968),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1026),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_957),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1062),
.B(n_531),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_958),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_996),
.B(n_1070),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_966),
.A2(n_825),
.B1(n_913),
.B2(n_650),
.Y(n_1211)
);

HAxp5_ASAP7_75t_L g1212 ( 
.A(n_1067),
.B(n_671),
.CON(n_1212),
.SN(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_959),
.B(n_950),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_958),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_958),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_958),
.Y(n_1216)
);

XNOR2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1039),
.B(n_562),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_959),
.B(n_950),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_957),
.B(n_923),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_996),
.B(n_1070),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1059),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_959),
.B(n_950),
.Y(n_1222)
);

INVx5_ASAP7_75t_SL g1223 ( 
.A(n_1040),
.Y(n_1223)
);

NOR2xp67_ASAP7_75t_L g1224 ( 
.A(n_1005),
.B(n_759),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1087),
.A2(n_939),
.B1(n_955),
.B2(n_950),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1026),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_966),
.B(n_650),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_956),
.B(n_1044),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1099),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1094),
.A2(n_1227),
.B1(n_1142),
.B2(n_1101),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1106),
.Y(n_1231)
);

AO21x2_ASAP7_75t_L g1232 ( 
.A1(n_1148),
.A2(n_1154),
.B(n_1118),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1202),
.A2(n_1211),
.B1(n_1115),
.B2(n_1136),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1127),
.A2(n_1195),
.B1(n_1213),
.B2(n_1218),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1193),
.A2(n_1120),
.B1(n_1186),
.B2(n_1213),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1159),
.Y(n_1236)
);

INVx6_ASAP7_75t_L g1237 ( 
.A(n_1157),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1146),
.A2(n_1139),
.B1(n_1133),
.B2(n_1225),
.Y(n_1238)
);

BUFx8_ASAP7_75t_L g1239 ( 
.A(n_1105),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1132),
.B(n_1124),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1156),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1102),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1192),
.Y(n_1243)
);

CKINVDCx16_ASAP7_75t_R g1244 ( 
.A(n_1122),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1134),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1128),
.Y(n_1246)
);

INVx6_ASAP7_75t_L g1247 ( 
.A(n_1134),
.Y(n_1247)
);

BUFx4f_ASAP7_75t_L g1248 ( 
.A(n_1112),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_1138),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1093),
.A2(n_1199),
.B(n_1183),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1146),
.A2(n_1133),
.B1(n_1139),
.B2(n_1225),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1186),
.B(n_1195),
.Y(n_1252)
);

BUFx2_ASAP7_75t_R g1253 ( 
.A(n_1153),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1174),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1206),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1200),
.Y(n_1256)
);

BUFx2_ASAP7_75t_R g1257 ( 
.A(n_1140),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1218),
.A2(n_1222),
.B1(n_1110),
.B2(n_1108),
.Y(n_1258)
);

BUFx8_ASAP7_75t_L g1259 ( 
.A(n_1092),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1152),
.A2(n_1128),
.B1(n_1179),
.B2(n_1222),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1104),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1116),
.Y(n_1262)
);

BUFx2_ASAP7_75t_R g1263 ( 
.A(n_1197),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1152),
.A2(n_1144),
.B1(n_1208),
.B2(n_1119),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1108),
.B(n_1110),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1124),
.B(n_1164),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1119),
.A2(n_1114),
.B1(n_1161),
.B2(n_1162),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1138),
.A2(n_1160),
.B1(n_1158),
.B2(n_1114),
.Y(n_1268)
);

BUFx4f_ASAP7_75t_SL g1269 ( 
.A(n_1204),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1178),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1226),
.Y(n_1271)
);

BUFx8_ASAP7_75t_L g1272 ( 
.A(n_1198),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1217),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1184),
.A2(n_1129),
.B1(n_1190),
.B2(n_1194),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1095),
.B(n_1097),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1141),
.A2(n_1109),
.B1(n_1177),
.B2(n_1091),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1141),
.A2(n_1224),
.B1(n_1221),
.B2(n_1116),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1161),
.A2(n_1151),
.B1(n_1147),
.B2(n_1172),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1150),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1182),
.B(n_1228),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1117),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1221),
.A2(n_1125),
.B1(n_1191),
.B2(n_1196),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1163),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_SL g1284 ( 
.A1(n_1175),
.A2(n_1147),
.B(n_1219),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1151),
.A2(n_1168),
.B1(n_1176),
.B2(n_1121),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1209),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1137),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1176),
.A2(n_1125),
.B1(n_1169),
.B2(n_1123),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1178),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1185),
.B(n_1187),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1096),
.B(n_1187),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1100),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1104),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1149),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1104),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_SL g1296 ( 
.A(n_1143),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1173),
.A2(n_1170),
.B1(n_1171),
.B2(n_1175),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1214),
.A2(n_1201),
.B1(n_1215),
.B2(n_1216),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1111),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1170),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1096),
.B(n_1103),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1145),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1103),
.A2(n_1210),
.B1(n_1220),
.B2(n_1158),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1212),
.B(n_1220),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1210),
.A2(n_1113),
.B1(n_1223),
.B2(n_1166),
.Y(n_1305)
);

INVx6_ASAP7_75t_L g1306 ( 
.A(n_1107),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1165),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1165),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1155),
.B(n_1098),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1131),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1131),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1131),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1135),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1223),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1173),
.A2(n_1167),
.B1(n_1180),
.B2(n_1203),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1098),
.B(n_1188),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1188),
.B(n_1203),
.Y(n_1317)
);

BUFx8_ASAP7_75t_SL g1318 ( 
.A(n_1189),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1126),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1207),
.A2(n_1189),
.B1(n_1205),
.B2(n_1181),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1094),
.A2(n_825),
.B1(n_913),
.B2(n_909),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1096),
.B(n_1103),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1095),
.B(n_1097),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1099),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1099),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1099),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1096),
.B(n_1103),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1096),
.B(n_1103),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1099),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1095),
.B(n_1097),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1094),
.A2(n_913),
.B1(n_943),
.B2(n_942),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1095),
.B(n_1097),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1094),
.A2(n_913),
.B1(n_943),
.B2(n_942),
.Y(n_1333)
);

BUFx2_ASAP7_75t_SL g1334 ( 
.A(n_1193),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1300),
.B(n_1238),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1259),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1262),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1300),
.B(n_1278),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1275),
.Y(n_1339)
);

INVxp33_ASAP7_75t_L g1340 ( 
.A(n_1280),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1230),
.A2(n_1233),
.B1(n_1331),
.B2(n_1333),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1238),
.B(n_1251),
.Y(n_1342)
);

BUFx2_ASAP7_75t_SL g1343 ( 
.A(n_1296),
.Y(n_1343)
);

CKINVDCx6p67_ASAP7_75t_R g1344 ( 
.A(n_1314),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1240),
.Y(n_1345)
);

AND2x4_ASAP7_75t_SL g1346 ( 
.A(n_1266),
.B(n_1240),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1252),
.B(n_1265),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1277),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1323),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1278),
.B(n_1267),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1267),
.B(n_1264),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1264),
.B(n_1251),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1252),
.B(n_1234),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1258),
.B(n_1276),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1241),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1274),
.B(n_1331),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1282),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1256),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1260),
.B(n_1240),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1319),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1333),
.A2(n_1321),
.B1(n_1268),
.B2(n_1260),
.Y(n_1361)
);

BUFx2_ASAP7_75t_SL g1362 ( 
.A(n_1296),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1319),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1281),
.B(n_1236),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1242),
.B(n_1243),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1236),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1246),
.A2(n_1250),
.B(n_1284),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1290),
.A2(n_1303),
.B(n_1304),
.C(n_1305),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1279),
.B(n_1283),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1297),
.B(n_1285),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1254),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1297),
.B(n_1285),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1254),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1266),
.B(n_1288),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1269),
.Y(n_1375)
);

AO21x2_ASAP7_75t_L g1376 ( 
.A1(n_1232),
.A2(n_1289),
.B(n_1270),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1266),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1288),
.B(n_1325),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1232),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1315),
.A2(n_1320),
.B(n_1302),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1229),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1231),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1324),
.Y(n_1383)
);

BUFx4f_ASAP7_75t_SL g1384 ( 
.A(n_1314),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1294),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1286),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1326),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1329),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1330),
.B(n_1332),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1299),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1255),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1259),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1259),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1271),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1308),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1291),
.B(n_1257),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1298),
.B(n_1235),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1301),
.B(n_1328),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1316),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1309),
.Y(n_1400)
);

NOR2x1_ASAP7_75t_L g1401 ( 
.A(n_1316),
.B(n_1317),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1307),
.A2(n_1311),
.B(n_1312),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1309),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1301),
.B(n_1328),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1249),
.A2(n_1273),
.B1(n_1334),
.B2(n_1247),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1301),
.B(n_1328),
.Y(n_1406)
);

AO21x1_ASAP7_75t_L g1407 ( 
.A1(n_1356),
.A2(n_1253),
.B(n_1310),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1376),
.Y(n_1408)
);

BUFx12f_ASAP7_75t_L g1409 ( 
.A(n_1392),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1345),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1360),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1353),
.B(n_1292),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1335),
.B(n_1322),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1345),
.Y(n_1414)
);

NOR2x1_ASAP7_75t_L g1415 ( 
.A(n_1402),
.B(n_1313),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1363),
.B(n_1335),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1355),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1341),
.A2(n_1350),
.B1(n_1361),
.B2(n_1351),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1341),
.A2(n_1273),
.B1(n_1263),
.B2(n_1245),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1379),
.B(n_1327),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1379),
.B(n_1327),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1402),
.Y(n_1422)
);

INVx5_ASAP7_75t_L g1423 ( 
.A(n_1379),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1338),
.B(n_1245),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1350),
.A2(n_1248),
.B(n_1295),
.C(n_1293),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1338),
.B(n_1245),
.Y(n_1426)
);

NAND2x1_ASAP7_75t_L g1427 ( 
.A(n_1377),
.B(n_1306),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1370),
.B(n_1372),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1370),
.B(n_1293),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1354),
.B(n_1352),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1378),
.B(n_1261),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1378),
.B(n_1261),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1352),
.B(n_1247),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1347),
.B(n_1247),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1351),
.A2(n_1249),
.B1(n_1272),
.B2(n_1269),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1346),
.B(n_1287),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1342),
.B(n_1244),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1428),
.B(n_1348),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1428),
.B(n_1359),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1430),
.B(n_1385),
.Y(n_1440)
);

OAI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1418),
.A2(n_1368),
.B1(n_1405),
.B2(n_1397),
.C(n_1396),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1431),
.B(n_1371),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1407),
.B(n_1401),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1430),
.B(n_1357),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1418),
.B(n_1397),
.C(n_1358),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1431),
.B(n_1371),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1419),
.A2(n_1346),
.B(n_1392),
.Y(n_1447)
);

AOI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1415),
.A2(n_1407),
.B(n_1427),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1431),
.B(n_1373),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1419),
.A2(n_1340),
.B1(n_1349),
.B2(n_1339),
.C(n_1390),
.Y(n_1450)
);

OAI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1435),
.A2(n_1398),
.B1(n_1404),
.B2(n_1386),
.C(n_1248),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1432),
.B(n_1373),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1412),
.B(n_1337),
.Y(n_1453)
);

OAI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1435),
.A2(n_1386),
.B1(n_1393),
.B2(n_1401),
.C(n_1343),
.Y(n_1454)
);

OAI221xp5_ASAP7_75t_L g1455 ( 
.A1(n_1425),
.A2(n_1393),
.B1(n_1362),
.B2(n_1343),
.C(n_1400),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1412),
.B(n_1388),
.Y(n_1456)
);

NAND3xp33_ASAP7_75t_L g1457 ( 
.A(n_1437),
.B(n_1387),
.C(n_1383),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1413),
.B(n_1365),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1413),
.B(n_1432),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1434),
.B(n_1344),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1437),
.B(n_1387),
.C(n_1382),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1420),
.B(n_1374),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1420),
.B(n_1402),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1413),
.B(n_1365),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1420),
.B(n_1389),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1437),
.B(n_1366),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1421),
.B(n_1389),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1429),
.B(n_1381),
.Y(n_1468)
);

OAI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1434),
.A2(n_1362),
.B1(n_1403),
.B2(n_1400),
.C(n_1336),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1433),
.A2(n_1344),
.B1(n_1336),
.B2(n_1426),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1422),
.B(n_1382),
.C(n_1383),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1421),
.B(n_1399),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1407),
.A2(n_1336),
.B1(n_1406),
.B2(n_1384),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1411),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1422),
.B(n_1394),
.C(n_1391),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1415),
.A2(n_1380),
.B(n_1367),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1424),
.A2(n_1369),
.B1(n_1395),
.B2(n_1403),
.C(n_1364),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1463),
.B(n_1408),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1474),
.B(n_1411),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1457),
.B(n_1461),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1463),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1474),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1440),
.B(n_1417),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1471),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1471),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1475),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1457),
.B(n_1436),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1472),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1444),
.B(n_1438),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1475),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1468),
.B(n_1416),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1466),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1462),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1476),
.B(n_1423),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1476),
.B(n_1410),
.Y(n_1497)
);

INVx4_ASAP7_75t_L g1498 ( 
.A(n_1442),
.Y(n_1498)
);

AND2x2_ASAP7_75t_SL g1499 ( 
.A(n_1439),
.B(n_1436),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1442),
.Y(n_1500)
);

NOR2xp67_ASAP7_75t_R g1501 ( 
.A(n_1473),
.B(n_1409),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1446),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1449),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1496),
.B(n_1448),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1481),
.B(n_1484),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1498),
.B(n_1452),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1482),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1482),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1479),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1498),
.B(n_1452),
.Y(n_1510)
);

NAND2x1_ASAP7_75t_SL g1511 ( 
.A(n_1485),
.B(n_1448),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1479),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1500),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1494),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1490),
.B(n_1453),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1499),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1500),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1489),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1519)
);

AOI21xp33_ASAP7_75t_L g1520 ( 
.A1(n_1480),
.A2(n_1470),
.B(n_1469),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1481),
.B(n_1459),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1498),
.B(n_1414),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1490),
.B(n_1456),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1498),
.B(n_1414),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1499),
.B(n_1414),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1481),
.B(n_1458),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1503),
.Y(n_1527)
);

NOR2x1_ASAP7_75t_L g1528 ( 
.A(n_1480),
.B(n_1461),
.Y(n_1528)
);

NOR2x1p5_ASAP7_75t_L g1529 ( 
.A(n_1501),
.B(n_1445),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1496),
.B(n_1436),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1499),
.B(n_1414),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1496),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1494),
.B(n_1464),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1483),
.B(n_1460),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1481),
.B(n_1484),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1503),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1502),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1507),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1519),
.B(n_1478),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1519),
.B(n_1496),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1533),
.B(n_1493),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1528),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1529),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1507),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1516),
.B(n_1478),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1514),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1521),
.B(n_1493),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1521),
.B(n_1493),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1518),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1520),
.A2(n_1445),
.B1(n_1447),
.B2(n_1454),
.Y(n_1550)
);

INVxp33_ASAP7_75t_L g1551 ( 
.A(n_1534),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1515),
.B(n_1486),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1518),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_SL g1554 ( 
.A(n_1532),
.B(n_1455),
.Y(n_1554)
);

AOI32xp33_ASAP7_75t_L g1555 ( 
.A1(n_1516),
.A2(n_1488),
.A3(n_1491),
.B1(n_1487),
.B2(n_1485),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_SL g1556 ( 
.A(n_1532),
.B(n_1447),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1496),
.Y(n_1557)
);

OAI32xp33_ASAP7_75t_L g1558 ( 
.A1(n_1532),
.A2(n_1491),
.A3(n_1488),
.B1(n_1487),
.B2(n_1443),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1523),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1526),
.B(n_1495),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1530),
.B(n_1478),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1526),
.B(n_1495),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1530),
.B(n_1486),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1508),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1509),
.B(n_1495),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1509),
.B(n_1492),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1512),
.A2(n_1441),
.B(n_1491),
.C(n_1497),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1525),
.B(n_1492),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1525),
.B(n_1492),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1504),
.B(n_1496),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1508),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1512),
.B(n_1409),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1513),
.Y(n_1573)
);

NAND3xp33_ASAP7_75t_L g1574 ( 
.A(n_1505),
.B(n_1450),
.C(n_1470),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1513),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1505),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1504),
.B(n_1497),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1517),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1531),
.B(n_1497),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1517),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1538),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1544),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1542),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1577),
.B(n_1504),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_SL g1585 ( 
.A(n_1543),
.B(n_1511),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_1554),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1546),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1577),
.B(n_1563),
.Y(n_1588)
);

INVx3_ASAP7_75t_SL g1589 ( 
.A(n_1543),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1549),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1556),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1541),
.B(n_1535),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1549),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1564),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1577),
.B(n_1531),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1553),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1563),
.B(n_1506),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1571),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1551),
.A2(n_1550),
.B1(n_1574),
.B2(n_1559),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1551),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1568),
.B(n_1506),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1568),
.B(n_1510),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1572),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1575),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1578),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1580),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1576),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1569),
.B(n_1579),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1565),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1566),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1545),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1552),
.B(n_1535),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1558),
.A2(n_1451),
.B1(n_1501),
.B2(n_1497),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1572),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1607),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1607),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1600),
.A2(n_1567),
.B(n_1511),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1608),
.Y(n_1620)
);

NOR2x1_ASAP7_75t_L g1621 ( 
.A(n_1602),
.B(n_1570),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1602),
.B(n_1547),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1588),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1588),
.B(n_1540),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1589),
.B(n_1287),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1587),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1588),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1596),
.Y(n_1628)
);

OAI31xp33_ASAP7_75t_L g1629 ( 
.A1(n_1585),
.A2(n_1555),
.A3(n_1477),
.B(n_1570),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1589),
.B(n_1583),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1608),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1601),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1601),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1583),
.B(n_1569),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1606),
.Y(n_1635)
);

AND2x6_ASAP7_75t_L g1636 ( 
.A(n_1591),
.B(n_1239),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1596),
.Y(n_1637)
);

OAI32xp33_ASAP7_75t_L g1638 ( 
.A1(n_1586),
.A2(n_1591),
.A3(n_1605),
.B1(n_1616),
.B2(n_1613),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1609),
.B(n_1548),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1606),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1586),
.A2(n_1540),
.B(n_1557),
.Y(n_1641)
);

NOR4xp25_ASAP7_75t_SL g1642 ( 
.A(n_1609),
.B(n_1537),
.C(n_1527),
.D(n_1536),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1617),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1624),
.B(n_1589),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1634),
.B(n_1613),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1618),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1620),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1634),
.B(n_1613),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1624),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1621),
.B(n_1605),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1630),
.B(n_1616),
.Y(n_1651)
);

INVxp67_ASAP7_75t_SL g1652 ( 
.A(n_1625),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1628),
.Y(n_1653)
);

NOR2xp67_ASAP7_75t_L g1654 ( 
.A(n_1626),
.B(n_1610),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1637),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1623),
.B(n_1610),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1627),
.B(n_1610),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_L g1658 ( 
.A(n_1619),
.B(n_1629),
.C(n_1615),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1629),
.B(n_1615),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1641),
.B(n_1596),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1636),
.B(n_1598),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1636),
.B(n_1603),
.Y(n_1662)
);

AOI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1658),
.A2(n_1638),
.B(n_1619),
.C(n_1622),
.Y(n_1663)
);

AOI221x1_ASAP7_75t_L g1664 ( 
.A1(n_1651),
.A2(n_1631),
.B1(n_1632),
.B2(n_1640),
.C(n_1635),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1654),
.B(n_1636),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1659),
.A2(n_1633),
.B1(n_1639),
.B2(n_1612),
.C(n_1611),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_L g1667 ( 
.A(n_1650),
.B(n_1642),
.C(n_1582),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1656),
.Y(n_1668)
);

NOR3xp33_ASAP7_75t_L g1669 ( 
.A(n_1652),
.B(n_1612),
.C(n_1636),
.Y(n_1669)
);

O2A1O1Ixp5_ASAP7_75t_L g1670 ( 
.A1(n_1660),
.A2(n_1611),
.B(n_1584),
.C(n_1597),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1646),
.A2(n_1581),
.B1(n_1582),
.B2(n_1595),
.C(n_1599),
.Y(n_1671)
);

NOR4xp25_ASAP7_75t_L g1672 ( 
.A(n_1643),
.B(n_1595),
.C(n_1581),
.D(n_1599),
.Y(n_1672)
);

AOI21xp33_ASAP7_75t_SL g1673 ( 
.A1(n_1660),
.A2(n_1592),
.B(n_1614),
.Y(n_1673)
);

OAI21xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1661),
.A2(n_1584),
.B(n_1598),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1668),
.B(n_1643),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1667),
.A2(n_1662),
.B1(n_1649),
.B2(n_1657),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_SL g1677 ( 
.A(n_1663),
.B(n_1644),
.C(n_1661),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1669),
.B(n_1644),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1670),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1664),
.Y(n_1680)
);

OAI31xp33_ASAP7_75t_L g1681 ( 
.A1(n_1665),
.A2(n_1656),
.A3(n_1647),
.B(n_1649),
.Y(n_1681)
);

NOR2x1p5_ASAP7_75t_L g1682 ( 
.A(n_1673),
.B(n_1653),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_SL g1683 ( 
.A(n_1674),
.B(n_1655),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1666),
.B(n_1653),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1671),
.A2(n_1655),
.B1(n_1647),
.B2(n_1648),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1672),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1675),
.Y(n_1687)
);

NAND4xp25_ASAP7_75t_L g1688 ( 
.A(n_1681),
.B(n_1648),
.C(n_1645),
.D(n_1584),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1678),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1682),
.B(n_1645),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1676),
.A2(n_1594),
.B1(n_1590),
.B2(n_1593),
.C(n_1597),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1677),
.B(n_1592),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1675),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1690),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1692),
.B(n_1679),
.Y(n_1695)
);

INVxp33_ASAP7_75t_SL g1696 ( 
.A(n_1689),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1688),
.A2(n_1680),
.B1(n_1686),
.B2(n_1683),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1691),
.A2(n_1684),
.B1(n_1685),
.B2(n_1540),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1687),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1693),
.Y(n_1700)
);

OR2x6_ASAP7_75t_L g1701 ( 
.A(n_1694),
.B(n_1237),
.Y(n_1701)
);

AOI211x1_ASAP7_75t_L g1702 ( 
.A1(n_1695),
.A2(n_1604),
.B(n_1603),
.C(n_1598),
.Y(n_1702)
);

AND3x4_ASAP7_75t_L g1703 ( 
.A(n_1696),
.B(n_1557),
.C(n_1239),
.Y(n_1703)
);

NAND2x1p5_ASAP7_75t_L g1704 ( 
.A(n_1699),
.B(n_1239),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1700),
.Y(n_1705)
);

NOR4xp25_ASAP7_75t_L g1706 ( 
.A(n_1705),
.B(n_1697),
.C(n_1698),
.D(n_1590),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1702),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1701),
.B(n_1603),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1708),
.Y(n_1709)
);

OAI322xp33_ASAP7_75t_L g1710 ( 
.A1(n_1709),
.A2(n_1707),
.A3(n_1704),
.B1(n_1706),
.B2(n_1703),
.C1(n_1593),
.C2(n_1590),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1710),
.A2(n_1597),
.B1(n_1594),
.B2(n_1593),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1710),
.A2(n_1375),
.B1(n_1594),
.B2(n_1237),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1557),
.B1(n_1604),
.B2(n_1409),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1711),
.A2(n_1642),
.B1(n_1614),
.B2(n_1604),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1713),
.A2(n_1579),
.B(n_1272),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1714),
.A2(n_1539),
.B1(n_1545),
.B2(n_1561),
.Y(n_1716)
);

INVxp33_ASAP7_75t_L g1717 ( 
.A(n_1715),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1717),
.A2(n_1716),
.B(n_1539),
.Y(n_1718)
);

OAI221xp5_ASAP7_75t_R g1719 ( 
.A1(n_1718),
.A2(n_1318),
.B1(n_1561),
.B2(n_1562),
.C(n_1560),
.Y(n_1719)
);

AOI211xp5_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1318),
.B(n_1524),
.C(n_1522),
.Y(n_1720)
);


endmodule