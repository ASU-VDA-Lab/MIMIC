module fake_netlist_6_2902_n_106 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_106);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_106;

wire n_52;
wire n_91;
wire n_46;
wire n_18;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

OA21x2_ASAP7_75t_L g42 ( 
.A1(n_24),
.A2(n_0),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_0),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_30),
.Y(n_46)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_30),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2x1p5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp67_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_35),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_39),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_42),
.B1(n_43),
.B2(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_49),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_47),
.B1(n_52),
.B2(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2x1p5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

CKINVDCx11_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_47),
.B1(n_55),
.B2(n_41),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_57),
.B1(n_51),
.B2(n_52),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_63),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_51),
.B1(n_64),
.B2(n_60),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_60),
.B1(n_29),
.B2(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.C(n_38),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

OAI33xp33_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_40),
.A3(n_37),
.B1(n_36),
.B2(n_50),
.B3(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_58),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_58),
.C(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_81),
.A2(n_42),
.B(n_34),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_SL g89 ( 
.A(n_85),
.B(n_53),
.C(n_79),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_84),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_2),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_86),
.A3(n_38),
.B1(n_87),
.B2(n_3),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_91),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_89),
.B1(n_38),
.B2(n_49),
.Y(n_95)
);

OAI31xp33_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_4),
.A3(n_53),
.B(n_12),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

NAND4xp25_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_93),
.C(n_13),
.D(n_8),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_44),
.C(n_97),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_99),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

NAND4xp25_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_44),
.C(n_99),
.D(n_93),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_100),
.B(n_101),
.Y(n_106)
);


endmodule