module fake_jpeg_16254_n_81 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_81);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_81;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx2_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_16),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_11),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_13),
.B1(n_15),
.B2(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_10),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_12),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_24),
.C(n_22),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_42),
.C(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_13),
.B1(n_19),
.B2(n_21),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_42),
.B(n_14),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_9),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_46),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_49),
.B1(n_51),
.B2(n_24),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_1),
.B(n_2),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_32),
.B(n_35),
.Y(n_55)
);

AND2x6_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_1),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_52),
.B1(n_10),
.B2(n_14),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_56),
.B1(n_59),
.B2(n_5),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_58),
.B(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_39),
.B1(n_21),
.B2(n_7),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_19),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_18),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_60),
.A2(n_45),
.B1(n_48),
.B2(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_58),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_64),
.B(n_66),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_55),
.B(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_70),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_72),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_65),
.B1(n_5),
.B2(n_8),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_73),
.A2(n_24),
.B(n_2),
.C(n_8),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_2),
.B(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_77),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_76),
.Y(n_81)
);


endmodule