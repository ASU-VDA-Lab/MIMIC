module real_jpeg_18341_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_8),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_1),
.B(n_53),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_1),
.B(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_2),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_2),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_2),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_3),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_3),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_3),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_3),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_4),
.B(n_53),
.Y(n_52)
);

AND2x4_ASAP7_75t_SL g83 ( 
.A(n_4),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_5),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_5),
.A2(n_12),
.B1(n_113),
.B2(n_118),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_5),
.B(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_5),
.Y(n_186)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_6),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_7),
.B(n_151),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_9),
.Y(n_138)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_9),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_10),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_11),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_11),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_11),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_11),
.B(n_115),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_12),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_12),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_12),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_12),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_12),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_12),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_12),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_13),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_13),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_13),
.B(n_96),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g103 ( 
.A(n_13),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_13),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_13),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_13),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_14),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_14),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_15),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_15),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_15),
.B(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_15),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_15),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_15),
.B(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_16),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_16),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_18),
.Y(n_148)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_206),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_172),
.B(n_203),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_25),
.B(n_173),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_99),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_66),
.C(n_87),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_27),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.C(n_57),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_29),
.B(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_30),
.B(n_40),
.C(n_46),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_38),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_47),
.B(n_57),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_48),
.B(n_52),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_51),
.Y(n_194)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_51),
.Y(n_257)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_56),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.C(n_63),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_58),
.A2(n_61),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_58),
.Y(n_215)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_61),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_61),
.A2(n_216),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_61),
.B(n_283),
.C(n_287),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_62),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_63),
.B(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_66),
.B(n_87),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_67),
.B(n_78),
.C(n_85),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.C(n_75),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_68),
.A2(n_75),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_68),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_71),
.B(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_75),
.Y(n_180)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_76),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_81),
.Y(n_184)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_93),
.C(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_90),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_95),
.A2(n_97),
.B1(n_219),
.B2(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_97),
.B(n_219),
.C(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_142),
.B1(n_170),
.B2(n_171),
.Y(n_99)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_125),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_111),
.C(n_124),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_102),
.B(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_106),
.C(n_110),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_111),
.A2(n_112),
.B1(n_124),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_112),
.A2(n_182),
.B(n_185),
.Y(n_181)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_135),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_129),
.A2(n_130),
.B1(n_196),
.B2(n_197),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_130),
.B(n_191),
.C(n_196),
.Y(n_190)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_157),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_150),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_151),
.Y(n_253)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_151),
.Y(n_281)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_155),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_199),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_176),
.B(n_200),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_190),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_181),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_179),
.B(n_237),
.C(n_241),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_191),
.B(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_SL g271 ( 
.A(n_192),
.B(n_195),
.Y(n_271)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_192),
.A2(n_278),
.B1(n_279),
.B2(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_228),
.B(n_328),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_226),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_SL g329 ( 
.A(n_209),
.B(n_226),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.C(n_224),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_210),
.B(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_212),
.B(n_224),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.C(n_222),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_213),
.B(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_218),
.B(n_223),
.Y(n_320)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_219),
.Y(n_267)
);

XOR2x1_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_323),
.B(n_327),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_309),
.B(n_322),
.Y(n_231)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_274),
.B(n_308),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_262),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_234),
.B(n_262),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_245),
.C(n_254),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_235),
.B(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_245),
.A2(n_246),
.B1(n_254),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_252),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_247),
.B(n_252),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_254),
.Y(n_305)
);

AO22x1_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_254)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_255),
.Y(n_260)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_258),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_260),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_268),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_265),
.C(n_268),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_271),
.C(n_272),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_302),
.B(n_307),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_290),
.B(n_301),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_282),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_297),
.B(n_300),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_295),
.Y(n_300)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_306),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_321),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_SL g322 ( 
.A(n_310),
.B(n_321),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_318),
.B2(n_319),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_317),
.C(n_318),
.Y(n_326)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_326),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);


endmodule