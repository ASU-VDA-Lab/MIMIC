module fake_jpeg_31336_n_365 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_365);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_365;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_40),
.B(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_43),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_23),
.B(n_21),
.CON(n_43),
.SN(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_16),
.C(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_17),
.B(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_65),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_13),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_13),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_20),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_29),
.B1(n_31),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_76),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_29),
.B1(n_31),
.B2(n_30),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_97),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_38),
.B1(n_19),
.B2(n_20),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_39),
.B1(n_34),
.B2(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_92),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_35),
.B1(n_63),
.B2(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_82),
.A2(n_93),
.B1(n_101),
.B2(n_56),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_34),
.B1(n_36),
.B2(n_22),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_36),
.B1(n_28),
.B2(n_32),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_18),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_35),
.B1(n_22),
.B2(n_28),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_96),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_36),
.B1(n_25),
.B2(n_32),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_94),
.A2(n_107),
.B1(n_106),
.B2(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_26),
.B1(n_25),
.B2(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_26),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_46),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_2),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_37),
.B1(n_16),
.B2(n_11),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_50),
.A2(n_37),
.B1(n_16),
.B2(n_4),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_41),
.A2(n_37),
.B1(n_18),
.B2(n_4),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_54),
.B1(n_58),
.B2(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_150),
.B1(n_74),
.B2(n_73),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_65),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_60),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_124),
.Y(n_159)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_88),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_55),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_130),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_51),
.B1(n_37),
.B2(n_18),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_140),
.Y(n_152)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_37),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_76),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_136),
.Y(n_171)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

OR2x2_ASAP7_75t_SL g133 ( 
.A(n_71),
.B(n_58),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_R g178 ( 
.A(n_133),
.B(n_149),
.Y(n_178)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_147),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_55),
.B(n_44),
.C(n_58),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_44),
.B(n_37),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_107),
.C(n_67),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx5_ASAP7_75t_SL g166 ( 
.A(n_142),
.Y(n_166)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_72),
.B(n_18),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_78),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_89),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_81),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_153),
.A2(n_176),
.B1(n_177),
.B2(n_120),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_71),
.B(n_72),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_184),
.B(n_137),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_106),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_160),
.B(n_126),
.C(n_3),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_75),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_111),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_67),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_167),
.A2(n_168),
.B(n_169),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_96),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_95),
.B(n_89),
.C(n_90),
.Y(n_170)
);

AO22x1_ASAP7_75t_L g210 ( 
.A1(n_170),
.A2(n_174),
.B1(n_138),
.B2(n_135),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_139),
.A2(n_100),
.B1(n_109),
.B2(n_105),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_144),
.A2(n_105),
.B1(n_56),
.B2(n_103),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_125),
.B(n_103),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_125),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_134),
.A2(n_108),
.B(n_81),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_143),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_103),
.B1(n_81),
.B2(n_18),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_128),
.B1(n_133),
.B2(n_121),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_197),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_188),
.A2(n_191),
.B1(n_193),
.B2(n_195),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_189),
.B(n_192),
.Y(n_232)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_111),
.B1(n_121),
.B2(n_134),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_152),
.A2(n_111),
.B1(n_123),
.B2(n_147),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_194),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_152),
.A2(n_114),
.B1(n_122),
.B2(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_114),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_202),
.Y(n_245)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_129),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_161),
.B(n_113),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_112),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_208),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_159),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_112),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_136),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_209),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_216),
.B(n_174),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_211),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_212),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_155),
.B(n_148),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_222),
.C(n_185),
.Y(n_229)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_214),
.Y(n_246)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

INVxp33_ASAP7_75t_SL g247 ( 
.A(n_215),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_153),
.A2(n_178),
.B1(n_170),
.B2(n_186),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_178),
.B1(n_182),
.B2(n_184),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_182),
.A2(n_142),
.B1(n_126),
.B2(n_18),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_228),
.B1(n_234),
.B2(n_188),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_170),
.B(n_167),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_225),
.B(n_229),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_167),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_235),
.C(n_250),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_169),
.B1(n_165),
.B2(n_176),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_185),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_165),
.B(n_185),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_245),
.Y(n_262)
);

AOI22x1_ASAP7_75t_L g243 ( 
.A1(n_210),
.A2(n_169),
.B1(n_177),
.B2(n_166),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_214),
.B(n_210),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_209),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_197),
.B(n_217),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_191),
.A2(n_162),
.B(n_157),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_253),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_255),
.A2(n_260),
.B1(n_268),
.B2(n_273),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_194),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_261),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_247),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_258),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_223),
.A2(n_228),
.B1(n_246),
.B2(n_245),
.Y(n_260)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_206),
.C(n_211),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_262),
.A2(n_239),
.B(n_230),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_187),
.Y(n_263)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_226),
.C(n_235),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_266),
.C(n_270),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_208),
.B1(n_190),
.B2(n_196),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_274),
.B1(n_278),
.B2(n_258),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_198),
.C(n_222),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_193),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_269),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_195),
.B1(n_219),
.B2(n_215),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_240),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_201),
.C(n_199),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_241),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_229),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_204),
.B1(n_181),
.B2(n_166),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_230),
.A2(n_164),
.B1(n_216),
.B2(n_175),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_276),
.Y(n_298)
);

BUFx12f_ASAP7_75t_SL g277 ( 
.A(n_225),
.Y(n_277)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_239),
.A2(n_166),
.B1(n_164),
.B2(n_175),
.Y(n_278)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_282),
.A2(n_293),
.B1(n_254),
.B2(n_260),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_283),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_242),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_294),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_285),
.B(n_292),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_264),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_297),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_244),
.B(n_236),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_290),
.A2(n_172),
.B(n_179),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_243),
.B1(n_253),
.B2(n_249),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_276),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_254),
.A2(n_243),
.B1(n_233),
.B2(n_241),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_278),
.B1(n_272),
.B2(n_273),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_242),
.C(n_227),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_281),
.C(n_285),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_252),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_300),
.A2(n_307),
.B1(n_311),
.B2(n_286),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_270),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_291),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_304),
.A2(n_316),
.B1(n_287),
.B2(n_280),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_259),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_312),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_255),
.B1(n_262),
.B2(n_268),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_310),
.C(n_292),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_266),
.C(n_227),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_282),
.A2(n_252),
.B1(n_248),
.B2(n_216),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_296),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_248),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_284),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_279),
.B(n_294),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_286),
.A2(n_172),
.B1(n_179),
.B2(n_156),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_326),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_299),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_324),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_319),
.A2(n_321),
.B1(n_316),
.B2(n_315),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_287),
.B1(n_283),
.B2(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_300),
.B1(n_295),
.B2(n_311),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_327),
.C(n_328),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_325),
.A2(n_317),
.B(n_321),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_291),
.C(n_298),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_312),
.C(n_305),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_306),
.C(n_313),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_330),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_301),
.A2(n_298),
.B1(n_179),
.B2(n_156),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_333),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_325),
.A2(n_314),
.B(n_306),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_334),
.A2(n_340),
.B(n_319),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_303),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_339),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_156),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_4),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_329),
.A2(n_2),
.B(n_3),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_348),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_328),
.B(n_322),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_343),
.A2(n_337),
.B(n_338),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_341),
.B(n_322),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_345),
.Y(n_352)
);

XNOR2x1_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_2),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_347),
.B(n_349),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_4),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_5),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_350),
.A2(n_334),
.B(n_340),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_351),
.B(n_350),
.C(n_344),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_332),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_346),
.A2(n_332),
.B(n_6),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_354),
.B(n_5),
.Y(n_358)
);

MAJx2_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_359),
.C(n_360),
.Y(n_361)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_358),
.A2(n_356),
.B(n_355),
.C(n_9),
.Y(n_362)
);

AOI322xp5_ASAP7_75t_L g360 ( 
.A1(n_352),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_360)
);

OAI321xp33_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_361),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_8),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_8),
.Y(n_365)
);


endmodule