module fake_jpeg_7090_n_184 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_32),
.B(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_18),
.B(n_16),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_33),
.A2(n_41),
.B(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_21),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_3),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_22),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_3),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_50),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_24),
.B(n_20),
.C(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_48),
.B(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_52),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_29),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_57),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_24),
.C(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_63),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_30),
.B1(n_15),
.B2(n_22),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_19),
.B1(n_17),
.B2(n_7),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_22),
.B1(n_30),
.B2(n_15),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_69),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_38),
.B(n_23),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_11),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_15),
.B(n_23),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_98),
.B1(n_99),
.B2(n_102),
.Y(n_107)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_21),
.A3(n_19),
.B1(n_17),
.B2(n_8),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_12),
.C(n_13),
.Y(n_123)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_48),
.Y(n_117)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_96),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_62),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_53),
.B1(n_67),
.B2(n_71),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_55),
.B(n_61),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_112),
.B(n_118),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_75),
.B(n_74),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_119),
.Y(n_128)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_73),
.B1(n_47),
.B2(n_71),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_122),
.B1(n_89),
.B2(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_120),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_57),
.B(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_56),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_91),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_63),
.B1(n_62),
.B2(n_67),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_126),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_125),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_85),
.A2(n_91),
.B1(n_98),
.B2(n_99),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_132),
.C(n_141),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_111),
.C(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_139),
.Y(n_153)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_104),
.B(n_84),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_104),
.C(n_84),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_83),
.C(n_103),
.Y(n_155)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_109),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_150),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_126),
.B1(n_107),
.B2(n_120),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_112),
.B(n_113),
.C(n_117),
.D(n_107),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_133),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_123),
.B1(n_105),
.B2(n_89),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_154),
.B(n_130),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_151),
.C(n_140),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_137),
.A2(n_83),
.B1(n_72),
.B2(n_86),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_162),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_133),
.B1(n_137),
.B2(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_161),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_140),
.Y(n_161)
);

AO221x1_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_139),
.B1(n_142),
.B2(n_90),
.C(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_128),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

BUFx4f_ASAP7_75t_SL g170 ( 
.A(n_159),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_170),
.B(n_156),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_174),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_147),
.A3(n_165),
.B1(n_148),
.B2(n_160),
.C1(n_164),
.C2(n_157),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_165),
.B1(n_152),
.B2(n_131),
.Y(n_174)
);

BUFx12f_ASAP7_75t_SL g179 ( 
.A(n_175),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_167),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_142),
.B(n_59),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_170),
.A3(n_176),
.B1(n_174),
.B2(n_167),
.C1(n_149),
.C2(n_139),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_178),
.C(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);


endmodule