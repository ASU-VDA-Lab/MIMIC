module fake_jpeg_8572_n_269 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_29),
.B1(n_18),
.B2(n_30),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_47),
.B(n_25),
.Y(n_80)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_54),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_29),
.B1(n_18),
.B2(n_30),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_29),
.B1(n_22),
.B2(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_53),
.B1(n_60),
.B2(n_27),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_28),
.B(n_22),
.C(n_20),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_55),
.B(n_59),
.C(n_45),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_17),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_28),
.B(n_25),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_22),
.B(n_20),
.C(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_25),
.B1(n_17),
.B2(n_26),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_59),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_76),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_63),
.B1(n_77),
.B2(n_86),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_32),
.B1(n_31),
.B2(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_84),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_41),
.B1(n_40),
.B2(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_71),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_74),
.Y(n_91)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_36),
.C(n_38),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_48),
.C(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_32),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_42),
.A2(n_25),
.B1(n_31),
.B2(n_27),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_80),
.B(n_83),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_2),
.B(n_3),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_27),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_48),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_101),
.B(n_80),
.Y(n_129)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_82),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_54),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_98),
.C(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_105),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_69),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_68),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_46),
.B1(n_56),
.B2(n_50),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_79),
.B1(n_77),
.B2(n_56),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_74),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_38),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_2),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_128),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_75),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_125),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_76),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_132),
.B(n_135),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_138),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_64),
.Y(n_133)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

NOR2xp67_ASAP7_75t_SL g134 ( 
.A(n_89),
.B(n_70),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_111),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_3),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_84),
.C(n_33),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_102),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_93),
.B(n_56),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_112),
.B1(n_79),
.B2(n_21),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_50),
.B1(n_79),
.B2(n_38),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_141),
.A2(n_109),
.B1(n_106),
.B2(n_96),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_3),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_142),
.A2(n_90),
.B(n_102),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_143),
.A2(n_169),
.B1(n_135),
.B2(n_21),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_142),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_165),
.B(n_142),
.Y(n_187)
);

OAI21x1_ASAP7_75t_R g149 ( 
.A1(n_122),
.A2(n_110),
.B(n_112),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_155),
.B(n_156),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_164),
.C(n_166),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_90),
.B(n_105),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_100),
.B(n_114),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_130),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_99),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_164),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_99),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_141),
.B1(n_132),
.B2(n_127),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_38),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_52),
.B1(n_33),
.B2(n_21),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_172),
.B(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_175),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_187),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_136),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_185),
.C(n_189),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_181),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_191),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_115),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_170),
.B1(n_165),
.B2(n_155),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_153),
.B1(n_33),
.B2(n_7),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_124),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_146),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_161),
.C(n_144),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_144),
.C(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_199),
.C(n_209),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_143),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_124),
.B1(n_152),
.B2(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_207),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_145),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_208),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_124),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_157),
.C(n_162),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_171),
.B1(n_188),
.B2(n_7),
.Y(n_227)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_212),
.B(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_153),
.C(n_6),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_186),
.C(n_190),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_187),
.B(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

BUFx12_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_220),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_221),
.B(n_222),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_192),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_225),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_227),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_173),
.B(n_171),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_206),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_194),
.C(n_198),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_202),
.B(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_217),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_240),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_194),
.C(n_209),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.C(n_226),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_205),
.C(n_189),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_210),
.B(n_201),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_224),
.B1(n_220),
.B2(n_221),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_232),
.B1(n_233),
.B2(n_240),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_245),
.C(n_246),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_4),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_215),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_230),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_215),
.C(n_6),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_4),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_244),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_254),
.B(n_256),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_243),
.B(n_238),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_246),
.C(n_234),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_260),
.B(n_8),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_259),
.A3(n_255),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_4),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_14),
.C(n_7),
.Y(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_8),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

AOI321xp33_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_264),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C(n_9),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_266),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_268),
.Y(n_269)
);


endmodule