module fake_jpeg_4349_n_150 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_150);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_4),
.B(n_11),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_12),
.B(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_20),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_34),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_20),
.B(n_17),
.C(n_24),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_42),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_21),
.B1(n_22),
.B2(n_12),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_26),
.A2(n_21),
.B1(n_22),
.B2(n_12),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_30),
.B(n_25),
.C(n_29),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_52),
.Y(n_79)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

HAxp5_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_32),
.CON(n_53),
.SN(n_53)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_32),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_31),
.B(n_34),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_32),
.B1(n_17),
.B2(n_25),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_64),
.B1(n_44),
.B2(n_41),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_18),
.B1(n_21),
.B2(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_39),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_18),
.B1(n_28),
.B2(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_46),
.B1(n_28),
.B2(n_33),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_44),
.B1(n_52),
.B2(n_41),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_94),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_48),
.C(n_59),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_59),
.C(n_48),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_73),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_103),
.Y(n_115)
);

OAI221xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_72),
.B1(n_68),
.B2(n_74),
.C(n_66),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_100),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_76),
.C(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_104),
.Y(n_116)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_53),
.B(n_75),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_100),
.B(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_83),
.B1(n_93),
.B2(n_87),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_114),
.B1(n_121),
.B2(n_46),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_71),
.B1(n_78),
.B2(n_46),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_120),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_116),
.B(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_102),
.B1(n_110),
.B2(n_101),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_111),
.B1(n_114),
.B2(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_35),
.B(n_69),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_127),
.B(n_14),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_112),
.C(n_113),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_128),
.C(n_129),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_82),
.C(n_32),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_32),
.C(n_29),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_27),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_130),
.B(n_27),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_134),
.B(n_137),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_17),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_126),
.B(n_124),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_135),
.A2(n_13),
.B(n_2),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_0),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_141),
.B(n_140),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_15),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_132),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_23),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_1),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_2),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_7),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_146)
);

OAI21x1_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_144),
.B(n_10),
.Y(n_147)
);

AOI21x1_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_9),
.B(n_11),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_16),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_16),
.Y(n_150)
);


endmodule