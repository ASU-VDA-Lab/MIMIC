module fake_jpeg_3105_n_96 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_46),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_30),
.B1(n_35),
.B2(n_29),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_35),
.B1(n_27),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_40),
.B1(n_31),
.B2(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_56),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_31),
.B1(n_34),
.B2(n_2),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_34),
.B1(n_2),
.B2(n_3),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_0),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_67),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_1),
.B(n_3),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_5),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_73),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_15),
.B1(n_23),
.B2(n_22),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_17),
.B1(n_21),
.B2(n_9),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_6),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_64),
.B(n_16),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_78),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_11),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_74),
.B(n_26),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_72),
.B1(n_10),
.B2(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_84),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_87),
.B1(n_80),
.B2(n_83),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_83),
.B1(n_81),
.B2(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_8),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_8),
.Y(n_96)
);


endmodule