module fake_ariane_411_n_923 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_923);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_923;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_885;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_731;
wire n_336;
wire n_665;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_839;
wire n_770;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_238;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_260;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_847;
wire n_772;
wire n_741;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_856;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_767;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_95),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_80),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_57),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_75),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_25),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_65),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_53),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_2),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_157),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_26),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_29),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_107),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_154),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_160),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_40),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_97),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_105),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_69),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_126),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_12),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_88),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_60),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_79),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_35),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_46),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_18),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_55),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_61),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_21),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_15),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_58),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_101),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_164),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_30),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_140),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_182),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_122),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_92),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_39),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_103),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_24),
.Y(n_242)
);

BUFx4f_ASAP7_75t_SL g243 ( 
.A(n_84),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_36),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_13),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_82),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_26),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_110),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_121),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_85),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_135),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_23),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_22),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_42),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_81),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_176),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_49),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_145),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_33),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_54),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_4),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_169),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_4),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_128),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_3),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_38),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_64),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_68),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_151),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_165),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_170),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_52),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_168),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_134),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_21),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_124),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_115),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_159),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_138),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_63),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_137),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_56),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_172),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_207),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_204),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_209),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_212),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

BUFx2_ASAP7_75t_SL g290 ( 
.A(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_252),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_276),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_255),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_211),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_255),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_232),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_0),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_206),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_190),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_0),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_190),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_224),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_224),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_215),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_190),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_200),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_196),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_240),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_196),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_196),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_196),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_214),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_214),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_214),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_214),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_278),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_191),
.B(n_1),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_278),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_257),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_248),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_253),
.B(n_1),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_233),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_262),
.B(n_2),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_198),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_264),
.B(n_3),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_203),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_284),
.B(n_5),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_227),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_189),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_228),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_192),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_199),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_210),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_243),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_193),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_283),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_233),
.B(n_5),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_195),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_282),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_217),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_195),
.B(n_6),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_218),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_219),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_303),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_289),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_295),
.Y(n_354)
);

NAND2xp33_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_251),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_309),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_221),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_220),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_219),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_350),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_229),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_334),
.Y(n_366)
);

OA21x2_ASAP7_75t_L g367 ( 
.A1(n_350),
.A2(n_237),
.B(n_235),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_331),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_340),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_335),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_292),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_313),
.Y(n_373)
);

AND2x6_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_230),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_296),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_304),
.B(n_261),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_329),
.B(n_239),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_R g379 ( 
.A(n_341),
.B(n_194),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_315),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_317),
.Y(n_382)
);

NAND2xp33_ASAP7_75t_L g383 ( 
.A(n_298),
.B(n_251),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_326),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_319),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_L g386 ( 
.A1(n_298),
.A2(n_249),
.B1(n_230),
.B2(n_241),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_343),
.Y(n_388)
);

CKINVDCx6p67_ASAP7_75t_R g389 ( 
.A(n_290),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_R g390 ( 
.A(n_336),
.B(n_197),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_325),
.B(n_244),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_346),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_320),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_307),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_290),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_336),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_345),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_286),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_301),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_338),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_338),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_342),
.B(n_250),
.Y(n_407)
);

NOR2x1p5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_285),
.Y(n_408)
);

OR2x6_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_337),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_353),
.Y(n_410)
);

AND2x2_ASAP7_75t_SL g411 ( 
.A(n_355),
.B(n_241),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_342),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_363),
.B1(n_367),
.B2(n_386),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_377),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_249),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_304),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_393),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_311),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_406),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_359),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_395),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_354),
.B(n_297),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_285),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_287),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_393),
.Y(n_428)
);

AND2x6_ASAP7_75t_SL g429 ( 
.A(n_407),
.B(n_259),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_388),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_366),
.B(n_306),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_287),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_401),
.A2(n_344),
.B1(n_288),
.B2(n_294),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_368),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_360),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_366),
.B(n_306),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_405),
.B(n_288),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_365),
.B(n_310),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_374),
.A2(n_305),
.B1(n_330),
.B2(n_328),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_383),
.A2(n_294),
.B1(n_322),
.B2(n_310),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_370),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_361),
.B(n_302),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_322),
.Y(n_447)
);

NAND2x1p5_ASAP7_75t_L g448 ( 
.A(n_369),
.B(n_332),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_401),
.B(n_251),
.Y(n_449)
);

AND2x2_ASAP7_75t_SL g450 ( 
.A(n_355),
.B(n_383),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_401),
.B(n_251),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_403),
.B(n_327),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_389),
.B(n_327),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_360),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_403),
.B(n_300),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_403),
.B(n_263),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_392),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_379),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_364),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_403),
.B(n_265),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_379),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_370),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_352),
.B(n_268),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_372),
.B(n_274),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_399),
.B(n_201),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_382),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_385),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_385),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_396),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_374),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_374),
.B(n_202),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_358),
.A2(n_299),
.B1(n_281),
.B2(n_280),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_390),
.B(n_205),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_430),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_351),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_391),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_363),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_363),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_414),
.B(n_442),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_432),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_445),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_428),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_414),
.B(n_363),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_363),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_451),
.B(n_367),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_416),
.B(n_390),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_418),
.B(n_357),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_415),
.A2(n_260),
.B1(n_213),
.B2(n_216),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_L g494 ( 
.A(n_415),
.B(n_208),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_416),
.B(n_378),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_462),
.B(n_456),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_468),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_432),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_381),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_428),
.A2(n_367),
.B(n_223),
.Y(n_500)
);

O2A1O1Ixp33_ASAP7_75t_L g501 ( 
.A1(n_412),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_433),
.B(n_373),
.Y(n_502)
);

A2O1A1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_457),
.A2(n_267),
.B(n_225),
.C(n_226),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_467),
.B(n_415),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_415),
.B(n_222),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_413),
.A2(n_384),
.B1(n_375),
.B2(n_371),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_413),
.A2(n_375),
.B1(n_371),
.B2(n_279),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_446),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_435),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_409),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_415),
.B(n_231),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_417),
.B(n_234),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_417),
.B(n_236),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_425),
.B(n_7),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_440),
.B(n_238),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_471),
.B(n_247),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_410),
.B(n_256),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_446),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_451),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_438),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_419),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_422),
.B(n_258),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_466),
.A2(n_277),
.B1(n_275),
.B2(n_273),
.Y(n_526)
);

NOR2x1p5_ASAP7_75t_L g527 ( 
.A(n_424),
.B(n_270),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_466),
.A2(n_272),
.B1(n_271),
.B2(n_10),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_437),
.B(n_8),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_454),
.B(n_186),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_471),
.B(n_9),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_444),
.B(n_9),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_459),
.B(n_10),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_431),
.B(n_11),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_431),
.B(n_11),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_411),
.B(n_12),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_409),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_SL g538 ( 
.A(n_434),
.B(n_13),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_423),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_466),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_427),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_441),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_411),
.B(n_14),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_458),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_421),
.B(n_16),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_460),
.Y(n_546)
);

AOI22x1_ASAP7_75t_L g547 ( 
.A1(n_472),
.A2(n_477),
.B1(n_439),
.B2(n_455),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_522),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_522),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_483),
.A2(n_491),
.B1(n_480),
.B2(n_482),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_506),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_544),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_524),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_478),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_480),
.B(n_421),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_517),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_489),
.B(n_450),
.Y(n_559)
);

NOR3xp33_ASAP7_75t_SL g560 ( 
.A(n_538),
.B(n_436),
.C(n_475),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_521),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_484),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_492),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_489),
.B(n_450),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_485),
.Y(n_565)
);

AOI21x1_ASAP7_75t_L g566 ( 
.A1(n_500),
.A2(n_461),
.B(n_457),
.Y(n_566)
);

BUFx4f_ASAP7_75t_L g567 ( 
.A(n_492),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_486),
.B(n_464),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_479),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_522),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_508),
.A2(n_466),
.B1(n_443),
.B2(n_472),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_539),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_541),
.B(n_464),
.Y(n_574)
);

CKINVDCx8_ASAP7_75t_R g575 ( 
.A(n_511),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_499),
.B(n_461),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_537),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_487),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_542),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_481),
.B(n_426),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_515),
.B(n_448),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_R g582 ( 
.A(n_509),
.B(n_418),
.Y(n_582)
);

AND2x2_ASAP7_75t_SL g583 ( 
.A(n_508),
.B(n_528),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_481),
.B(n_443),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_498),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_482),
.B(n_466),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_510),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_520),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_545),
.B(n_476),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_R g590 ( 
.A(n_494),
.B(n_429),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_496),
.B(n_476),
.Y(n_591)
);

BUFx4f_ASAP7_75t_L g592 ( 
.A(n_490),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_545),
.B(n_448),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_536),
.Y(n_594)
);

BUFx12f_ASAP7_75t_L g595 ( 
.A(n_527),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_SL g596 ( 
.A(n_543),
.B(n_408),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_523),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_529),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_490),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_487),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_497),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_507),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_495),
.B(n_468),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_546),
.Y(n_604)
);

BUFx4f_ASAP7_75t_L g605 ( 
.A(n_530),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_504),
.B(n_474),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_555),
.B(n_507),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_566),
.A2(n_547),
.B(n_488),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_583),
.A2(n_540),
.B1(n_528),
.B2(n_532),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_559),
.A2(n_535),
.B(n_534),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_564),
.A2(n_535),
.B(n_534),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_550),
.B(n_439),
.Y(n_612)
);

OA21x2_ASAP7_75t_L g613 ( 
.A1(n_606),
.A2(n_566),
.B(n_586),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_580),
.B(n_455),
.Y(n_614)
);

OAI21x1_ASAP7_75t_L g615 ( 
.A1(n_551),
.A2(n_477),
.B(n_470),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_551),
.A2(n_473),
.B(n_470),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_576),
.A2(n_503),
.B(n_540),
.Y(n_617)
);

AO32x2_ASAP7_75t_L g618 ( 
.A1(n_583),
.A2(n_501),
.A3(n_449),
.B1(n_452),
.B2(n_533),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_553),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_502),
.Y(n_620)
);

AO31x2_ASAP7_75t_L g621 ( 
.A1(n_584),
.A2(n_473),
.A3(n_512),
.B(n_505),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_573),
.Y(n_622)
);

AOI211x1_ASAP7_75t_L g623 ( 
.A1(n_574),
.A2(n_531),
.B(n_525),
.C(n_519),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_556),
.A2(n_514),
.B(n_513),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_602),
.B(n_526),
.Y(n_625)
);

AOI21x1_ASAP7_75t_L g626 ( 
.A1(n_589),
.A2(n_593),
.B(n_603),
.Y(n_626)
);

AOI221x1_ASAP7_75t_L g627 ( 
.A1(n_596),
.A2(n_469),
.B1(n_465),
.B2(n_449),
.C(n_452),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_556),
.A2(n_516),
.B(n_518),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_594),
.B(n_526),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_557),
.Y(n_630)
);

OAI21x1_ASAP7_75t_SL g631 ( 
.A1(n_578),
.A2(n_493),
.B(n_452),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_572),
.A2(n_560),
.B1(n_598),
.B2(n_602),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_557),
.A2(n_469),
.B(n_465),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_561),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_591),
.B(n_449),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_605),
.A2(n_469),
.B(n_465),
.Y(n_636)
);

OAI21xp33_ASAP7_75t_SL g637 ( 
.A1(n_578),
.A2(n_17),
.B(n_18),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_594),
.B(n_465),
.Y(n_638)
);

OAI21x1_ASAP7_75t_SL g639 ( 
.A1(n_578),
.A2(n_449),
.B(n_452),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_587),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_597),
.B(n_469),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_561),
.A2(n_452),
.B(n_449),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_597),
.A2(n_17),
.B(n_19),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_548),
.A2(n_108),
.B(n_184),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_562),
.B(n_19),
.Y(n_645)
);

OAI21x1_ASAP7_75t_L g646 ( 
.A1(n_548),
.A2(n_106),
.B(n_183),
.Y(n_646)
);

AOI21x1_ASAP7_75t_L g647 ( 
.A1(n_562),
.A2(n_104),
.B(n_181),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_585),
.Y(n_648)
);

NOR2x1_ASAP7_75t_L g649 ( 
.A(n_554),
.B(n_185),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_548),
.A2(n_102),
.B(n_177),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g651 ( 
.A1(n_585),
.A2(n_100),
.B(n_174),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_569),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_600),
.A2(n_109),
.B(n_173),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_610),
.A2(n_605),
.B(n_596),
.C(n_581),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_608),
.A2(n_600),
.B(n_601),
.Y(n_655)
);

A2O1A1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_610),
.A2(n_605),
.B(n_581),
.C(n_567),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_609),
.A2(n_632),
.B1(n_625),
.B2(n_607),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_628),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_634),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_630),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_648),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_624),
.A2(n_600),
.B(n_601),
.Y(n_662)
);

BUFx8_ASAP7_75t_L g663 ( 
.A(n_618),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_633),
.A2(n_599),
.B(n_592),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_626),
.A2(n_599),
.B(n_592),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_615),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_638),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_611),
.A2(n_592),
.B(n_567),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_609),
.A2(n_590),
.B1(n_604),
.B2(n_567),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_612),
.A2(n_571),
.B(n_549),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_612),
.A2(n_599),
.B(n_571),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_620),
.B(n_565),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_651),
.A2(n_599),
.B(n_571),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_638),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_632),
.B(n_579),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_611),
.A2(n_549),
.B(n_570),
.Y(n_676)
);

OAI21x1_ASAP7_75t_SL g677 ( 
.A1(n_631),
.A2(n_549),
.B(n_570),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_613),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_616),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_617),
.A2(n_604),
.B(n_563),
.C(n_579),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_617),
.A2(n_570),
.B(n_563),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_640),
.B(n_599),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_645),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_642),
.A2(n_571),
.B(n_558),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_653),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_619),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_622),
.B(n_565),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_629),
.Y(n_688)
);

NAND2x1p5_ASAP7_75t_L g689 ( 
.A(n_649),
.B(n_571),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_641),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_629),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_645),
.Y(n_692)
);

OAI22x1_ASAP7_75t_L g693 ( 
.A1(n_652),
.A2(n_588),
.B1(n_595),
.B2(n_575),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_644),
.Y(n_694)
);

OAI211xp5_ASAP7_75t_L g695 ( 
.A1(n_643),
.A2(n_554),
.B(n_552),
.C(n_582),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_641),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_686),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_687),
.B(n_577),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_577),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_686),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_657),
.A2(n_643),
.B1(n_614),
.B2(n_595),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_659),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_675),
.B(n_552),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_669),
.A2(n_635),
.B1(n_637),
.B2(n_614),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_659),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_657),
.A2(n_623),
.B1(n_575),
.B2(n_636),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_670),
.A2(n_627),
.B(n_613),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_660),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_680),
.A2(n_650),
.B(n_646),
.C(n_618),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_667),
.Y(n_710)
);

AOI221xp5_ASAP7_75t_L g711 ( 
.A1(n_693),
.A2(n_618),
.B1(n_639),
.B2(n_25),
.C(n_27),
.Y(n_711)
);

NOR2x1_ASAP7_75t_SL g712 ( 
.A(n_695),
.B(n_647),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_R g713 ( 
.A(n_671),
.B(n_621),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_654),
.A2(n_621),
.B(n_24),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_668),
.A2(n_621),
.B(n_27),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_660),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_682),
.B(n_20),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_676),
.A2(n_28),
.B(n_29),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

AO21x2_ASAP7_75t_L g720 ( 
.A1(n_662),
.A2(n_679),
.B(n_666),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_672),
.B(n_28),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_661),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_663),
.A2(n_693),
.B1(n_688),
.B2(n_683),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_687),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_683),
.B(n_30),
.C(n_31),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_682),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_682),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_691),
.Y(n_728)
);

O2A1O1Ixp33_ASAP7_75t_SL g729 ( 
.A1(n_656),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_671),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_663),
.A2(n_37),
.B1(n_41),
.B2(n_43),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_674),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_692),
.B(n_179),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_692),
.B(n_44),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_689),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_696),
.Y(n_736)
);

OAI21x1_ASAP7_75t_L g737 ( 
.A1(n_673),
.A2(n_47),
.B(n_48),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_696),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_689),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_SL g740 ( 
.A1(n_663),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_740)
);

NOR2x1_ASAP7_75t_SL g741 ( 
.A(n_690),
.B(n_62),
.Y(n_741)
);

AO21x2_ASAP7_75t_L g742 ( 
.A1(n_662),
.A2(n_66),
.B(n_67),
.Y(n_742)
);

NAND2x1p5_ASAP7_75t_L g743 ( 
.A(n_664),
.B(n_70),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_681),
.B(n_71),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_685),
.A2(n_171),
.B(n_73),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_724),
.B(n_698),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_719),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_710),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_710),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_701),
.A2(n_663),
.B1(n_690),
.B2(n_689),
.Y(n_750)
);

OAI211xp5_ASAP7_75t_SL g751 ( 
.A1(n_721),
.A2(n_658),
.B(n_678),
.C(n_679),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_701),
.A2(n_740),
.B1(n_731),
.B2(n_714),
.Y(n_752)
);

OAI211xp5_ASAP7_75t_L g753 ( 
.A1(n_718),
.A2(n_658),
.B(n_678),
.C(n_694),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_728),
.Y(n_754)
);

OAI31xp33_ASAP7_75t_L g755 ( 
.A1(n_706),
.A2(n_678),
.A3(n_658),
.B(n_666),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_722),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_732),
.B(n_700),
.Y(n_757)
);

O2A1O1Ixp5_ASAP7_75t_L g758 ( 
.A1(n_733),
.A2(n_677),
.B(n_684),
.C(n_694),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_731),
.A2(n_665),
.B1(n_694),
.B2(n_685),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_740),
.A2(n_665),
.B1(n_694),
.B2(n_685),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_711),
.A2(n_673),
.B(n_684),
.C(n_664),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_703),
.A2(n_694),
.B1(n_685),
.B2(n_677),
.Y(n_762)
);

NOR2x1_ASAP7_75t_L g763 ( 
.A(n_725),
.B(n_703),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_709),
.A2(n_685),
.B(n_655),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_717),
.A2(n_655),
.B1(n_74),
.B2(n_76),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_717),
.Y(n_766)
);

OA21x2_ASAP7_75t_L g767 ( 
.A1(n_707),
.A2(n_72),
.B(n_77),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_726),
.B(n_78),
.Y(n_768)
);

AOI21x1_ASAP7_75t_L g769 ( 
.A1(n_733),
.A2(n_83),
.B(n_86),
.Y(n_769)
);

AOI221xp5_ASAP7_75t_L g770 ( 
.A1(n_715),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.C(n_91),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_699),
.Y(n_771)
);

OAI21x1_ASAP7_75t_SL g772 ( 
.A1(n_712),
.A2(n_93),
.B(n_94),
.Y(n_772)
);

AOI221xp5_ASAP7_75t_L g773 ( 
.A1(n_729),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.C(n_111),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_702),
.B(n_112),
.Y(n_774)
);

OAI221xp5_ASAP7_75t_L g775 ( 
.A1(n_704),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.C(n_117),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_723),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_SL g777 ( 
.A1(n_723),
.A2(n_123),
.B(n_125),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_726),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_705),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_697),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_738),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_726),
.B(n_129),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_744),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_747),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_747),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_749),
.B(n_738),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_781),
.Y(n_787)
);

NOR2x1_ASAP7_75t_L g788 ( 
.A(n_751),
.B(n_739),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_756),
.B(n_779),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_756),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_780),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_757),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_748),
.B(n_730),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_746),
.B(n_730),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_762),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_778),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_767),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_778),
.B(n_730),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_778),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_763),
.B(n_736),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_778),
.B(n_730),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_758),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_767),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_766),
.B(n_720),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_766),
.B(n_720),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_767),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_752),
.A2(n_727),
.B1(n_726),
.B2(n_716),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_771),
.B(n_742),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_771),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_761),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_774),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_785),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_810),
.A2(n_752),
.B1(n_777),
.B2(n_776),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_800),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_787),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_800),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_785),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_794),
.B(n_755),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_785),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_794),
.B(n_764),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_784),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_784),
.Y(n_822)
);

NOR4xp25_ASAP7_75t_SL g823 ( 
.A(n_802),
.B(n_754),
.C(n_775),
.D(n_713),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_804),
.B(n_761),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_786),
.B(n_759),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_786),
.B(n_699),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_790),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_804),
.B(n_759),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_824),
.B(n_805),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_824),
.B(n_805),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_815),
.B(n_802),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_821),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_815),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_821),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_814),
.B(n_789),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_820),
.B(n_793),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_820),
.B(n_793),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_824),
.B(n_809),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_824),
.B(n_795),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_822),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_839),
.B(n_818),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_839),
.Y(n_842)
);

AND2x2_ASAP7_75t_SL g843 ( 
.A(n_829),
.B(n_810),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_838),
.B(n_813),
.Y(n_844)
);

AO22x1_ASAP7_75t_L g845 ( 
.A1(n_829),
.A2(n_816),
.B1(n_828),
.B2(n_818),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_835),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_842),
.B(n_831),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_841),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_846),
.B(n_833),
.Y(n_849)
);

NAND2x1_ASAP7_75t_L g850 ( 
.A(n_841),
.B(n_838),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_844),
.B(n_831),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_844),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_852),
.B(n_843),
.Y(n_853)
);

NAND2x1_ASAP7_75t_L g854 ( 
.A(n_847),
.B(n_829),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_849),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_SL g856 ( 
.A1(n_851),
.A2(n_845),
.B1(n_825),
.B2(n_830),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_851),
.A2(n_843),
.B1(n_828),
.B2(n_830),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_855),
.Y(n_858)
);

OAI32xp33_ASAP7_75t_L g859 ( 
.A1(n_853),
.A2(n_848),
.A3(n_825),
.B1(n_850),
.B2(n_795),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_857),
.A2(n_848),
.B1(n_830),
.B2(n_837),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_856),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_861),
.B(n_854),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_858),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_860),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_859),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_858),
.B(n_836),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_863),
.Y(n_867)
);

XNOR2xp5_ASAP7_75t_L g868 ( 
.A(n_862),
.B(n_828),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_862),
.B(n_836),
.Y(n_869)
);

NOR3x1_ASAP7_75t_L g870 ( 
.A(n_865),
.B(n_753),
.C(n_799),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_866),
.Y(n_871)
);

AOI21xp33_ASAP7_75t_L g872 ( 
.A1(n_864),
.A2(n_811),
.B(n_772),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_863),
.B(n_837),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_865),
.B(n_770),
.C(n_773),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_874),
.A2(n_823),
.B(n_783),
.Y(n_875)
);

AOI221xp5_ASAP7_75t_L g876 ( 
.A1(n_868),
.A2(n_806),
.B1(n_797),
.B2(n_803),
.C(n_828),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_R g877 ( 
.A(n_871),
.B(n_769),
.Y(n_877)
);

OAI211xp5_ASAP7_75t_SL g878 ( 
.A1(n_867),
.A2(n_776),
.B(n_765),
.C(n_788),
.Y(n_878)
);

AOI221xp5_ASAP7_75t_L g879 ( 
.A1(n_869),
.A2(n_797),
.B1(n_806),
.B2(n_803),
.C(n_811),
.Y(n_879)
);

AOI222xp33_ASAP7_75t_L g880 ( 
.A1(n_873),
.A2(n_797),
.B1(n_803),
.B2(n_806),
.C1(n_811),
.C2(n_807),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_870),
.B(n_826),
.Y(n_881)
);

AOI221xp5_ASAP7_75t_L g882 ( 
.A1(n_872),
.A2(n_760),
.B1(n_834),
.B2(n_832),
.C(n_840),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_871),
.Y(n_883)
);

AOI221xp5_ASAP7_75t_L g884 ( 
.A1(n_874),
.A2(n_760),
.B1(n_834),
.B2(n_832),
.C(n_840),
.Y(n_884)
);

AOI211xp5_ASAP7_75t_L g885 ( 
.A1(n_883),
.A2(n_745),
.B(n_734),
.C(n_823),
.Y(n_885)
);

XNOR2x1_ASAP7_75t_L g886 ( 
.A(n_881),
.B(n_768),
.Y(n_886)
);

AO21x2_ASAP7_75t_L g887 ( 
.A1(n_877),
.A2(n_875),
.B(n_878),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_879),
.A2(n_788),
.B(n_808),
.C(n_750),
.Y(n_888)
);

AND2x2_ASAP7_75t_SL g889 ( 
.A(n_882),
.B(n_768),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_884),
.Y(n_890)
);

AOI31xp33_ASAP7_75t_L g891 ( 
.A1(n_876),
.A2(n_768),
.A3(n_782),
.B(n_799),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_880),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_883),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_893),
.B(n_887),
.Y(n_894)
);

NAND4xp25_ASAP7_75t_L g895 ( 
.A(n_890),
.B(n_892),
.C(n_885),
.D(n_888),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_887),
.B(n_789),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_886),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_889),
.B(n_827),
.Y(n_898)
);

OAI22xp33_ASAP7_75t_L g899 ( 
.A1(n_891),
.A2(n_827),
.B1(n_822),
.B2(n_796),
.Y(n_899)
);

NAND4xp75_ASAP7_75t_L g900 ( 
.A(n_889),
.B(n_808),
.C(n_798),
.D(n_801),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_SL g901 ( 
.A(n_894),
.B(n_743),
.C(n_750),
.Y(n_901)
);

AOI211xp5_ASAP7_75t_L g902 ( 
.A1(n_895),
.A2(n_737),
.B(n_801),
.C(n_798),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_900),
.Y(n_903)
);

AOI221xp5_ASAP7_75t_SL g904 ( 
.A1(n_896),
.A2(n_796),
.B1(n_817),
.B2(n_812),
.C(n_819),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_897),
.Y(n_905)
);

NAND4xp25_ASAP7_75t_SL g906 ( 
.A(n_898),
.B(n_792),
.C(n_817),
.D(n_812),
.Y(n_906)
);

BUFx8_ASAP7_75t_L g907 ( 
.A(n_905),
.Y(n_907)
);

OAI221xp5_ASAP7_75t_L g908 ( 
.A1(n_902),
.A2(n_899),
.B1(n_743),
.B2(n_796),
.C(n_819),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_903),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_904),
.B(n_796),
.Y(n_910)
);

OA22x2_ASAP7_75t_L g911 ( 
.A1(n_909),
.A2(n_901),
.B1(n_906),
.B2(n_792),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_907),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_908),
.A2(n_910),
.B1(n_742),
.B2(n_792),
.Y(n_913)
);

OA21x2_ASAP7_75t_L g914 ( 
.A1(n_913),
.A2(n_790),
.B(n_791),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_912),
.A2(n_911),
.B(n_791),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_R g916 ( 
.A1(n_915),
.A2(n_741),
.B1(n_791),
.B2(n_735),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_914),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_917),
.Y(n_918)
);

OAI22xp33_ASAP7_75t_L g919 ( 
.A1(n_916),
.A2(n_739),
.B1(n_713),
.B2(n_708),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_R g920 ( 
.A1(n_918),
.A2(n_133),
.B1(n_136),
.B2(n_139),
.Y(n_920)
);

AOI322xp5_ASAP7_75t_L g921 ( 
.A1(n_920),
.A2(n_919),
.A3(n_142),
.B1(n_143),
.B2(n_144),
.C1(n_146),
.C2(n_147),
.Y(n_921)
);

OAI221xp5_ASAP7_75t_L g922 ( 
.A1(n_921),
.A2(n_141),
.B1(n_150),
.B2(n_152),
.C(n_155),
.Y(n_922)
);

AOI211xp5_ASAP7_75t_L g923 ( 
.A1(n_922),
.A2(n_156),
.B(n_158),
.C(n_162),
.Y(n_923)
);


endmodule