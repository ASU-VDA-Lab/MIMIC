module fake_jpeg_8797_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

CKINVDCx11_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_53),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_65),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_68),
.Y(n_85)
);

NAND2x1_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_35),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_89),
.B1(n_99),
.B2(n_45),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_72),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_75),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_47),
.B1(n_38),
.B2(n_22),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_74),
.A2(n_77),
.B1(n_68),
.B2(n_63),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_47),
.B1(n_38),
.B2(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_87),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_39),
.Y(n_101)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_22),
.B1(n_29),
.B2(n_47),
.Y(n_89)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_95),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_22),
.B1(n_29),
.B2(n_32),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_93),
.B1(n_70),
.B2(n_98),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_103),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_39),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_114),
.B1(n_119),
.B2(n_127),
.Y(n_147)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_110),
.Y(n_150)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

AO22x2_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_48),
.B1(n_45),
.B2(n_37),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_48),
.B(n_37),
.C(n_40),
.Y(n_137)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_116),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_90),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_39),
.B1(n_55),
.B2(n_44),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_124),
.B1(n_126),
.B2(n_92),
.Y(n_155)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_81),
.A2(n_32),
.B1(n_36),
.B2(n_18),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_129),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_60),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_134),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_139),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_105),
.B1(n_87),
.B2(n_83),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_33),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_33),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_152),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_75),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_40),
.B(n_41),
.Y(n_172)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_148),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_153),
.B(n_113),
.Y(n_158)
);

CKINVDCx10_ASAP7_75t_R g151 ( 
.A(n_110),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_46),
.C(n_81),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_156),
.C(n_46),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_73),
.B1(n_88),
.B2(n_96),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_40),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_126),
.B(n_58),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_157),
.A2(n_163),
.B(n_167),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_173),
.B(n_179),
.Y(n_198)
);

OAI22x1_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_100),
.B1(n_106),
.B2(n_35),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_159),
.A2(n_183),
.B1(n_27),
.B2(n_24),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_61),
.B(n_58),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_165),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_105),
.A3(n_93),
.B1(n_98),
.B2(n_106),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_169),
.B(n_175),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_133),
.C(n_148),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_174),
.B1(n_177),
.B2(n_144),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_24),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_145),
.B(n_134),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_121),
.B1(n_120),
.B2(n_48),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_186),
.B1(n_188),
.B2(n_135),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_95),
.B(n_35),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_21),
.B1(n_31),
.B2(n_23),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_31),
.B1(n_95),
.B2(n_27),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_0),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_26),
.B(n_1),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_141),
.A2(n_35),
.B1(n_23),
.B2(n_27),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_190),
.A2(n_34),
.B1(n_25),
.B2(n_26),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_211),
.B(n_213),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_138),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_193),
.B(n_203),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_206),
.C(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_133),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_160),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_209),
.B(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_138),
.Y(n_205)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_146),
.C(n_144),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_217),
.B1(n_34),
.B2(n_25),
.Y(n_241)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_16),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_219),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_27),
.C(n_24),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_234),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_186),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_214),
.C(n_194),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_164),
.B1(n_176),
.B2(n_188),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_238),
.B1(n_216),
.B2(n_217),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_187),
.B(n_182),
.Y(n_230)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_187),
.B(n_183),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_237),
.B1(n_1),
.B2(n_2),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

AO22x1_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_161),
.B1(n_182),
.B2(n_24),
.Y(n_235)
);

NAND2xp67_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_3),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_202),
.A2(n_34),
.B1(n_25),
.B2(n_16),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_26),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_240),
.B(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

CKINVDCx6p67_ASAP7_75t_R g244 ( 
.A(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_0),
.Y(n_245)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_247),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_206),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_191),
.C(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_256),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_209),
.C(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_2),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_262),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_261),
.A2(n_266),
.B(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_244),
.Y(n_263)
);

INVx13_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_265),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_4),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_236),
.B(n_220),
.Y(n_271)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_222),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_252),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_227),
.B1(n_232),
.B2(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_283),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_254),
.A2(n_231),
.B1(n_237),
.B2(n_243),
.Y(n_282)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_SL g283 ( 
.A(n_251),
.B(n_230),
.C(n_235),
.Y(n_283)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_288),
.B(n_269),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_259),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_299),
.C(n_280),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_267),
.Y(n_290)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_250),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_297),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_284),
.B(n_260),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_300),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_273),
.B(n_223),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_256),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_268),
.C(n_247),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_238),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_304),
.C(n_313),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_282),
.C(n_270),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_306),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_286),
.A2(n_272),
.B1(n_276),
.B2(n_249),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_293),
.B(n_271),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_287),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_310),
.B(n_5),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_278),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_4),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_278),
.C(n_221),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_307),
.A2(n_296),
.B1(n_291),
.B2(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_320),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_15),
.B1(n_6),
.B2(n_7),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_5),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_5),
.Y(n_322)
);

NOR4xp25_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_9),
.C(n_11),
.D(n_12),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_302),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_328),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_8),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_301),
.B1(n_11),
.B2(n_12),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_327),
.C(n_325),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_330),
.A2(n_321),
.B(n_315),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.C(n_327),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_324),
.B1(n_316),
.B2(n_331),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_316),
.C(n_11),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_337),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_9),
.Y(n_339)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_13),
.B(n_327),
.Y(n_340)
);


endmodule