module fake_ariane_857_n_2846 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_620, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2846);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2846;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2461;
wire n_2207;
wire n_2702;
wire n_2731;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2529;
wire n_2238;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2271;
wire n_2116;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2495;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1053;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_727;
wire n_699;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1614;
wire n_1162;
wire n_1377;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_887;
wire n_729;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1860;
wire n_1734;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_791;
wire n_876;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1603;
wire n_1370;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2441;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_2503;
wire n_1758;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2723;
wire n_1271;
wire n_2096;
wire n_2556;
wire n_2440;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2324;
wire n_2153;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_2101;
wire n_1934;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2552;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2432;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_2188;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_110),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_391),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_574),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_74),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_393),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_506),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_493),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_10),
.Y(n_635)
);

CKINVDCx14_ASAP7_75t_R g636 ( 
.A(n_43),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_123),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_427),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_402),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_224),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_480),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_588),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_324),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_587),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_222),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_549),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_282),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_552),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_22),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_526),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_600),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_524),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_463),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_501),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_292),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_240),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_508),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_477),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_485),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_182),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_581),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_448),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_113),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_416),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_624),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_189),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_30),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_444),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_428),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_218),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_578),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_583),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_182),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_77),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_229),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_163),
.Y(n_676)
);

CKINVDCx16_ASAP7_75t_R g677 ( 
.A(n_360),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_593),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_59),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_503),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_527),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_490),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_342),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_192),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_387),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_188),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_187),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_376),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_291),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_436),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_335),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_306),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_7),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_449),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_51),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_270),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_509),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_377),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_194),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_254),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_505),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_291),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_32),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_484),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_461),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_539),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_56),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_105),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_76),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_429),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_308),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_96),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_352),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_614),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_550),
.Y(n_715)
);

BUFx5_ASAP7_75t_L g716 ( 
.A(n_5),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_424),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_282),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_145),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_250),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_434),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_8),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_240),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_478),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_560),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_339),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_34),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_404),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_589),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_530),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_32),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_98),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_253),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_285),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_620),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_284),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_123),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_294),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_219),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_3),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_294),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_438),
.Y(n_742)
);

CKINVDCx16_ASAP7_75t_R g743 ( 
.A(n_256),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_460),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_458),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_515),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_270),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_555),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_244),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_479),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_556),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_198),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_613),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_488),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_462),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_18),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_542),
.Y(n_757)
);

CKINVDCx16_ASAP7_75t_R g758 ( 
.A(n_597),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_95),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_143),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_40),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_400),
.Y(n_762)
);

CKINVDCx14_ASAP7_75t_R g763 ( 
.A(n_74),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_121),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_25),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_365),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_544),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_321),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_445),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_586),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_612),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_495),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_222),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_132),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_446),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_231),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_374),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_450),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_529),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_491),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_100),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_439),
.Y(n_782)
);

CKINVDCx14_ASAP7_75t_R g783 ( 
.A(n_437),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_28),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_499),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_390),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_179),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_516),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_611),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_310),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_337),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_546),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_47),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_137),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_623),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_296),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_37),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_415),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_573),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_324),
.Y(n_800)
);

BUFx10_ASAP7_75t_L g801 ( 
.A(n_440),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_105),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_364),
.Y(n_803)
);

CKINVDCx16_ASAP7_75t_R g804 ( 
.A(n_200),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_602),
.Y(n_805)
);

CKINVDCx16_ASAP7_75t_R g806 ( 
.A(n_112),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_510),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_525),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_502),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_221),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_44),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_418),
.Y(n_812)
);

BUFx10_ASAP7_75t_L g813 ( 
.A(n_367),
.Y(n_813)
);

CKINVDCx16_ASAP7_75t_R g814 ( 
.A(n_88),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_441),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_290),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_252),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_205),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_61),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_570),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_442),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_85),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_38),
.Y(n_823)
);

BUFx10_ASAP7_75t_L g824 ( 
.A(n_132),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_266),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_1),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_423),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_519),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_609),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_482),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_251),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_494),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_469),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_409),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_120),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_410),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_347),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_75),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_470),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_507),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_520),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_350),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_51),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_401),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_617),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_604),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_146),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_465),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_474),
.Y(n_849)
);

CKINVDCx16_ASAP7_75t_R g850 ( 
.A(n_172),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_155),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_183),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_197),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_381),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_143),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_265),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_53),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_406),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_73),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_106),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_292),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_134),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_471),
.Y(n_863)
);

BUFx5_ASAP7_75t_L g864 ( 
.A(n_599),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_592),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_594),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_590),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_35),
.Y(n_868)
);

BUFx10_ASAP7_75t_L g869 ( 
.A(n_170),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_497),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_27),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_385),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_475),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_489),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_618),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_625),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_627),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_399),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_464),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_451),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_276),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_26),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_483),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_605),
.Y(n_884)
);

BUFx5_ASAP7_75t_L g885 ( 
.A(n_165),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_398),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_104),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_345),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_621),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_212),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_457),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_64),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_603),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_34),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_619),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_147),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_380),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_22),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_562),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_426),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_548),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_116),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_498),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_204),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_20),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_225),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_566),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_43),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_229),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_414),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_161),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_536),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_511),
.Y(n_913)
);

CKINVDCx16_ASAP7_75t_R g914 ( 
.A(n_348),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_532),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_136),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_8),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_131),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_321),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_185),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_571),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_453),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_243),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_237),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_622),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_540),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_517),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_223),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_41),
.Y(n_929)
);

BUFx10_ASAP7_75t_L g930 ( 
.A(n_541),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_432),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_301),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_94),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_411),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_71),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_537),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_18),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_15),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_230),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_373),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_278),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_431),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_163),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_435),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_20),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_179),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_492),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_545),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_579),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_13),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_208),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_194),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_615),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_181),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_610),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_86),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_150),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_71),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_386),
.Y(n_959)
);

CKINVDCx16_ASAP7_75t_R g960 ( 
.A(n_30),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_591),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_467),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_10),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_226),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_514),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_274),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_49),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_576),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_54),
.Y(n_969)
);

BUFx5_ASAP7_75t_L g970 ( 
.A(n_413),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_500),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_452),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_173),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_580),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_89),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_481),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_241),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_0),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_383),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_454),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_69),
.Y(n_981)
);

BUFx2_ASAP7_75t_SL g982 ( 
.A(n_596),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_553),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_357),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_235),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_9),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_226),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_487),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_60),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_267),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_21),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_372),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_344),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_353),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_521),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_558),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_141),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_60),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_405),
.Y(n_999)
);

BUFx10_ASAP7_75t_L g1000 ( 
.A(n_585),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_565),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_165),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_433),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_504),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_569),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_551),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_21),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_157),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_547),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_326),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_108),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_595),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_616),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_27),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_533),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_472),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_171),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_601),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_24),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_235),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_250),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_110),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_188),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_208),
.Y(n_1024)
);

BUFx10_ASAP7_75t_L g1025 ( 
.A(n_19),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_567),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_420),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_456),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_412),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_512),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_606),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_237),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_189),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_178),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_125),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_199),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_584),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_75),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_626),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_564),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_543),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_252),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_195),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_53),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_486),
.Y(n_1045)
);

CKINVDCx16_ASAP7_75t_R g1046 ( 
.A(n_259),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_210),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_102),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_76),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_161),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_26),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_320),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_598),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_218),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_523),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_216),
.Y(n_1056)
);

INVxp33_ASAP7_75t_SL g1057 ( 
.A(n_128),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_559),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_248),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_5),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_278),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_534),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_407),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_358),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_355),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_473),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_176),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_341),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_275),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_23),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_563),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_572),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_11),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_214),
.Y(n_1074)
);

CKINVDCx14_ASAP7_75t_R g1075 ( 
.A(n_496),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_326),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_134),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_262),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_575),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_211),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_19),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_528),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_45),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_90),
.Y(n_1084)
);

BUFx5_ASAP7_75t_L g1085 ( 
.A(n_568),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_257),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_455),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_169),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_233),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_63),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_35),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_476),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_557),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_140),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_37),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_9),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_397),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_522),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_554),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_443),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_330),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_447),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_518),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_513),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_466),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_531),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_175),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_535),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_538),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_184),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_287),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_29),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_155),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_98),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_318),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_6),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_561),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_459),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_468),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_77),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_138),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_104),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_320),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_608),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_68),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_152),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_135),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_140),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_241),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_39),
.Y(n_1130)
);

CKINVDCx16_ASAP7_75t_R g1131 ( 
.A(n_577),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_58),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_300),
.Y(n_1133)
);

BUFx10_ASAP7_75t_L g1134 ( 
.A(n_170),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_39),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_582),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_607),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_164),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_70),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_164),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_752),
.B(n_0),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_798),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_SL g1143 ( 
.A(n_677),
.B(n_331),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_712),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_SL g1145 ( 
.A(n_758),
.B(n_332),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_712),
.B(n_1),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_822),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_760),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_822),
.Y(n_1149)
);

BUFx8_ASAP7_75t_SL g1150 ( 
.A(n_673),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_878),
.B(n_2),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_760),
.Y(n_1152)
);

BUFx8_ASAP7_75t_L g1153 ( 
.A(n_638),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_801),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_801),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1014),
.B(n_2),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_716),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_716),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_716),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_716),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1014),
.B(n_3),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_878),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1104),
.B(n_4),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_707),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_760),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1104),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_760),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_887),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_716),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_707),
.Y(n_1170)
);

BUFx8_ASAP7_75t_SL g1171 ( 
.A(n_718),
.Y(n_1171)
);

AND2x6_ASAP7_75t_L g1172 ( 
.A(n_634),
.B(n_333),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_780),
.B(n_4),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_839),
.B(n_6),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1057),
.B(n_7),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1102),
.B(n_11),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_743),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_804),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_716),
.Y(n_1179)
);

XNOR2xp5_ASAP7_75t_L g1180 ( 
.A(n_727),
.B(n_12),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_887),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_885),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_636),
.B(n_12),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_798),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_885),
.B(n_630),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_908),
.B(n_13),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_813),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_885),
.B(n_14),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_887),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_806),
.B(n_14),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_634),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_885),
.B(n_15),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_816),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_887),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_SL g1195 ( 
.A(n_914),
.B(n_334),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_636),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_763),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_639),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_885),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_816),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_885),
.B(n_632),
.Y(n_1201)
);

NOR2x1_ASAP7_75t_L g1202 ( 
.A(n_639),
.B(n_336),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_814),
.B(n_16),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_652),
.B(n_16),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_896),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_763),
.B(n_17),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_654),
.B(n_661),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_896),
.Y(n_1208)
);

BUFx8_ASAP7_75t_SL g1209 ( 
.A(n_871),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_668),
.B(n_17),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_818),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_850),
.Y(n_1212)
);

INVx5_ASAP7_75t_L g1213 ( 
.A(n_813),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_960),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_896),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_896),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_678),
.B(n_23),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_989),
.Y(n_1218)
);

BUFx8_ASAP7_75t_SL g1219 ( 
.A(n_881),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_989),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_989),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_681),
.B(n_24),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_682),
.B(n_25),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_989),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1046),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_783),
.B(n_28),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_783),
.B(n_29),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_635),
.Y(n_1228)
);

INVx5_ASAP7_75t_L g1229 ( 
.A(n_930),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1048),
.Y(n_1230)
);

AND2x6_ASAP7_75t_L g1231 ( 
.A(n_767),
.B(n_338),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_911),
.B(n_31),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1075),
.B(n_31),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_688),
.B(n_33),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1075),
.B(n_33),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_690),
.B(n_36),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_957),
.B(n_986),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1094),
.B(n_36),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_704),
.B(n_38),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1048),
.Y(n_1240)
);

BUFx8_ASAP7_75t_SL g1241 ( 
.A(n_956),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1048),
.Y(n_1242)
);

AND2x6_ASAP7_75t_L g1243 ( 
.A(n_767),
.B(n_340),
.Y(n_1243)
);

AND2x6_ASAP7_75t_L g1244 ( 
.A(n_913),
.B(n_343),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_930),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_710),
.B(n_40),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1000),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_724),
.B(n_41),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1048),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_725),
.B(n_42),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_824),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1067),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1116),
.B(n_42),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_628),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1067),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_730),
.B(n_44),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1067),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1067),
.Y(n_1258)
);

BUFx12f_ASAP7_75t_L g1259 ( 
.A(n_1000),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_913),
.B(n_45),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1140),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1027),
.B(n_46),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1140),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_824),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1140),
.Y(n_1265)
);

INVx5_ASAP7_75t_L g1266 ( 
.A(n_1140),
.Y(n_1266)
);

BUFx12f_ASAP7_75t_L g1267 ( 
.A(n_869),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1027),
.B(n_46),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_745),
.B(n_47),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1131),
.B(n_346),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_746),
.B(n_48),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_717),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_717),
.Y(n_1273)
);

INVx5_ASAP7_75t_L g1274 ( 
.A(n_717),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1124),
.B(n_48),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_717),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_751),
.B(n_49),
.Y(n_1277)
);

BUFx12f_ASAP7_75t_L g1278 ( 
.A(n_869),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1124),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_675),
.B(n_50),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_753),
.B(n_50),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_631),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_640),
.Y(n_1283)
);

AND2x6_ASAP7_75t_L g1284 ( 
.A(n_729),
.B(n_349),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_754),
.B(n_52),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1025),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_645),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_675),
.B(n_52),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_762),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1025),
.B(n_54),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_766),
.Y(n_1291)
);

INVx5_ASAP7_75t_L g1292 ( 
.A(n_858),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_676),
.B(n_55),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_676),
.B(n_55),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_696),
.B(n_768),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_696),
.B(n_768),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_649),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1134),
.B(n_56),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_769),
.B(n_57),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_772),
.B(n_57),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_858),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_656),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_666),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_779),
.B(n_58),
.Y(n_1304)
);

INVx4_ASAP7_75t_L g1305 ( 
.A(n_858),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_786),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_803),
.B(n_59),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_692),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_796),
.B(n_61),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1134),
.B(n_729),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_796),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_693),
.Y(n_1312)
);

INVx5_ASAP7_75t_L g1313 ( 
.A(n_858),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1196),
.B(n_853),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1226),
.A2(n_1089),
.B1(n_1081),
.B2(n_1047),
.Y(n_1315)
);

OR2x6_ASAP7_75t_L g1316 ( 
.A(n_1264),
.B(n_924),
.Y(n_1316)
);

OAI22xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1151),
.A2(n_709),
.B1(n_774),
.B2(n_708),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1226),
.A2(n_1107),
.B1(n_1086),
.B2(n_1019),
.Y(n_1318)
);

AO22x2_ASAP7_75t_L g1319 ( 
.A1(n_1162),
.A2(n_920),
.B1(n_987),
.B2(n_793),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1227),
.A2(n_1112),
.B1(n_1137),
.B2(n_691),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1143),
.A2(n_1128),
.B1(n_643),
.B2(n_647),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_SL g1322 ( 
.A(n_1237),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1227),
.A2(n_697),
.B1(n_735),
.B2(n_714),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1233),
.A2(n_820),
.B1(n_841),
.B2(n_778),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1233),
.A2(n_863),
.B1(n_893),
.B2(n_846),
.Y(n_1325)
);

AO22x2_ASAP7_75t_L g1326 ( 
.A1(n_1166),
.A2(n_951),
.B1(n_998),
.B2(n_853),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1235),
.A2(n_922),
.B1(n_974),
.B2(n_910),
.Y(n_1327)
);

AO22x2_ASAP7_75t_L g1328 ( 
.A1(n_1235),
.A2(n_1038),
.B1(n_1061),
.B2(n_998),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1267),
.B(n_1061),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1145),
.A2(n_655),
.B1(n_660),
.B2(n_637),
.Y(n_1330)
);

AO22x2_ASAP7_75t_L g1331 ( 
.A1(n_1183),
.A2(n_1115),
.B1(n_1126),
.B2(n_1038),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1214),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1191),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1212),
.A2(n_1270),
.B1(n_1195),
.B2(n_1177),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1212),
.A2(n_983),
.B1(n_1031),
.B2(n_979),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1196),
.B(n_1115),
.Y(n_1336)
);

OA22x2_ASAP7_75t_L g1337 ( 
.A1(n_1178),
.A2(n_722),
.B1(n_732),
.B2(n_699),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1197),
.B(n_736),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1148),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1183),
.A2(n_1065),
.B1(n_1058),
.B2(n_674),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1197),
.B(n_1126),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1187),
.B(n_904),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1211),
.A2(n_667),
.B1(n_670),
.B2(n_663),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1187),
.B(n_1245),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1163),
.A2(n_686),
.B1(n_687),
.B2(n_679),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1213),
.B(n_973),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1225),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1206),
.A2(n_749),
.B1(n_838),
.B2(n_703),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1148),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1152),
.Y(n_1350)
);

AO22x2_ASAP7_75t_L g1351 ( 
.A1(n_1206),
.A2(n_737),
.B1(n_738),
.B2(n_734),
.Y(n_1351)
);

OAI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1190),
.A2(n_689),
.B1(n_695),
.B2(n_684),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1173),
.A2(n_851),
.B1(n_861),
.B2(n_731),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1203),
.A2(n_1174),
.B1(n_1310),
.B2(n_1141),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1213),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1176),
.A2(n_784),
.B1(n_906),
.B2(n_733),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1290),
.A2(n_797),
.B1(n_810),
.B2(n_739),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1152),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1165),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1290),
.A2(n_773),
.B1(n_800),
.B2(n_740),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1308),
.A2(n_702),
.B1(n_711),
.B2(n_700),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1180),
.A2(n_720),
.B1(n_723),
.B2(n_719),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1182),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1229),
.B(n_1096),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1142),
.B(n_827),
.Y(n_1365)
);

OA22x2_ASAP7_75t_L g1366 ( 
.A1(n_1297),
.A2(n_765),
.B1(n_776),
.B2(n_756),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1298),
.A2(n_856),
.B1(n_950),
.B2(n_823),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1229),
.B(n_787),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1199),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1165),
.Y(n_1370)
);

AO22x2_ASAP7_75t_L g1371 ( 
.A1(n_1298),
.A2(n_794),
.B1(n_817),
.B2(n_790),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1167),
.Y(n_1372)
);

AO22x2_ASAP7_75t_L g1373 ( 
.A1(n_1186),
.A2(n_831),
.B1(n_835),
.B2(n_819),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1279),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1167),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1175),
.A2(n_747),
.B1(n_759),
.B2(n_741),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1207),
.A2(n_764),
.B1(n_802),
.B2(n_781),
.Y(n_1377)
);

OAI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1164),
.A2(n_1129),
.B1(n_1130),
.B2(n_1127),
.Y(n_1378)
);

AO22x2_ASAP7_75t_L g1379 ( 
.A1(n_1232),
.A2(n_847),
.B1(n_852),
.B2(n_843),
.Y(n_1379)
);

OR2x6_ASAP7_75t_L g1380 ( 
.A(n_1278),
.B(n_1139),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1180),
.A2(n_761),
.B1(n_825),
.B2(n_811),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1245),
.B(n_859),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1247),
.B(n_882),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1168),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1184),
.B(n_875),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1254),
.A2(n_1042),
.B1(n_1074),
.B2(n_963),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1247),
.B(n_890),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1204),
.A2(n_855),
.B1(n_857),
.B2(n_826),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1170),
.A2(n_1200),
.B1(n_1251),
.B2(n_1193),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1282),
.B(n_902),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1238),
.A2(n_894),
.B1(n_919),
.B2(n_868),
.Y(n_1391)
);

NAND2xp33_ASAP7_75t_SL g1392 ( 
.A(n_1260),
.B(n_860),
.Y(n_1392)
);

OAI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1286),
.A2(n_892),
.B1(n_898),
.B2(n_862),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1168),
.Y(n_1394)
);

NAND2xp33_ASAP7_75t_SL g1395 ( 
.A(n_1262),
.B(n_916),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1154),
.A2(n_1121),
.B1(n_1122),
.B2(n_1120),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1181),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1289),
.B(n_905),
.Y(n_1398)
);

AO22x2_ASAP7_75t_L g1399 ( 
.A1(n_1253),
.A2(n_917),
.B1(n_923),
.B2(n_909),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1228),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1181),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1189),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1189),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1150),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1155),
.A2(n_928),
.B1(n_929),
.B2(n_918),
.Y(n_1405)
);

AO22x2_ASAP7_75t_L g1406 ( 
.A1(n_1280),
.A2(n_941),
.B1(n_943),
.B2(n_939),
.Y(n_1406)
);

AO22x2_ASAP7_75t_L g1407 ( 
.A1(n_1288),
.A2(n_952),
.B1(n_964),
.B2(n_945),
.Y(n_1407)
);

OR2x6_ASAP7_75t_L g1408 ( 
.A(n_1259),
.B(n_1113),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1198),
.B(n_808),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1291),
.B(n_967),
.Y(n_1410)
);

OAI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1210),
.A2(n_1223),
.B1(n_1234),
.B2(n_1217),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1306),
.Y(n_1412)
);

AO22x2_ASAP7_75t_L g1413 ( 
.A1(n_1293),
.A2(n_985),
.B1(n_1002),
.B2(n_978),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1194),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1268),
.A2(n_1077),
.B1(n_954),
.B2(n_933),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1144),
.B(n_1011),
.Y(n_1416)
);

AO22x2_ASAP7_75t_L g1417 ( 
.A1(n_1294),
.A2(n_1023),
.B1(n_1032),
.B2(n_1022),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1222),
.A2(n_1111),
.B1(n_1114),
.B2(n_1110),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1147),
.B(n_1033),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1283),
.Y(n_1420)
);

OR2x6_ASAP7_75t_L g1421 ( 
.A(n_1311),
.B(n_1135),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1239),
.A2(n_1133),
.B1(n_1138),
.B2(n_1123),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1250),
.A2(n_935),
.B1(n_937),
.B2(n_932),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1275),
.A2(n_990),
.B1(n_1020),
.B2(n_975),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1236),
.A2(n_1095),
.B1(n_1051),
.B2(n_946),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1287),
.Y(n_1426)
);

AOI22x1_ASAP7_75t_SL g1427 ( 
.A1(n_1171),
.A2(n_1076),
.B1(n_977),
.B2(n_958),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1256),
.A2(n_966),
.B1(n_969),
.B2(n_938),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1246),
.A2(n_1036),
.B1(n_1049),
.B2(n_1021),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1269),
.A2(n_991),
.B1(n_997),
.B2(n_981),
.Y(n_1430)
);

AND2x2_ASAP7_75t_SL g1431 ( 
.A(n_1309),
.B(n_1146),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1156),
.B(n_744),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1194),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1271),
.A2(n_1008),
.B1(n_1010),
.B2(n_1007),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1248),
.A2(n_1307),
.B1(n_1277),
.B2(n_1285),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1299),
.A2(n_1024),
.B1(n_1034),
.B2(n_1017),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1281),
.A2(n_1090),
.B1(n_1060),
.B2(n_1069),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1303),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1149),
.B(n_1035),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1157),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1208),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1161),
.A2(n_1070),
.B1(n_1073),
.B2(n_1059),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1272),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1209),
.A2(n_1091),
.B1(n_1088),
.B2(n_1125),
.Y(n_1444)
);

AO22x2_ASAP7_75t_L g1445 ( 
.A1(n_1295),
.A2(n_1044),
.B1(n_1050),
.B2(n_1043),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1208),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1300),
.A2(n_1054),
.B1(n_1056),
.B2(n_1052),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1266),
.B(n_809),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1304),
.A2(n_1080),
.B1(n_1083),
.B2(n_1078),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1296),
.B(n_1084),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1188),
.A2(n_1132),
.B1(n_971),
.B2(n_1026),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1215),
.Y(n_1452)
);

AO22x2_ASAP7_75t_L g1453 ( 
.A1(n_1311),
.A2(n_658),
.B1(n_680),
.B2(n_657),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1158),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1192),
.A2(n_921),
.B1(n_1136),
.B2(n_897),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1215),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1302),
.B(n_791),
.Y(n_1457)
);

AO22x2_ASAP7_75t_L g1458 ( 
.A1(n_1312),
.A2(n_884),
.B1(n_961),
.B2(n_867),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1172),
.A2(n_1040),
.B1(n_650),
.B2(n_651),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1266),
.B(n_982),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1185),
.B(n_840),
.Y(n_1461)
);

AO22x2_ASAP7_75t_L g1462 ( 
.A1(n_1201),
.A2(n_744),
.B1(n_994),
.B2(n_830),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1273),
.B(n_642),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1216),
.Y(n_1464)
);

AO22x2_ASAP7_75t_L g1465 ( 
.A1(n_1205),
.A2(n_994),
.B1(n_1029),
.B2(n_830),
.Y(n_1465)
);

AO22x2_ASAP7_75t_L g1466 ( 
.A1(n_1218),
.A2(n_1045),
.B1(n_1064),
.B2(n_1029),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1216),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1153),
.A2(n_1064),
.B1(n_1045),
.B2(n_785),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1273),
.B(n_972),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1313),
.B(n_1274),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1202),
.A2(n_845),
.B1(n_865),
.B2(n_849),
.Y(n_1471)
);

AO22x2_ASAP7_75t_L g1472 ( 
.A1(n_1220),
.A2(n_953),
.B1(n_872),
.B2(n_874),
.Y(n_1472)
);

AND2x2_ASAP7_75t_SL g1473 ( 
.A(n_1219),
.B(n_671),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1159),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1172),
.A2(n_879),
.B1(n_888),
.B2(n_866),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1241),
.A2(n_903),
.B1(n_907),
.B2(n_899),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1172),
.A2(n_984),
.B1(n_992),
.B2(n_940),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1240),
.A2(n_996),
.B1(n_1009),
.B2(n_995),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1305),
.B(n_1053),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1231),
.A2(n_1055),
.B1(n_1063),
.B2(n_1018),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1221),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1242),
.A2(n_1093),
.B1(n_1100),
.B2(n_1082),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_R g1483 ( 
.A1(n_1258),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1160),
.A2(n_1106),
.B1(n_1087),
.B2(n_633),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1221),
.A2(n_641),
.B1(n_644),
.B2(n_629),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_R g1486 ( 
.A1(n_1169),
.A2(n_66),
.B1(n_62),
.B2(n_65),
.Y(n_1486)
);

OAI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1179),
.A2(n_653),
.B1(n_659),
.B2(n_646),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1274),
.B(n_891),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1231),
.A2(n_664),
.B1(n_665),
.B2(n_648),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1224),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1292),
.B(n_1117),
.Y(n_1491)
);

OAI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1231),
.A2(n_672),
.B1(n_683),
.B2(n_662),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1243),
.A2(n_685),
.B1(n_694),
.B2(n_669),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1224),
.A2(n_701),
.B1(n_705),
.B2(n_698),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1292),
.B(n_706),
.Y(n_1495)
);

OAI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1230),
.A2(n_715),
.B1(n_721),
.B2(n_713),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1230),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1249),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1249),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1252),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1252),
.Y(n_1501)
);

CKINVDCx6p67_ASAP7_75t_R g1502 ( 
.A(n_1243),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1255),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1243),
.A2(n_728),
.B1(n_742),
.B2(n_726),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1244),
.A2(n_750),
.B1(n_755),
.B2(n_748),
.Y(n_1505)
);

AO22x2_ASAP7_75t_L g1506 ( 
.A1(n_1244),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1255),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1244),
.A2(n_770),
.B1(n_771),
.B2(n_757),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1284),
.A2(n_777),
.B1(n_782),
.B2(n_775),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_SL g1510 ( 
.A1(n_1257),
.A2(n_789),
.B1(n_792),
.B2(n_788),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1313),
.B(n_795),
.Y(n_1511)
);

OR2x6_ASAP7_75t_L g1512 ( 
.A(n_1257),
.B(n_891),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1261),
.B(n_799),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1261),
.B(n_805),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1263),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1284),
.A2(n_812),
.B1(n_815),
.B2(n_807),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1263),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1265),
.B(n_821),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1265),
.B(n_828),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1272),
.A2(n_832),
.B1(n_833),
.B2(n_829),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1284),
.A2(n_836),
.B1(n_837),
.B2(n_834),
.Y(n_1521)
);

AND2x2_ASAP7_75t_SL g1522 ( 
.A(n_1276),
.B(n_891),
.Y(n_1522)
);

OAI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1276),
.A2(n_844),
.B1(n_848),
.B2(n_842),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1301),
.A2(n_870),
.B1(n_873),
.B2(n_854),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1301),
.A2(n_876),
.B1(n_880),
.B2(n_877),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1182),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1212),
.A2(n_886),
.B1(n_889),
.B2(n_883),
.Y(n_1527)
);

OAI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1151),
.A2(n_900),
.B1(n_901),
.B2(n_895),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1182),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1196),
.B(n_912),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1180),
.A2(n_915),
.B1(n_926),
.B2(n_925),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1177),
.B(n_67),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1264),
.B(n_891),
.Y(n_1533)
);

INVx8_ASAP7_75t_L g1534 ( 
.A(n_1154),
.Y(n_1534)
);

AO22x2_ASAP7_75t_L g1535 ( 
.A1(n_1162),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1535)
);

OAI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1212),
.A2(n_934),
.B1(n_936),
.B2(n_927),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1142),
.B(n_942),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1191),
.Y(n_1538)
);

OA22x2_ASAP7_75t_L g1539 ( 
.A1(n_1162),
.A2(n_947),
.B1(n_948),
.B2(n_944),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1148),
.Y(n_1540)
);

OAI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1212),
.A2(n_949),
.B1(n_959),
.B2(n_955),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1214),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1148),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1142),
.B(n_962),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1196),
.B(n_931),
.Y(n_1545)
);

AO22x2_ASAP7_75t_L g1546 ( 
.A1(n_1162),
.A2(n_78),
.B1(n_72),
.B2(n_73),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1180),
.A2(n_965),
.B1(n_976),
.B2(n_968),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1272),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1151),
.A2(n_988),
.B1(n_993),
.B2(n_980),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1226),
.A2(n_1001),
.B1(n_1004),
.B2(n_999),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1151),
.A2(n_1006),
.B1(n_1013),
.B2(n_1005),
.Y(n_1551)
);

OAI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1212),
.A2(n_1016),
.B1(n_1028),
.B2(n_1015),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1142),
.B(n_1037),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1196),
.B(n_1039),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1142),
.B(n_1041),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1226),
.A2(n_1066),
.B1(n_1068),
.B2(n_1062),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1212),
.A2(n_1072),
.B1(n_1079),
.B2(n_1071),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1226),
.A2(n_1097),
.B1(n_1098),
.B2(n_1092),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1182),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1182),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1196),
.B(n_1099),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1177),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1148),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1182),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1226),
.A2(n_1103),
.B1(n_1105),
.B2(n_1101),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1148),
.Y(n_1566)
);

AO22x2_ASAP7_75t_L g1567 ( 
.A1(n_1162),
.A2(n_79),
.B1(n_72),
.B2(n_78),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_SL g1568 ( 
.A(n_1183),
.B(n_931),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1191),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1212),
.A2(n_1109),
.B1(n_1118),
.B2(n_1108),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1182),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1151),
.A2(n_1119),
.B1(n_81),
.B2(n_79),
.Y(n_1572)
);

AO22x2_ASAP7_75t_L g1573 ( 
.A1(n_1162),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1148),
.Y(n_1574)
);

OAI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1151),
.A2(n_83),
.B1(n_80),
.B2(n_82),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1148),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1180),
.A2(n_1003),
.B1(n_1012),
.B2(n_931),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1226),
.A2(n_931),
.B1(n_1012),
.B2(n_1003),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1177),
.B(n_83),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1226),
.A2(n_1012),
.B1(n_1030),
.B2(n_1003),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1226),
.A2(n_1012),
.B1(n_1030),
.B2(n_1003),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1148),
.Y(n_1582)
);

AO22x2_ASAP7_75t_L g1583 ( 
.A1(n_1162),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1196),
.B(n_1030),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1187),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1180),
.A2(n_1030),
.B1(n_88),
.B2(n_84),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_SL g1587 ( 
.A(n_1143),
.B(n_864),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1142),
.B(n_864),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1226),
.A2(n_970),
.B1(n_1085),
.B2(n_864),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1148),
.Y(n_1590)
);

AO22x2_ASAP7_75t_L g1591 ( 
.A1(n_1162),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1180),
.A2(n_92),
.B1(n_87),
.B2(n_91),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1182),
.Y(n_1593)
);

AO22x2_ASAP7_75t_L g1594 ( 
.A1(n_1162),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1182),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1151),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1196),
.B(n_864),
.Y(n_1597)
);

AO22x2_ASAP7_75t_L g1598 ( 
.A1(n_1162),
.A2(n_99),
.B1(n_96),
.B2(n_97),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1177),
.B(n_97),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_SL g1600 ( 
.A(n_1237),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1142),
.B(n_864),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1226),
.A2(n_970),
.B1(n_1085),
.B2(n_864),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1182),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1182),
.Y(n_1604)
);

BUFx10_ASAP7_75t_L g1605 ( 
.A(n_1190),
.Y(n_1605)
);

AO22x2_ASAP7_75t_L g1606 ( 
.A1(n_1162),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1606)
);

AO22x2_ASAP7_75t_L g1607 ( 
.A1(n_1162),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1182),
.Y(n_1608)
);

OAI22xp33_ASAP7_75t_R g1609 ( 
.A1(n_1175),
.A2(n_107),
.B1(n_103),
.B2(n_106),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1226),
.A2(n_1085),
.B1(n_970),
.B2(n_109),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1226),
.A2(n_1085),
.B1(n_970),
.B2(n_109),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1196),
.B(n_970),
.Y(n_1612)
);

OAI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1212),
.A2(n_111),
.B1(n_107),
.B2(n_108),
.Y(n_1613)
);

AO22x2_ASAP7_75t_L g1614 ( 
.A1(n_1162),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1182),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1142),
.B(n_1085),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1196),
.B(n_970),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1182),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1196),
.B(n_1085),
.Y(n_1619)
);

OA22x2_ASAP7_75t_L g1620 ( 
.A1(n_1162),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1620)
);

AO22x2_ASAP7_75t_L g1621 ( 
.A1(n_1162),
.A2(n_117),
.B1(n_114),
.B2(n_115),
.Y(n_1621)
);

AO22x2_ASAP7_75t_L g1622 ( 
.A1(n_1162),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1180),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1148),
.Y(n_1624)
);

AO22x2_ASAP7_75t_L g1625 ( 
.A1(n_1162),
.A2(n_124),
.B1(n_121),
.B2(n_122),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1148),
.Y(n_1626)
);

OAI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1212),
.A2(n_125),
.B1(n_122),
.B2(n_124),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1196),
.B(n_126),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1187),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1196),
.B(n_126),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1226),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1187),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1148),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1226),
.A2(n_130),
.B1(n_127),
.B2(n_129),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1148),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1182),
.Y(n_1636)
);

INVx4_ASAP7_75t_L g1637 ( 
.A(n_1187),
.Y(n_1637)
);

AO22x2_ASAP7_75t_L g1638 ( 
.A1(n_1162),
.A2(n_133),
.B1(n_130),
.B2(n_131),
.Y(n_1638)
);

OA22x2_ASAP7_75t_L g1639 ( 
.A1(n_1162),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1182),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1177),
.B(n_137),
.Y(n_1641)
);

OAI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1212),
.A2(n_141),
.B1(n_138),
.B2(n_139),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1148),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1148),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1226),
.A2(n_144),
.B1(n_139),
.B2(n_142),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1212),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_1646)
);

AOI22x1_ASAP7_75t_L g1647 ( 
.A1(n_1260),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1214),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1148),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1374),
.Y(n_1650)
);

XNOR2xp5_ASAP7_75t_L g1651 ( 
.A(n_1335),
.B(n_148),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1333),
.B(n_149),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1400),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1420),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1426),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1438),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1363),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1538),
.B(n_149),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1584),
.B(n_150),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1369),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1569),
.B(n_151),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1332),
.B(n_151),
.Y(n_1662)
);

XOR2xp5_ASAP7_75t_L g1663 ( 
.A(n_1323),
.B(n_152),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1597),
.B(n_153),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1526),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1529),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_SL g1667 ( 
.A(n_1587),
.B(n_153),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1440),
.Y(n_1668)
);

XOR2xp5_ASAP7_75t_L g1669 ( 
.A(n_1324),
.B(n_154),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1562),
.B(n_154),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1589),
.A2(n_354),
.B(n_351),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1559),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_1443),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1534),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1560),
.Y(n_1675)
);

XOR2xp5_ASAP7_75t_L g1676 ( 
.A(n_1325),
.B(n_156),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1411),
.B(n_156),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1564),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1412),
.B(n_157),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1571),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1593),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1602),
.A2(n_359),
.B(n_356),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1542),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1545),
.B(n_158),
.Y(n_1684)
);

XOR2x2_ASAP7_75t_L g1685 ( 
.A(n_1315),
.B(n_1318),
.Y(n_1685)
);

BUFx5_ASAP7_75t_L g1686 ( 
.A(n_1454),
.Y(n_1686)
);

XOR2xp5_ASAP7_75t_L g1687 ( 
.A(n_1327),
.B(n_158),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1347),
.B(n_159),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1595),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1474),
.Y(n_1690)
);

NAND2x1p5_ASAP7_75t_L g1691 ( 
.A(n_1522),
.B(n_159),
.Y(n_1691)
);

INVx3_ASAP7_75t_R g1692 ( 
.A(n_1648),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1443),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1537),
.B(n_160),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1603),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1604),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1608),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1615),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1544),
.B(n_160),
.Y(n_1699)
);

XOR2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1610),
.B(n_1611),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1618),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1534),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1636),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1640),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1419),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1588),
.A2(n_1616),
.B(n_1601),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1439),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1339),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_SL g1709 ( 
.A(n_1334),
.B(n_1577),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1457),
.B(n_162),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1416),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1450),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1532),
.B(n_162),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1612),
.B(n_166),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1398),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1410),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1488),
.Y(n_1717)
);

INVxp33_ASAP7_75t_L g1718 ( 
.A(n_1362),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1617),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1530),
.B(n_166),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1619),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1513),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_1518),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1404),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1490),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1498),
.Y(n_1726)
);

AND2x6_ASAP7_75t_L g1727 ( 
.A(n_1475),
.B(n_361),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_1531),
.Y(n_1728)
);

INVxp33_ASAP7_75t_L g1729 ( 
.A(n_1381),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1554),
.B(n_1561),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1503),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1507),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1349),
.Y(n_1733)
);

XOR2xp5_ASAP7_75t_L g1734 ( 
.A(n_1547),
.B(n_167),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1515),
.Y(n_1735)
);

AND2x2_ASAP7_75t_SL g1736 ( 
.A(n_1473),
.B(n_167),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1435),
.B(n_168),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1517),
.Y(n_1738)
);

XOR2xp5_ASAP7_75t_L g1739 ( 
.A(n_1320),
.B(n_168),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1421),
.B(n_169),
.Y(n_1740)
);

INVx2_ASAP7_75t_SL g1741 ( 
.A(n_1533),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1368),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1460),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1550),
.B(n_1556),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1382),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1383),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1387),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1314),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1527),
.B(n_171),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1336),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1341),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1533),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1350),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1649),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1358),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1359),
.Y(n_1756)
);

NOR2xp67_ASAP7_75t_L g1757 ( 
.A(n_1637),
.B(n_1355),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1461),
.A2(n_363),
.B(n_362),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1370),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1372),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1375),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1579),
.B(n_172),
.Y(n_1762)
);

NOR2xp67_ASAP7_75t_L g1763 ( 
.A(n_1585),
.B(n_366),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1384),
.Y(n_1764)
);

BUFx3_ASAP7_75t_L g1765 ( 
.A(n_1344),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1394),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1397),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1401),
.Y(n_1768)
);

XNOR2x2_ASAP7_75t_L g1769 ( 
.A(n_1458),
.B(n_173),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1402),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1403),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1433),
.Y(n_1772)
);

XNOR2xp5_ASAP7_75t_L g1773 ( 
.A(n_1340),
.B(n_174),
.Y(n_1773)
);

XOR2xp5_ASAP7_75t_L g1774 ( 
.A(n_1427),
.B(n_174),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1421),
.B(n_175),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1441),
.Y(n_1776)
);

NOR2xp67_ASAP7_75t_L g1777 ( 
.A(n_1629),
.B(n_368),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1452),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1456),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1605),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1464),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1558),
.B(n_176),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1553),
.B(n_1555),
.Y(n_1783)
);

AND2x2_ASAP7_75t_SL g1784 ( 
.A(n_1431),
.B(n_177),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1467),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1481),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1497),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1499),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1500),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1501),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1540),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1338),
.B(n_177),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1565),
.B(n_1365),
.Y(n_1793)
);

INVxp33_ASAP7_75t_L g1794 ( 
.A(n_1342),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1543),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1385),
.B(n_178),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1563),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1566),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1574),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1536),
.B(n_180),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1576),
.Y(n_1801)
);

INVx1_ASAP7_75t_SL g1802 ( 
.A(n_1346),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1541),
.B(n_180),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1582),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1590),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1624),
.Y(n_1806)
);

INVxp33_ASAP7_75t_L g1807 ( 
.A(n_1364),
.Y(n_1807)
);

INVxp67_ASAP7_75t_SL g1808 ( 
.A(n_1470),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1626),
.Y(n_1809)
);

INVxp33_ASAP7_75t_L g1810 ( 
.A(n_1390),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1633),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1635),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1406),
.B(n_181),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1406),
.B(n_183),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1469),
.B(n_184),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1643),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1644),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1407),
.B(n_185),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1552),
.B(n_186),
.Y(n_1819)
);

CKINVDCx16_ASAP7_75t_R g1820 ( 
.A(n_1408),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1414),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1446),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1548),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1557),
.B(n_186),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1432),
.A2(n_370),
.B(n_369),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1407),
.B(n_187),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1570),
.B(n_190),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1491),
.B(n_190),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1322),
.Y(n_1829)
);

CKINVDCx20_ASAP7_75t_R g1830 ( 
.A(n_1405),
.Y(n_1830)
);

INVx4_ASAP7_75t_L g1831 ( 
.A(n_1502),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1366),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1465),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1465),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1354),
.B(n_191),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1466),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1413),
.B(n_191),
.Y(n_1837)
);

XNOR2xp5_ASAP7_75t_L g1838 ( 
.A(n_1444),
.B(n_192),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_R g1839 ( 
.A(n_1329),
.B(n_193),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1389),
.B(n_193),
.Y(n_1840)
);

AND2x6_ASAP7_75t_L g1841 ( 
.A(n_1477),
.B(n_371),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1466),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1448),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1479),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1628),
.B(n_195),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1348),
.B(n_196),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1328),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1391),
.B(n_196),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1328),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1548),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1331),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1331),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1568),
.A2(n_378),
.B(n_375),
.Y(n_1853)
);

NAND2xp33_ASAP7_75t_R g1854 ( 
.A(n_1329),
.B(n_197),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1512),
.Y(n_1855)
);

INVx4_ASAP7_75t_SL g1856 ( 
.A(n_1600),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1512),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1463),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1409),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1630),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1326),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1326),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1495),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1337),
.Y(n_1864)
);

OR2x2_ASAP7_75t_SL g1865 ( 
.A(n_1599),
.B(n_198),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1511),
.B(n_199),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1506),
.Y(n_1867)
);

INVxp33_ASAP7_75t_SL g1868 ( 
.A(n_1510),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1413),
.B(n_200),
.Y(n_1869)
);

INVxp33_ASAP7_75t_L g1870 ( 
.A(n_1641),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1632),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1506),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1445),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1417),
.B(n_1351),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1459),
.B(n_201),
.Y(n_1875)
);

INVx3_ASAP7_75t_R g1876 ( 
.A(n_1316),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1445),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1514),
.Y(n_1878)
);

XOR2xp5_ASAP7_75t_L g1879 ( 
.A(n_1386),
.B(n_201),
.Y(n_1879)
);

XOR2x2_ASAP7_75t_L g1880 ( 
.A(n_1357),
.B(n_202),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1417),
.B(n_202),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1472),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1519),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1462),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1351),
.B(n_203),
.Y(n_1885)
);

OR2x6_ASAP7_75t_L g1886 ( 
.A(n_1380),
.B(n_203),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1462),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1371),
.B(n_204),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1472),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1447),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1449),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1539),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1415),
.B(n_205),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1424),
.B(n_1353),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1373),
.Y(n_1895)
);

BUFx6f_ASAP7_75t_SL g1896 ( 
.A(n_1316),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1371),
.B(n_206),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1373),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1379),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1379),
.Y(n_1900)
);

OR2x6_ASAP7_75t_L g1901 ( 
.A(n_1380),
.B(n_206),
.Y(n_1901)
);

XOR2xp5_ASAP7_75t_L g1902 ( 
.A(n_1442),
.B(n_1528),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1399),
.Y(n_1903)
);

INVxp33_ASAP7_75t_L g1904 ( 
.A(n_1319),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1480),
.B(n_207),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1408),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1399),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1451),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1493),
.B(n_207),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1360),
.B(n_209),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1455),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1356),
.B(n_209),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1487),
.B(n_210),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1647),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1631),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1634),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1645),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1578),
.Y(n_1918)
);

CKINVDCx20_ASAP7_75t_R g1919 ( 
.A(n_1367),
.Y(n_1919)
);

INVxp33_ASAP7_75t_L g1920 ( 
.A(n_1319),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1580),
.Y(n_1921)
);

AND2x6_ASAP7_75t_L g1922 ( 
.A(n_1504),
.B(n_379),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1581),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1425),
.B(n_211),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1330),
.Y(n_1925)
);

XOR2x2_ASAP7_75t_L g1926 ( 
.A(n_1321),
.B(n_212),
.Y(n_1926)
);

AND2x2_ASAP7_75t_SL g1927 ( 
.A(n_1505),
.B(n_213),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1478),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1508),
.B(n_213),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1429),
.B(n_214),
.Y(n_1930)
);

INVxp67_ASAP7_75t_L g1931 ( 
.A(n_1437),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1378),
.B(n_215),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1524),
.Y(n_1933)
);

XOR2xp5_ASAP7_75t_L g1934 ( 
.A(n_1549),
.B(n_215),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1551),
.B(n_216),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1620),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1639),
.Y(n_1937)
);

XNOR2xp5_ASAP7_75t_L g1938 ( 
.A(n_1458),
.B(n_217),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1482),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1471),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1418),
.B(n_217),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1453),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1453),
.B(n_1525),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1509),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1646),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1535),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_SL g1947 ( 
.A(n_1476),
.B(n_219),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1516),
.B(n_220),
.Y(n_1948)
);

XOR2x2_ASAP7_75t_L g1949 ( 
.A(n_1352),
.B(n_220),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1422),
.B(n_221),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1535),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1546),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1521),
.B(n_223),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1546),
.B(n_224),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1567),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1567),
.Y(n_1956)
);

XOR2xp5_ASAP7_75t_L g1957 ( 
.A(n_1376),
.B(n_225),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1573),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1573),
.B(n_227),
.Y(n_1959)
);

XNOR2xp5_ASAP7_75t_L g1960 ( 
.A(n_1468),
.B(n_227),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1583),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1583),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1591),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1591),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_SL g1965 ( 
.A(n_1343),
.B(n_228),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1428),
.B(n_228),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1520),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1594),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1489),
.B(n_230),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1594),
.Y(n_1970)
);

CKINVDCx20_ASAP7_75t_R g1971 ( 
.A(n_1392),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1598),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1668),
.Y(n_1973)
);

AND2x2_ASAP7_75t_SL g1974 ( 
.A(n_1927),
.B(n_1609),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1657),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1810),
.B(n_1598),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1673),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1690),
.Y(n_1978)
);

BUFx3_ASAP7_75t_L g1979 ( 
.A(n_1724),
.Y(n_1979)
);

BUFx6f_ASAP7_75t_L g1980 ( 
.A(n_1673),
.Y(n_1980)
);

INVx2_ASAP7_75t_SL g1981 ( 
.A(n_1683),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1730),
.B(n_1606),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1859),
.B(n_1492),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1741),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1844),
.B(n_1430),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1783),
.B(n_1436),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1829),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1708),
.Y(n_1988)
);

AND2x4_ASAP7_75t_L g1989 ( 
.A(n_1831),
.B(n_1395),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1711),
.B(n_1606),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1733),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1768),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1674),
.Y(n_1993)
);

BUFx3_ASAP7_75t_L g1994 ( 
.A(n_1702),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1660),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1831),
.B(n_231),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1793),
.B(n_1719),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1931),
.B(n_1396),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1721),
.B(n_1484),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1802),
.B(n_1607),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1944),
.B(n_1345),
.Y(n_2001)
);

INVxp67_ASAP7_75t_L g2002 ( 
.A(n_1662),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1665),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1748),
.B(n_1750),
.Y(n_2004)
);

INVx3_ASAP7_75t_L g2005 ( 
.A(n_1771),
.Y(n_2005)
);

INVx4_ASAP7_75t_L g2006 ( 
.A(n_1856),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1751),
.B(n_1607),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1786),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1666),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1816),
.Y(n_2010)
);

INVx3_ASAP7_75t_L g2011 ( 
.A(n_1673),
.Y(n_2011)
);

INVx4_ASAP7_75t_L g2012 ( 
.A(n_1856),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1692),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1878),
.B(n_1485),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1672),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1650),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1675),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1883),
.B(n_1494),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1744),
.B(n_1496),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1737),
.B(n_1572),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1870),
.B(n_1614),
.Y(n_2021)
);

BUFx4f_ASAP7_75t_L g2022 ( 
.A(n_1906),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1693),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1693),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1693),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1753),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_1740),
.Y(n_2027)
);

AND2x2_ASAP7_75t_SL g2028 ( 
.A(n_1784),
.B(n_1486),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1911),
.B(n_1317),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1678),
.Y(n_2030)
);

INVx4_ASAP7_75t_L g2031 ( 
.A(n_1906),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1752),
.B(n_1614),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1680),
.Y(n_2033)
);

INVx4_ASAP7_75t_L g2034 ( 
.A(n_1906),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1780),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_1740),
.Y(n_2036)
);

BUFx6f_ASAP7_75t_L g2037 ( 
.A(n_1743),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1754),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1684),
.B(n_232),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1688),
.B(n_1621),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1681),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1755),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_1765),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1794),
.B(n_1621),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1807),
.B(n_1622),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1689),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1914),
.B(n_1377),
.Y(n_2047)
);

INVx2_ASAP7_75t_SL g2048 ( 
.A(n_1684),
.Y(n_2048)
);

AND2x6_ASAP7_75t_L g2049 ( 
.A(n_1867),
.B(n_1483),
.Y(n_2049)
);

INVx1_ASAP7_75t_SL g2050 ( 
.A(n_1775),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1756),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1759),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1695),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1696),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1715),
.B(n_1622),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1760),
.Y(n_2056)
);

OR2x6_ASAP7_75t_L g2057 ( 
.A(n_1886),
.B(n_1586),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1761),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1697),
.B(n_1388),
.Y(n_2059)
);

AND2x2_ASAP7_75t_SL g2060 ( 
.A(n_1709),
.B(n_1592),
.Y(n_2060)
);

INVx4_ASAP7_75t_L g2061 ( 
.A(n_1775),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1716),
.B(n_1625),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1896),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1723),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_1894),
.B(n_1393),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1698),
.B(n_1423),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1764),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1967),
.B(n_1434),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1701),
.B(n_1575),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1703),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1766),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1823),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1767),
.Y(n_2073)
);

OAI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1706),
.A2(n_1523),
.B(n_1361),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1670),
.B(n_1625),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1704),
.B(n_1596),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1813),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1874),
.B(n_1638),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1814),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1667),
.B(n_1613),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1770),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1686),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_1818),
.Y(n_2083)
);

INVx2_ASAP7_75t_SL g2084 ( 
.A(n_1933),
.Y(n_2084)
);

BUFx3_ASAP7_75t_L g2085 ( 
.A(n_1850),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_1873),
.B(n_232),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_1712),
.B(n_1820),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1843),
.B(n_1638),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1808),
.B(n_1627),
.Y(n_2089)
);

OAI21xp5_ASAP7_75t_L g2090 ( 
.A1(n_1694),
.A2(n_1642),
.B(n_384),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1705),
.B(n_1707),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1912),
.B(n_1623),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1710),
.B(n_233),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1772),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1860),
.B(n_234),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_1965),
.B(n_234),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1653),
.B(n_236),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1654),
.B(n_236),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1686),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1655),
.Y(n_2100)
);

INVxp67_ASAP7_75t_L g2101 ( 
.A(n_1800),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1792),
.B(n_238),
.Y(n_2102)
);

INVxp67_ASAP7_75t_L g2103 ( 
.A(n_1803),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_1826),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1924),
.B(n_238),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1656),
.B(n_239),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1924),
.B(n_239),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1893),
.B(n_242),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1863),
.B(n_242),
.Y(n_2109)
);

AND2x2_ASAP7_75t_SL g2110 ( 
.A(n_1736),
.B(n_243),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_1871),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1908),
.B(n_1918),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1921),
.B(n_244),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1893),
.B(n_245),
.Y(n_2114)
);

BUFx3_ASAP7_75t_L g2115 ( 
.A(n_1821),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1686),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1888),
.B(n_245),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1923),
.B(n_246),
.Y(n_2118)
);

NAND2xp33_ASAP7_75t_SL g2119 ( 
.A(n_1876),
.B(n_246),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1897),
.B(n_247),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_1837),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1659),
.B(n_247),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1885),
.B(n_248),
.Y(n_2123)
);

BUFx4f_ASAP7_75t_L g2124 ( 
.A(n_1691),
.Y(n_2124)
);

INVx2_ASAP7_75t_SL g2125 ( 
.A(n_1720),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1718),
.B(n_249),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1729),
.B(n_249),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1677),
.B(n_251),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_1869),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_1877),
.B(n_253),
.Y(n_2130)
);

AND2x2_ASAP7_75t_SL g2131 ( 
.A(n_1947),
.B(n_254),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1782),
.B(n_255),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1796),
.B(n_1928),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_1776),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1778),
.Y(n_2135)
);

BUFx4f_ASAP7_75t_SL g2136 ( 
.A(n_1971),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1725),
.Y(n_2137)
);

AND2x2_ASAP7_75t_SL g2138 ( 
.A(n_1954),
.B(n_255),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_1895),
.B(n_256),
.Y(n_2139)
);

AND2x4_ASAP7_75t_L g2140 ( 
.A(n_1898),
.B(n_257),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_1679),
.Y(n_2141)
);

INVx4_ASAP7_75t_L g2142 ( 
.A(n_1922),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1779),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1726),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1881),
.B(n_1742),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1745),
.B(n_258),
.Y(n_2146)
);

BUFx3_ASAP7_75t_L g2147 ( 
.A(n_1822),
.Y(n_2147)
);

BUFx2_ASAP7_75t_L g2148 ( 
.A(n_1930),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_1896),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_1846),
.B(n_258),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1746),
.B(n_259),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1731),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1940),
.B(n_260),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1732),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_1899),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1686),
.Y(n_2156)
);

INVxp67_ASAP7_75t_L g2157 ( 
.A(n_1824),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1747),
.B(n_260),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1910),
.B(n_261),
.Y(n_2159)
);

BUFx3_ASAP7_75t_L g2160 ( 
.A(n_1855),
.Y(n_2160)
);

BUFx3_ASAP7_75t_L g2161 ( 
.A(n_1857),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1939),
.B(n_261),
.Y(n_2162)
);

HB1xp67_ASAP7_75t_L g2163 ( 
.A(n_1900),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1890),
.B(n_262),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1891),
.B(n_263),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1848),
.B(n_263),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1903),
.B(n_264),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_1907),
.B(n_264),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1686),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_1722),
.B(n_265),
.Y(n_2170)
);

AND2x2_ASAP7_75t_SL g2171 ( 
.A(n_1959),
.B(n_1827),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_1685),
.B(n_266),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1664),
.B(n_267),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1847),
.Y(n_2174)
);

HB1xp67_ASAP7_75t_L g2175 ( 
.A(n_1845),
.Y(n_2175)
);

NOR2xp67_ASAP7_75t_L g2176 ( 
.A(n_1757),
.B(n_382),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1840),
.B(n_268),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1915),
.B(n_268),
.Y(n_2178)
);

INVx3_ASAP7_75t_L g2179 ( 
.A(n_1781),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_1735),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_1916),
.B(n_269),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1738),
.Y(n_2182)
);

NOR2xp33_ASAP7_75t_L g2183 ( 
.A(n_1917),
.B(n_269),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1714),
.B(n_271),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1785),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1943),
.B(n_271),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1835),
.B(n_272),
.Y(n_2187)
);

AND2x6_ASAP7_75t_L g2188 ( 
.A(n_1872),
.B(n_1884),
.Y(n_2188)
);

NAND2x1p5_ASAP7_75t_L g2189 ( 
.A(n_1849),
.B(n_272),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1845),
.B(n_273),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1787),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1941),
.B(n_273),
.Y(n_2192)
);

OAI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_1699),
.A2(n_389),
.B(n_388),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_L g2194 ( 
.A(n_1868),
.B(n_1851),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_1936),
.B(n_274),
.Y(n_2195)
);

INVx3_ASAP7_75t_L g2196 ( 
.A(n_1788),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1815),
.B(n_275),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_1886),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_1852),
.B(n_276),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_1789),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1652),
.B(n_1658),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1833),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1937),
.B(n_277),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_1790),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1882),
.B(n_277),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_1901),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_1791),
.Y(n_2207)
);

INVx4_ASAP7_75t_L g2208 ( 
.A(n_1922),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1834),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_1713),
.B(n_1762),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_1889),
.B(n_279),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_1861),
.B(n_279),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_1864),
.B(n_280),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1661),
.B(n_280),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_1717),
.B(n_281),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_1862),
.B(n_281),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1795),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_L g2218 ( 
.A(n_1945),
.B(n_283),
.Y(n_2218)
);

NOR2xp33_ASAP7_75t_L g2219 ( 
.A(n_2065),
.B(n_1919),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1997),
.B(n_1970),
.Y(n_2220)
);

INVx3_ASAP7_75t_L g2221 ( 
.A(n_2006),
.Y(n_2221)
);

BUFx6f_ASAP7_75t_L g2222 ( 
.A(n_2022),
.Y(n_2222)
);

INVxp67_ASAP7_75t_L g2223 ( 
.A(n_1981),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2060),
.B(n_1972),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_2006),
.B(n_1832),
.Y(n_2225)
);

INVx2_ASAP7_75t_SL g2226 ( 
.A(n_2022),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2155),
.Y(n_2227)
);

BUFx12f_ASAP7_75t_L g2228 ( 
.A(n_2012),
.Y(n_2228)
);

BUFx6f_ASAP7_75t_L g2229 ( 
.A(n_2012),
.Y(n_2229)
);

AND2x6_ASAP7_75t_L g2230 ( 
.A(n_2086),
.B(n_1887),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1973),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1986),
.B(n_1946),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2171),
.B(n_1651),
.Y(n_2233)
);

CKINVDCx20_ASAP7_75t_R g2234 ( 
.A(n_1979),
.Y(n_2234)
);

AND2x4_ASAP7_75t_L g2235 ( 
.A(n_2111),
.B(n_1892),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2163),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2145),
.B(n_1951),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_2101),
.B(n_1952),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2202),
.Y(n_2239)
);

INVx1_ASAP7_75t_SL g2240 ( 
.A(n_2050),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2026),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2028),
.B(n_1955),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2103),
.B(n_2157),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2019),
.B(n_1956),
.Y(n_2244)
);

OR2x6_ASAP7_75t_L g2245 ( 
.A(n_2031),
.B(n_1901),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_2031),
.B(n_1858),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_2034),
.B(n_1728),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_L g2248 ( 
.A(n_1998),
.B(n_2092),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_2064),
.Y(n_2249)
);

AND2x4_ASAP7_75t_L g2250 ( 
.A(n_2034),
.B(n_1942),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2202),
.Y(n_2251)
);

BUFx2_ASAP7_75t_L g2252 ( 
.A(n_2061),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2078),
.B(n_1958),
.Y(n_2253)
);

INVx2_ASAP7_75t_SL g2254 ( 
.A(n_1994),
.Y(n_2254)
);

BUFx6f_ASAP7_75t_L g2255 ( 
.A(n_2064),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2133),
.B(n_1961),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1985),
.B(n_1962),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2209),
.Y(n_2258)
);

BUFx3_ASAP7_75t_L g2259 ( 
.A(n_2064),
.Y(n_2259)
);

NAND2x1_ASAP7_75t_SL g2260 ( 
.A(n_2172),
.B(n_1932),
.Y(n_2260)
);

HB1xp67_ASAP7_75t_L g2261 ( 
.A(n_2027),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2209),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2038),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_2061),
.B(n_1836),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2148),
.B(n_1773),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2002),
.B(n_1880),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2174),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2077),
.B(n_1963),
.Y(n_2268)
);

INVx3_ASAP7_75t_SL g2269 ( 
.A(n_1993),
.Y(n_2269)
);

NOR2xp67_ASAP7_75t_L g2270 ( 
.A(n_2035),
.B(n_1909),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2014),
.B(n_2018),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2174),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1975),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1975),
.Y(n_2274)
);

INVx5_ASAP7_75t_L g2275 ( 
.A(n_1987),
.Y(n_2275)
);

NOR2x1p5_ASAP7_75t_L g2276 ( 
.A(n_1989),
.B(n_1929),
.Y(n_2276)
);

BUFx2_ASAP7_75t_L g2277 ( 
.A(n_2036),
.Y(n_2277)
);

BUFx2_ASAP7_75t_L g2278 ( 
.A(n_2087),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2042),
.Y(n_2279)
);

AND2x2_ASAP7_75t_SL g2280 ( 
.A(n_2131),
.B(n_1974),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2112),
.B(n_1964),
.Y(n_2281)
);

NOR2xp33_ASAP7_75t_SL g2282 ( 
.A(n_2063),
.B(n_1830),
.Y(n_2282)
);

NAND2x1p5_ASAP7_75t_L g2283 ( 
.A(n_2037),
.B(n_2024),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2079),
.B(n_1904),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2054),
.B(n_2020),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_2084),
.B(n_1842),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_1977),
.Y(n_2287)
);

BUFx3_ASAP7_75t_L g2288 ( 
.A(n_2136),
.Y(n_2288)
);

AND2x6_ASAP7_75t_L g2289 ( 
.A(n_2086),
.B(n_1968),
.Y(n_2289)
);

NAND2xp33_ASAP7_75t_L g2290 ( 
.A(n_2201),
.B(n_1922),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_1977),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2054),
.B(n_1950),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_2175),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2218),
.B(n_1966),
.Y(n_2294)
);

CKINVDCx11_ASAP7_75t_R g2295 ( 
.A(n_2057),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2051),
.Y(n_2296)
);

OR2x2_ASAP7_75t_L g2297 ( 
.A(n_2083),
.B(n_1700),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2052),
.Y(n_2298)
);

BUFx6f_ASAP7_75t_L g2299 ( 
.A(n_1977),
.Y(n_2299)
);

NAND2x1p5_ASAP7_75t_L g2300 ( 
.A(n_2037),
.B(n_1749),
.Y(n_2300)
);

NAND2x1p5_ASAP7_75t_L g2301 ( 
.A(n_2037),
.B(n_1819),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2003),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_1980),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2003),
.Y(n_2304)
);

NAND2x1p5_ASAP7_75t_L g2305 ( 
.A(n_1989),
.B(n_1797),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2068),
.B(n_1948),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2056),
.Y(n_2307)
);

NAND2x1p5_ASAP7_75t_L g2308 ( 
.A(n_2043),
.B(n_1798),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2058),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2009),
.B(n_2015),
.Y(n_2310)
);

AND2x4_ASAP7_75t_L g2311 ( 
.A(n_2048),
.B(n_1925),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2104),
.B(n_1865),
.Y(n_2312)
);

OR2x6_ASAP7_75t_L g2313 ( 
.A(n_2057),
.B(n_1969),
.Y(n_2313)
);

INVxp67_ASAP7_75t_L g2314 ( 
.A(n_2194),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2009),
.Y(n_2315)
);

BUFx3_ASAP7_75t_L g2316 ( 
.A(n_2160),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2015),
.B(n_2030),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2030),
.B(n_1953),
.Y(n_2318)
);

NAND2x1p5_ASAP7_75t_L g2319 ( 
.A(n_2205),
.B(n_1799),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2186),
.B(n_1935),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2033),
.B(n_2041),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2159),
.B(n_1913),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2033),
.B(n_1875),
.Y(n_2323)
);

INVx1_ASAP7_75t_SL g2324 ( 
.A(n_2013),
.Y(n_2324)
);

BUFx6f_ASAP7_75t_L g2325 ( 
.A(n_1980),
.Y(n_2325)
);

INVx3_ASAP7_75t_L g2326 ( 
.A(n_1980),
.Y(n_2326)
);

BUFx4f_ASAP7_75t_L g2327 ( 
.A(n_1996),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2041),
.Y(n_2328)
);

CKINVDCx8_ASAP7_75t_R g2329 ( 
.A(n_2149),
.Y(n_2329)
);

BUFx2_ASAP7_75t_L g2330 ( 
.A(n_2039),
.Y(n_2330)
);

BUFx12f_ASAP7_75t_L g2331 ( 
.A(n_1984),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2046),
.Y(n_2332)
);

INVx2_ASAP7_75t_SL g2333 ( 
.A(n_2124),
.Y(n_2333)
);

NOR2x1_ASAP7_75t_L g2334 ( 
.A(n_2142),
.B(n_1905),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2046),
.B(n_1828),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2100),
.B(n_1866),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_2023),
.Y(n_2337)
);

NAND2x1p5_ASAP7_75t_L g2338 ( 
.A(n_2205),
.B(n_2211),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_2161),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2053),
.B(n_1922),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2067),
.Y(n_2341)
);

INVx3_ASAP7_75t_L g2342 ( 
.A(n_2023),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2053),
.B(n_1920),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2080),
.B(n_1902),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2071),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_2091),
.B(n_1801),
.Y(n_2346)
);

INVx1_ASAP7_75t_SL g2347 ( 
.A(n_2039),
.Y(n_2347)
);

INVxp67_ASAP7_75t_L g2348 ( 
.A(n_2181),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_1983),
.B(n_2089),
.Y(n_2349)
);

INVx5_ASAP7_75t_L g2350 ( 
.A(n_1996),
.Y(n_2350)
);

INVx6_ASAP7_75t_L g2351 ( 
.A(n_2023),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2073),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_2004),
.B(n_1804),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2121),
.B(n_1663),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_2198),
.B(n_1805),
.Y(n_2355)
);

HB1xp67_ASAP7_75t_L g2356 ( 
.A(n_2130),
.Y(n_2356)
);

CKINVDCx8_ASAP7_75t_R g2357 ( 
.A(n_2049),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2129),
.B(n_1669),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_2025),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2070),
.B(n_1727),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2070),
.Y(n_2361)
);

BUFx8_ASAP7_75t_SL g2362 ( 
.A(n_2124),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2100),
.B(n_1727),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2100),
.B(n_1727),
.Y(n_2364)
);

AND2x4_ASAP7_75t_L g2365 ( 
.A(n_2206),
.B(n_1806),
.Y(n_2365)
);

BUFx2_ASAP7_75t_L g2366 ( 
.A(n_2049),
.Y(n_2366)
);

OR2x2_ASAP7_75t_L g2367 ( 
.A(n_2210),
.B(n_1676),
.Y(n_2367)
);

HB1xp67_ASAP7_75t_L g2368 ( 
.A(n_2130),
.Y(n_2368)
);

BUFx4f_ASAP7_75t_L g2369 ( 
.A(n_2110),
.Y(n_2369)
);

OR2x6_ASAP7_75t_L g2370 ( 
.A(n_2139),
.B(n_1839),
.Y(n_2370)
);

BUFx8_ASAP7_75t_SL g2371 ( 
.A(n_2047),
.Y(n_2371)
);

INVx3_ASAP7_75t_L g2372 ( 
.A(n_2025),
.Y(n_2372)
);

NAND2x1p5_ASAP7_75t_L g2373 ( 
.A(n_2211),
.B(n_1809),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_2115),
.Y(n_2374)
);

INVxp67_ASAP7_75t_SL g2375 ( 
.A(n_2139),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1995),
.B(n_1727),
.Y(n_2376)
);

INVxp67_ASAP7_75t_L g2377 ( 
.A(n_2183),
.Y(n_2377)
);

INVxp67_ASAP7_75t_L g2378 ( 
.A(n_2109),
.Y(n_2378)
);

INVx6_ASAP7_75t_SL g2379 ( 
.A(n_2245),
.Y(n_2379)
);

BUFx4_ASAP7_75t_SL g2380 ( 
.A(n_2234),
.Y(n_2380)
);

INVx2_ASAP7_75t_SL g2381 ( 
.A(n_2288),
.Y(n_2381)
);

INVx3_ASAP7_75t_L g2382 ( 
.A(n_2228),
.Y(n_2382)
);

INVx2_ASAP7_75t_SL g2383 ( 
.A(n_2275),
.Y(n_2383)
);

INVx1_ASAP7_75t_SL g2384 ( 
.A(n_2339),
.Y(n_2384)
);

INVx3_ASAP7_75t_L g2385 ( 
.A(n_2222),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2239),
.Y(n_2386)
);

BUFx6f_ASAP7_75t_L g2387 ( 
.A(n_2222),
.Y(n_2387)
);

BUFx3_ASAP7_75t_L g2388 ( 
.A(n_2316),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2251),
.Y(n_2389)
);

INVxp67_ASAP7_75t_SL g2390 ( 
.A(n_2375),
.Y(n_2390)
);

INVx2_ASAP7_75t_SL g2391 ( 
.A(n_2275),
.Y(n_2391)
);

OR2x2_ASAP7_75t_L g2392 ( 
.A(n_2367),
.B(n_2000),
.Y(n_2392)
);

INVx5_ASAP7_75t_SL g2393 ( 
.A(n_2245),
.Y(n_2393)
);

OAI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2294),
.A2(n_2128),
.B1(n_2093),
.B2(n_2190),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_2366),
.B(n_2140),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2258),
.Y(n_2396)
);

OR2x2_ASAP7_75t_L g2397 ( 
.A(n_2219),
.B(n_2266),
.Y(n_2397)
);

BUFx6f_ASAP7_75t_L g2398 ( 
.A(n_2229),
.Y(n_2398)
);

INVx4_ASAP7_75t_L g2399 ( 
.A(n_2269),
.Y(n_2399)
);

INVx6_ASAP7_75t_SL g2400 ( 
.A(n_2370),
.Y(n_2400)
);

BUFx3_ASAP7_75t_L g2401 ( 
.A(n_2362),
.Y(n_2401)
);

NOR2xp67_ASAP7_75t_SL g2402 ( 
.A(n_2357),
.B(n_2142),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2262),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2280),
.B(n_2138),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2241),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2263),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_2333),
.B(n_2140),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_2329),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2267),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2272),
.Y(n_2410)
);

INVx2_ASAP7_75t_SL g2411 ( 
.A(n_2327),
.Y(n_2411)
);

INVxp67_ASAP7_75t_SL g2412 ( 
.A(n_2338),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2279),
.Y(n_2413)
);

BUFx12f_ASAP7_75t_L g2414 ( 
.A(n_2295),
.Y(n_2414)
);

BUFx4f_ASAP7_75t_SL g2415 ( 
.A(n_2331),
.Y(n_2415)
);

BUFx12f_ASAP7_75t_L g2416 ( 
.A(n_2374),
.Y(n_2416)
);

INVxp67_ASAP7_75t_L g2417 ( 
.A(n_2293),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2296),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2298),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2273),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2307),
.Y(n_2421)
);

INVx4_ASAP7_75t_L g2422 ( 
.A(n_2229),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2224),
.B(n_2126),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2278),
.Y(n_2424)
);

BUFx2_ASAP7_75t_L g2425 ( 
.A(n_2277),
.Y(n_2425)
);

INVx4_ASAP7_75t_L g2426 ( 
.A(n_2350),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2274),
.Y(n_2427)
);

BUFx2_ASAP7_75t_L g2428 ( 
.A(n_2330),
.Y(n_2428)
);

INVx1_ASAP7_75t_SL g2429 ( 
.A(n_2240),
.Y(n_2429)
);

HB1xp67_ASAP7_75t_L g2430 ( 
.A(n_2261),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_2350),
.B(n_2212),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2309),
.Y(n_2432)
);

AOI22xp33_ASAP7_75t_SL g2433 ( 
.A1(n_2344),
.A2(n_2127),
.B1(n_2107),
.B2(n_2105),
.Y(n_2433)
);

BUFx3_ASAP7_75t_L g2434 ( 
.A(n_2259),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2302),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_2249),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_2249),
.Y(n_2437)
);

BUFx12f_ASAP7_75t_L g2438 ( 
.A(n_2247),
.Y(n_2438)
);

AND2x4_ASAP7_75t_L g2439 ( 
.A(n_2264),
.B(n_2212),
.Y(n_2439)
);

INVx6_ASAP7_75t_SL g2440 ( 
.A(n_2370),
.Y(n_2440)
);

BUFx12f_ASAP7_75t_L g2441 ( 
.A(n_2254),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2233),
.A2(n_1687),
.B1(n_1739),
.B2(n_2177),
.Y(n_2442)
);

INVx2_ASAP7_75t_SL g2443 ( 
.A(n_2255),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2304),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2315),
.Y(n_2445)
);

INVx2_ASAP7_75t_SL g2446 ( 
.A(n_2255),
.Y(n_2446)
);

CKINVDCx20_ASAP7_75t_R g2447 ( 
.A(n_2324),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2224),
.B(n_2162),
.Y(n_2448)
);

OAI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2248),
.A2(n_2090),
.B1(n_2096),
.B2(n_2132),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2341),
.Y(n_2450)
);

NAND2x1p5_ASAP7_75t_L g2451 ( 
.A(n_2226),
.B(n_2025),
.Y(n_2451)
);

OAI22xp5_ASAP7_75t_SL g2452 ( 
.A1(n_2314),
.A2(n_1734),
.B1(n_1879),
.B2(n_1838),
.Y(n_2452)
);

NAND2x1p5_ASAP7_75t_L g2453 ( 
.A(n_2221),
.B(n_2011),
.Y(n_2453)
);

INVx1_ASAP7_75t_SL g2454 ( 
.A(n_2347),
.Y(n_2454)
);

INVx1_ASAP7_75t_SL g2455 ( 
.A(n_2297),
.Y(n_2455)
);

AOI22xp33_ASAP7_75t_L g2456 ( 
.A1(n_2265),
.A2(n_2114),
.B1(n_2108),
.B2(n_2049),
.Y(n_2456)
);

BUFx3_ASAP7_75t_L g2457 ( 
.A(n_2235),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2225),
.Y(n_2458)
);

BUFx6f_ASAP7_75t_L g2459 ( 
.A(n_2287),
.Y(n_2459)
);

BUFx2_ASAP7_75t_L g2460 ( 
.A(n_2356),
.Y(n_2460)
);

BUFx3_ASAP7_75t_L g2461 ( 
.A(n_2355),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2287),
.Y(n_2462)
);

INVx8_ASAP7_75t_L g2463 ( 
.A(n_2289),
.Y(n_2463)
);

BUFx3_ASAP7_75t_L g2464 ( 
.A(n_2365),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2328),
.Y(n_2465)
);

BUFx12f_ASAP7_75t_L g2466 ( 
.A(n_2311),
.Y(n_2466)
);

BUFx2_ASAP7_75t_L g2467 ( 
.A(n_2368),
.Y(n_2467)
);

BUFx2_ASAP7_75t_R g2468 ( 
.A(n_2371),
.Y(n_2468)
);

AND2x4_ASAP7_75t_L g2469 ( 
.A(n_2276),
.B(n_2182),
.Y(n_2469)
);

INVx2_ASAP7_75t_SL g2470 ( 
.A(n_2369),
.Y(n_2470)
);

INVx4_ASAP7_75t_L g2471 ( 
.A(n_2291),
.Y(n_2471)
);

AND2x4_ASAP7_75t_L g2472 ( 
.A(n_2253),
.B(n_2208),
.Y(n_2472)
);

BUFx3_ASAP7_75t_L g2473 ( 
.A(n_2283),
.Y(n_2473)
);

BUFx3_ASAP7_75t_L g2474 ( 
.A(n_2346),
.Y(n_2474)
);

BUFx3_ASAP7_75t_L g2475 ( 
.A(n_2353),
.Y(n_2475)
);

INVx6_ASAP7_75t_L g2476 ( 
.A(n_2246),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2349),
.B(n_2049),
.Y(n_2477)
);

INVx5_ASAP7_75t_L g2478 ( 
.A(n_2289),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2271),
.B(n_1982),
.Y(n_2479)
);

BUFx10_ASAP7_75t_L g2480 ( 
.A(n_2381),
.Y(n_2480)
);

INVx6_ASAP7_75t_L g2481 ( 
.A(n_2416),
.Y(n_2481)
);

INVxp67_ASAP7_75t_SL g2482 ( 
.A(n_2390),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2386),
.Y(n_2483)
);

AOI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2433),
.A2(n_2442),
.B1(n_2452),
.B2(n_2423),
.Y(n_2484)
);

AOI22xp33_ASAP7_75t_SL g2485 ( 
.A1(n_2404),
.A2(n_1769),
.B1(n_2320),
.B2(n_2322),
.Y(n_2485)
);

BUFx10_ASAP7_75t_L g2486 ( 
.A(n_2411),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2389),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2405),
.Y(n_2488)
);

INVx1_ASAP7_75t_SL g2489 ( 
.A(n_2447),
.Y(n_2489)
);

INVx1_ASAP7_75t_SL g2490 ( 
.A(n_2380),
.Y(n_2490)
);

HB1xp67_ASAP7_75t_L g2491 ( 
.A(n_2424),
.Y(n_2491)
);

AND2x4_ASAP7_75t_SL g2492 ( 
.A(n_2399),
.B(n_2291),
.Y(n_2492)
);

AOI22xp33_ASAP7_75t_L g2493 ( 
.A1(n_2449),
.A2(n_2320),
.B1(n_2322),
.B2(n_2166),
.Y(n_2493)
);

NAND2x1p5_ASAP7_75t_L g2494 ( 
.A(n_2478),
.B(n_2252),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2403),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2406),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2409),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2435),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2465),
.Y(n_2499)
);

CKINVDCx11_ASAP7_75t_R g2500 ( 
.A(n_2414),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2396),
.Y(n_2501)
);

INVx4_ASAP7_75t_L g2502 ( 
.A(n_2415),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2396),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2410),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2410),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2413),
.Y(n_2506)
);

BUFx6f_ASAP7_75t_L g2507 ( 
.A(n_2463),
.Y(n_2507)
);

INVxp67_ASAP7_75t_L g2508 ( 
.A(n_2424),
.Y(n_2508)
);

BUFx10_ASAP7_75t_L g2509 ( 
.A(n_2431),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2420),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2420),
.Y(n_2511)
);

AOI22xp33_ASAP7_75t_L g2512 ( 
.A1(n_2448),
.A2(n_2150),
.B1(n_2358),
.B2(n_2354),
.Y(n_2512)
);

OAI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2394),
.A2(n_2348),
.B1(n_2377),
.B2(n_2378),
.Y(n_2513)
);

INVx1_ASAP7_75t_SL g2514 ( 
.A(n_2429),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2427),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2397),
.A2(n_1926),
.B1(n_1938),
.B2(n_1949),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2418),
.Y(n_2517)
);

INVxp67_ASAP7_75t_SL g2518 ( 
.A(n_2417),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2477),
.A2(n_2187),
.B1(n_2192),
.B2(n_1854),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2479),
.B(n_2244),
.Y(n_2520)
);

AOI22xp33_ASAP7_75t_L g2521 ( 
.A1(n_2456),
.A2(n_2117),
.B1(n_2123),
.B2(n_2120),
.Y(n_2521)
);

INVx1_ASAP7_75t_SL g2522 ( 
.A(n_2384),
.Y(n_2522)
);

BUFx3_ASAP7_75t_L g2523 ( 
.A(n_2388),
.Y(n_2523)
);

BUFx2_ASAP7_75t_L g2524 ( 
.A(n_2474),
.Y(n_2524)
);

OAI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2425),
.A2(n_2243),
.B1(n_2317),
.B2(n_2310),
.Y(n_2525)
);

INVx1_ASAP7_75t_SL g2526 ( 
.A(n_2425),
.Y(n_2526)
);

AOI22xp33_ASAP7_75t_L g2527 ( 
.A1(n_2392),
.A2(n_2284),
.B1(n_2001),
.B2(n_2230),
.Y(n_2527)
);

INVx6_ASAP7_75t_L g2528 ( 
.A(n_2441),
.Y(n_2528)
);

CKINVDCx6p67_ASAP7_75t_R g2529 ( 
.A(n_2401),
.Y(n_2529)
);

INVx2_ASAP7_75t_SL g2530 ( 
.A(n_2476),
.Y(n_2530)
);

AOI22xp33_ASAP7_75t_L g2531 ( 
.A1(n_2466),
.A2(n_2230),
.B1(n_2306),
.B2(n_2178),
.Y(n_2531)
);

BUFx12f_ASAP7_75t_L g2532 ( 
.A(n_2438),
.Y(n_2532)
);

BUFx6f_ASAP7_75t_L g2533 ( 
.A(n_2463),
.Y(n_2533)
);

OAI22xp5_ASAP7_75t_L g2534 ( 
.A1(n_2430),
.A2(n_2321),
.B1(n_2292),
.B2(n_2335),
.Y(n_2534)
);

BUFx4f_ASAP7_75t_SL g2535 ( 
.A(n_2379),
.Y(n_2535)
);

AOI22xp33_ASAP7_75t_SL g2536 ( 
.A1(n_2455),
.A2(n_2075),
.B1(n_2040),
.B2(n_2289),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2439),
.B(n_2242),
.Y(n_2537)
);

BUFx12f_ASAP7_75t_L g2538 ( 
.A(n_2426),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2454),
.B(n_2232),
.Y(n_2539)
);

AOI22xp5_ASAP7_75t_L g2540 ( 
.A1(n_2472),
.A2(n_1960),
.B1(n_2242),
.B2(n_2223),
.Y(n_2540)
);

CKINVDCx20_ASAP7_75t_R g2541 ( 
.A(n_2434),
.Y(n_2541)
);

BUFx3_ASAP7_75t_L g2542 ( 
.A(n_2461),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2427),
.Y(n_2543)
);

NAND2x1p5_ASAP7_75t_L g2544 ( 
.A(n_2478),
.B(n_2299),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2444),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2419),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2421),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_2478),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2444),
.Y(n_2549)
);

OR2x2_ASAP7_75t_L g2550 ( 
.A(n_2428),
.B(n_2268),
.Y(n_2550)
);

OAI22xp5_ASAP7_75t_L g2551 ( 
.A1(n_2445),
.A2(n_2285),
.B1(n_2214),
.B2(n_2102),
.Y(n_2551)
);

OAI21xp33_ASAP7_75t_L g2552 ( 
.A1(n_2445),
.A2(n_2184),
.B(n_2173),
.Y(n_2552)
);

BUFx2_ASAP7_75t_SL g2553 ( 
.A(n_2469),
.Y(n_2553)
);

AOI22xp5_ASAP7_75t_L g2554 ( 
.A1(n_2472),
.A2(n_2313),
.B1(n_2282),
.B2(n_2290),
.Y(n_2554)
);

NAND2x1p5_ASAP7_75t_L g2555 ( 
.A(n_2402),
.B(n_2299),
.Y(n_2555)
);

AOI22xp33_ASAP7_75t_L g2556 ( 
.A1(n_2475),
.A2(n_2230),
.B1(n_1957),
.B2(n_1934),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2439),
.B(n_2237),
.Y(n_2557)
);

AOI21xp33_ASAP7_75t_L g2558 ( 
.A1(n_2432),
.A2(n_2122),
.B(n_2197),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2489),
.B(n_2522),
.Y(n_2559)
);

OAI21xp5_ASAP7_75t_SL g2560 ( 
.A1(n_2493),
.A2(n_1774),
.B(n_2074),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2488),
.Y(n_2561)
);

AOI22xp33_ASAP7_75t_SL g2562 ( 
.A1(n_2525),
.A2(n_2208),
.B1(n_1841),
.B2(n_2313),
.Y(n_2562)
);

AOI22xp33_ASAP7_75t_L g2563 ( 
.A1(n_2516),
.A2(n_1841),
.B1(n_2352),
.B2(n_2345),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2557),
.B(n_2428),
.Y(n_2564)
);

OR2x2_ASAP7_75t_SL g2565 ( 
.A(n_2481),
.B(n_2312),
.Y(n_2565)
);

OAI21xp33_ASAP7_75t_L g2566 ( 
.A1(n_2552),
.A2(n_2551),
.B(n_2513),
.Y(n_2566)
);

OAI222xp33_ASAP7_75t_L g2567 ( 
.A1(n_2485),
.A2(n_2373),
.B1(n_2319),
.B2(n_2257),
.C1(n_2281),
.C2(n_2256),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2496),
.Y(n_2568)
);

AOI22xp33_ASAP7_75t_SL g2569 ( 
.A1(n_2534),
.A2(n_1841),
.B1(n_2032),
.B2(n_1976),
.Y(n_2569)
);

OAI22xp33_ASAP7_75t_L g2570 ( 
.A1(n_2519),
.A2(n_2189),
.B1(n_2318),
.B2(n_2153),
.Y(n_2570)
);

HB1xp67_ASAP7_75t_L g2571 ( 
.A(n_2491),
.Y(n_2571)
);

BUFx4f_ASAP7_75t_SL g2572 ( 
.A(n_2541),
.Y(n_2572)
);

INVx1_ASAP7_75t_SL g2573 ( 
.A(n_2514),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2506),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2483),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2537),
.B(n_2460),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2540),
.B(n_2460),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_L g2578 ( 
.A1(n_2484),
.A2(n_1841),
.B1(n_2450),
.B2(n_2231),
.Y(n_2578)
);

OAI21xp5_ASAP7_75t_SL g2579 ( 
.A1(n_2521),
.A2(n_2193),
.B(n_2170),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2517),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2556),
.A2(n_2180),
.B1(n_2440),
.B2(n_2400),
.Y(n_2581)
);

AOI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_2512),
.A2(n_2395),
.B1(n_2220),
.B2(n_2199),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_2500),
.Y(n_2583)
);

BUFx12f_ASAP7_75t_L g2584 ( 
.A(n_2502),
.Y(n_2584)
);

OAI22xp5_ASAP7_75t_L g2585 ( 
.A1(n_2526),
.A2(n_2508),
.B1(n_2518),
.B2(n_2531),
.Y(n_2585)
);

OAI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_2482),
.A2(n_2270),
.B(n_2340),
.Y(n_2586)
);

BUFx3_ASAP7_75t_L g2587 ( 
.A(n_2523),
.Y(n_2587)
);

OAI21xp33_ASAP7_75t_L g2588 ( 
.A1(n_2558),
.A2(n_2260),
.B(n_2095),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2487),
.Y(n_2589)
);

OAI21xp5_ASAP7_75t_SL g2590 ( 
.A1(n_2554),
.A2(n_2301),
.B(n_2300),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2550),
.B(n_2467),
.Y(n_2591)
);

BUFx2_ASAP7_75t_L g2592 ( 
.A(n_2524),
.Y(n_2592)
);

INVx6_ASAP7_75t_L g2593 ( 
.A(n_2502),
.Y(n_2593)
);

AOI22xp33_ASAP7_75t_L g2594 ( 
.A1(n_2527),
.A2(n_2536),
.B1(n_2520),
.B2(n_2180),
.Y(n_2594)
);

AOI22xp33_ASAP7_75t_L g2595 ( 
.A1(n_2546),
.A2(n_2180),
.B1(n_2440),
.B2(n_2400),
.Y(n_2595)
);

OAI22xp5_ASAP7_75t_L g2596 ( 
.A1(n_2501),
.A2(n_2332),
.B1(n_2361),
.B2(n_2125),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_2547),
.A2(n_2250),
.B1(n_2395),
.B2(n_2044),
.Y(n_2597)
);

INVx2_ASAP7_75t_SL g2598 ( 
.A(n_2492),
.Y(n_2598)
);

CKINVDCx14_ASAP7_75t_R g2599 ( 
.A(n_2529),
.Y(n_2599)
);

OAI21xp33_ASAP7_75t_L g2600 ( 
.A1(n_2503),
.A2(n_2098),
.B(n_2097),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2495),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2490),
.B(n_2470),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2539),
.B(n_2467),
.Y(n_2603)
);

OAI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2504),
.A2(n_2106),
.B1(n_2323),
.B2(n_2360),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2553),
.B(n_2021),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2497),
.Y(n_2606)
);

NOR2xp33_ASAP7_75t_L g2607 ( 
.A(n_2535),
.B(n_2408),
.Y(n_2607)
);

OAI21xp33_ASAP7_75t_L g2608 ( 
.A1(n_2505),
.A2(n_2118),
.B(n_2113),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2498),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_SL g2610 ( 
.A1(n_2553),
.A2(n_2216),
.B1(n_2029),
.B2(n_2045),
.Y(n_2610)
);

OAI22xp5_ASAP7_75t_L g2611 ( 
.A1(n_2510),
.A2(n_2376),
.B1(n_2017),
.B2(n_2165),
.Y(n_2611)
);

INVx6_ASAP7_75t_L g2612 ( 
.A(n_2532),
.Y(n_2612)
);

OAI21xp5_ASAP7_75t_SL g2613 ( 
.A1(n_2494),
.A2(n_2151),
.B(n_2146),
.Y(n_2613)
);

AOI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_2542),
.A2(n_2286),
.B1(n_2469),
.B2(n_2457),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2499),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2530),
.B(n_2237),
.Y(n_2616)
);

BUFx6f_ASAP7_75t_L g2617 ( 
.A(n_2507),
.Y(n_2617)
);

AOI22xp5_ASAP7_75t_L g2618 ( 
.A1(n_2511),
.A2(n_2431),
.B1(n_2402),
.B2(n_2407),
.Y(n_2618)
);

AOI22xp33_ASAP7_75t_L g2619 ( 
.A1(n_2515),
.A2(n_2094),
.B1(n_2135),
.B2(n_2081),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2543),
.B(n_2545),
.Y(n_2620)
);

OAI22xp5_ASAP7_75t_SL g2621 ( 
.A1(n_2481),
.A2(n_2164),
.B1(n_2059),
.B2(n_2066),
.Y(n_2621)
);

OAI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_2549),
.A2(n_2383),
.B1(n_2391),
.B2(n_2141),
.Y(n_2622)
);

CKINVDCx6p67_ASAP7_75t_R g2623 ( 
.A(n_2538),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_L g2624 ( 
.A1(n_2507),
.A2(n_2191),
.B1(n_2217),
.B2(n_2143),
.Y(n_2624)
);

OAI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2555),
.A2(n_2238),
.B1(n_2364),
.B2(n_2363),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2509),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2548),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2509),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2548),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2544),
.Y(n_2630)
);

HB1xp67_ASAP7_75t_L g2631 ( 
.A(n_2507),
.Y(n_2631)
);

OAI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2528),
.A2(n_1682),
.B1(n_1671),
.B2(n_2305),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2533),
.Y(n_2633)
);

AOI22xp33_ASAP7_75t_SL g2634 ( 
.A1(n_2528),
.A2(n_2393),
.B1(n_1990),
.B2(n_2007),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2533),
.A2(n_2393),
.B1(n_2069),
.B2(n_2076),
.Y(n_2635)
);

AOI22xp33_ASAP7_75t_L g2636 ( 
.A1(n_2621),
.A2(n_2204),
.B1(n_2343),
.B2(n_2062),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2603),
.B(n_2055),
.Y(n_2637)
);

NAND3xp33_ASAP7_75t_L g2638 ( 
.A(n_2566),
.B(n_2158),
.C(n_1999),
.Y(n_2638)
);

AOI22xp33_ASAP7_75t_SL g2639 ( 
.A1(n_2621),
.A2(n_2168),
.B1(n_2167),
.B2(n_2088),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2591),
.B(n_2436),
.Y(n_2640)
);

AOI22xp33_ASAP7_75t_L g2641 ( 
.A1(n_2578),
.A2(n_2204),
.B1(n_2336),
.B2(n_2207),
.Y(n_2641)
);

NAND2xp33_ASAP7_75t_SL g2642 ( 
.A(n_2583),
.B(n_2533),
.Y(n_2642)
);

AOI22xp33_ASAP7_75t_L g2643 ( 
.A1(n_2566),
.A2(n_2204),
.B1(n_2334),
.B2(n_2464),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2579),
.A2(n_2468),
.B1(n_2476),
.B2(n_2453),
.Y(n_2644)
);

OAI21xp5_ASAP7_75t_SL g2645 ( 
.A1(n_2613),
.A2(n_2215),
.B(n_2203),
.Y(n_2645)
);

AOI22xp33_ASAP7_75t_L g2646 ( 
.A1(n_2563),
.A2(n_2185),
.B1(n_1978),
.B2(n_2407),
.Y(n_2646)
);

AOI22xp33_ASAP7_75t_L g2647 ( 
.A1(n_2594),
.A2(n_1978),
.B1(n_2144),
.B2(n_2137),
.Y(n_2647)
);

AOI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_2569),
.A2(n_2588),
.B1(n_2581),
.B2(n_2610),
.Y(n_2648)
);

INVxp67_ASAP7_75t_L g2649 ( 
.A(n_2559),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2588),
.A2(n_2152),
.B1(n_2154),
.B2(n_2253),
.Y(n_2650)
);

OAI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2560),
.A2(n_2379),
.B1(n_2412),
.B2(n_2308),
.Y(n_2651)
);

AOI22xp33_ASAP7_75t_SL g2652 ( 
.A1(n_2577),
.A2(n_2195),
.B1(n_2213),
.B2(n_2458),
.Y(n_2652)
);

AOI22xp33_ASAP7_75t_L g2653 ( 
.A1(n_2608),
.A2(n_2188),
.B1(n_2072),
.B2(n_2085),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2576),
.B(n_2436),
.Y(n_2654)
);

AOI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2562),
.A2(n_2119),
.B1(n_2188),
.B2(n_2227),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2608),
.A2(n_2188),
.B1(n_2072),
.B2(n_1992),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2575),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2570),
.A2(n_2188),
.B1(n_2072),
.B2(n_2008),
.Y(n_2658)
);

AOI22xp33_ASAP7_75t_SL g2659 ( 
.A1(n_2632),
.A2(n_2134),
.B1(n_2196),
.B2(n_2179),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2582),
.A2(n_2634),
.B1(n_2597),
.B2(n_2635),
.Y(n_2660)
);

OA21x2_ASAP7_75t_L g2661 ( 
.A1(n_2600),
.A2(n_1758),
.B(n_1853),
.Y(n_2661)
);

OAI21xp5_ASAP7_75t_SL g2662 ( 
.A1(n_2567),
.A2(n_2382),
.B(n_2451),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2564),
.B(n_2437),
.Y(n_2663)
);

AO22x1_ASAP7_75t_L g2664 ( 
.A1(n_2626),
.A2(n_2628),
.B1(n_2573),
.B2(n_2633),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2589),
.Y(n_2665)
);

AOI22xp33_ASAP7_75t_L g2666 ( 
.A1(n_2582),
.A2(n_2010),
.B1(n_1988),
.B2(n_2005),
.Y(n_2666)
);

AOI221xp5_ASAP7_75t_SL g2667 ( 
.A1(n_2585),
.A2(n_2236),
.B1(n_1825),
.B2(n_2437),
.C(n_2387),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2561),
.A2(n_2005),
.B1(n_1991),
.B2(n_2134),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2571),
.B(n_2443),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2601),
.B(n_2446),
.Y(n_2670)
);

OAI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2618),
.A2(n_2099),
.B1(n_2116),
.B2(n_2082),
.Y(n_2671)
);

CKINVDCx11_ASAP7_75t_R g2672 ( 
.A(n_2584),
.Y(n_2672)
);

OA21x2_ASAP7_75t_L g2673 ( 
.A1(n_2600),
.A2(n_1812),
.B(n_1811),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2620),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_2568),
.A2(n_1991),
.B1(n_2196),
.B2(n_2179),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2606),
.B(n_2459),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2574),
.A2(n_2200),
.B1(n_2016),
.B2(n_2473),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2616),
.B(n_2459),
.Y(n_2678)
);

OAI22xp33_ASAP7_75t_L g2679 ( 
.A1(n_2618),
.A2(n_2462),
.B1(n_2337),
.B2(n_2325),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2609),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2615),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2580),
.Y(n_2682)
);

OAI22xp5_ASAP7_75t_SL g2683 ( 
.A1(n_2599),
.A2(n_2387),
.B1(n_2422),
.B2(n_2398),
.Y(n_2683)
);

AOI21xp5_ASAP7_75t_SL g2684 ( 
.A1(n_2586),
.A2(n_2398),
.B(n_2337),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2627),
.Y(n_2685)
);

AOI22xp33_ASAP7_75t_L g2686 ( 
.A1(n_2605),
.A2(n_2200),
.B1(n_2147),
.B2(n_1817),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2592),
.B(n_2462),
.Y(n_2687)
);

AOI22xp33_ASAP7_75t_L g2688 ( 
.A1(n_2625),
.A2(n_2082),
.B1(n_2116),
.B2(n_2099),
.Y(n_2688)
);

AOI222xp33_ASAP7_75t_L g2689 ( 
.A1(n_2596),
.A2(n_2385),
.B1(n_2176),
.B2(n_2486),
.C1(n_1763),
.C2(n_1777),
.Y(n_2689)
);

OAI21xp5_ASAP7_75t_SL g2690 ( 
.A1(n_2645),
.A2(n_2590),
.B(n_2607),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2674),
.B(n_2629),
.Y(n_2691)
);

OAI21xp5_ASAP7_75t_SL g2692 ( 
.A1(n_2644),
.A2(n_2590),
.B(n_2602),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2657),
.B(n_2587),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2665),
.B(n_2604),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2654),
.B(n_2631),
.Y(n_2695)
);

AO22x1_ASAP7_75t_L g2696 ( 
.A1(n_2680),
.A2(n_2598),
.B1(n_2617),
.B2(n_2622),
.Y(n_2696)
);

NAND4xp25_ASAP7_75t_L g2697 ( 
.A(n_2667),
.B(n_2614),
.C(n_2611),
.D(n_2595),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2663),
.B(n_2617),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2681),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_2649),
.B(n_2593),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_2638),
.B(n_2617),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2678),
.B(n_2480),
.Y(n_2702)
);

OAI21xp33_ASAP7_75t_SL g2703 ( 
.A1(n_2669),
.A2(n_2630),
.B(n_2471),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2640),
.B(n_2480),
.Y(n_2704)
);

OA211x2_ASAP7_75t_L g2705 ( 
.A1(n_2643),
.A2(n_2612),
.B(n_2623),
.C(n_2572),
.Y(n_2705)
);

AOI221xp5_ASAP7_75t_L g2706 ( 
.A1(n_2639),
.A2(n_2619),
.B1(n_2624),
.B2(n_2011),
.C(n_286),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2687),
.B(n_2593),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2685),
.B(n_283),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_SL g2709 ( 
.A(n_2679),
.B(n_2486),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2664),
.B(n_284),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2637),
.B(n_285),
.Y(n_2711)
);

NAND3xp33_ASAP7_75t_L g2712 ( 
.A(n_2659),
.B(n_2325),
.C(n_2303),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2676),
.B(n_286),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2670),
.B(n_2682),
.Y(n_2714)
);

AOI21x1_ASAP7_75t_L g2715 ( 
.A1(n_2673),
.A2(n_2169),
.B(n_2156),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2650),
.B(n_287),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2659),
.B(n_288),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2672),
.B(n_2612),
.Y(n_2718)
);

NAND3xp33_ASAP7_75t_L g2719 ( 
.A(n_2639),
.B(n_2342),
.C(n_2326),
.Y(n_2719)
);

AOI21xp5_ASAP7_75t_SL g2720 ( 
.A1(n_2671),
.A2(n_2169),
.B(n_2156),
.Y(n_2720)
);

OAI221xp5_ASAP7_75t_SL g2721 ( 
.A1(n_2660),
.A2(n_2565),
.B1(n_289),
.B2(n_290),
.C(n_293),
.Y(n_2721)
);

OAI21xp5_ASAP7_75t_SL g2722 ( 
.A1(n_2652),
.A2(n_288),
.B(n_289),
.Y(n_2722)
);

NAND3xp33_ASAP7_75t_L g2723 ( 
.A(n_2662),
.B(n_2372),
.C(n_2359),
.Y(n_2723)
);

OAI21xp5_ASAP7_75t_SL g2724 ( 
.A1(n_2652),
.A2(n_293),
.B(n_295),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2636),
.B(n_295),
.Y(n_2725)
);

AND2x4_ASAP7_75t_L g2726 ( 
.A(n_2691),
.B(n_2648),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2694),
.B(n_2699),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2714),
.B(n_2673),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2695),
.B(n_2684),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2707),
.B(n_2688),
.Y(n_2730)
);

AO21x2_ASAP7_75t_L g2731 ( 
.A1(n_2715),
.A2(n_2651),
.B(n_2655),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_L g2732 ( 
.A1(n_2706),
.A2(n_2647),
.B1(n_2689),
.B2(n_2666),
.Y(n_2732)
);

NOR2xp33_ASAP7_75t_L g2733 ( 
.A(n_2690),
.B(n_2700),
.Y(n_2733)
);

NAND3xp33_ASAP7_75t_L g2734 ( 
.A(n_2721),
.B(n_2653),
.C(n_2656),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2698),
.B(n_2658),
.Y(n_2735)
);

NAND3xp33_ASAP7_75t_L g2736 ( 
.A(n_2721),
.B(n_2642),
.C(n_2686),
.Y(n_2736)
);

NAND3xp33_ASAP7_75t_L g2737 ( 
.A(n_2710),
.B(n_2661),
.C(n_2641),
.Y(n_2737)
);

AO21x2_ASAP7_75t_L g2738 ( 
.A1(n_2701),
.A2(n_2661),
.B(n_2646),
.Y(n_2738)
);

INVx2_ASAP7_75t_SL g2739 ( 
.A(n_2718),
.Y(n_2739)
);

OR2x2_ASAP7_75t_L g2740 ( 
.A(n_2693),
.B(n_2683),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_SL g2741 ( 
.A(n_2703),
.B(n_2677),
.Y(n_2741)
);

NAND4xp75_ASAP7_75t_L g2742 ( 
.A(n_2705),
.B(n_2668),
.C(n_2675),
.D(n_298),
.Y(n_2742)
);

OA211x2_ASAP7_75t_L g2743 ( 
.A1(n_2701),
.A2(n_2709),
.B(n_2700),
.C(n_2717),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2704),
.B(n_296),
.Y(n_2744)
);

AO21x2_ASAP7_75t_L g2745 ( 
.A1(n_2716),
.A2(n_2708),
.B(n_2725),
.Y(n_2745)
);

NOR3xp33_ASAP7_75t_L g2746 ( 
.A(n_2722),
.B(n_297),
.C(n_298),
.Y(n_2746)
);

OR2x2_ASAP7_75t_L g2747 ( 
.A(n_2711),
.B(n_297),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2702),
.B(n_299),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2692),
.B(n_2713),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2727),
.B(n_2696),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2745),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2727),
.B(n_2697),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2739),
.B(n_2720),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2745),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2728),
.Y(n_2755)
);

NAND4xp75_ASAP7_75t_L g2756 ( 
.A(n_2743),
.B(n_2706),
.C(n_2724),
.D(n_2723),
.Y(n_2756)
);

AOI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2746),
.A2(n_2719),
.B1(n_2712),
.B2(n_2351),
.Y(n_2757)
);

XNOR2xp5_ASAP7_75t_L g2758 ( 
.A(n_2749),
.B(n_299),
.Y(n_2758)
);

NAND4xp75_ASAP7_75t_L g2759 ( 
.A(n_2741),
.B(n_300),
.C(n_301),
.D(n_302),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2726),
.B(n_302),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2729),
.B(n_2733),
.Y(n_2761)
);

XNOR2xp5_ASAP7_75t_L g2762 ( 
.A(n_2748),
.B(n_303),
.Y(n_2762)
);

OA22x2_ASAP7_75t_L g2763 ( 
.A1(n_2758),
.A2(n_2762),
.B1(n_2757),
.B2(n_2761),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2751),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2755),
.Y(n_2765)
);

XOR2xp5_ASAP7_75t_L g2766 ( 
.A(n_2756),
.B(n_2740),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2752),
.Y(n_2767)
);

XOR2xp5_ASAP7_75t_L g2768 ( 
.A(n_2759),
.B(n_2742),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2754),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2767),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2764),
.Y(n_2771)
);

AOI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2766),
.A2(n_2746),
.B1(n_2726),
.B2(n_2741),
.Y(n_2772)
);

AOI22x1_ASAP7_75t_L g2773 ( 
.A1(n_2768),
.A2(n_2753),
.B1(n_2744),
.B2(n_2747),
.Y(n_2773)
);

BUFx2_ASAP7_75t_L g2774 ( 
.A(n_2765),
.Y(n_2774)
);

OAI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2763),
.A2(n_2733),
.B1(n_2757),
.B2(n_2736),
.Y(n_2775)
);

OA22x2_ASAP7_75t_L g2776 ( 
.A1(n_2763),
.A2(n_2760),
.B1(n_2750),
.B2(n_2728),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2770),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2774),
.Y(n_2778)
);

HB1xp67_ASAP7_75t_L g2779 ( 
.A(n_2775),
.Y(n_2779)
);

BUFx2_ASAP7_75t_L g2780 ( 
.A(n_2772),
.Y(n_2780)
);

BUFx2_ASAP7_75t_L g2781 ( 
.A(n_2776),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2771),
.Y(n_2782)
);

AOI22xp5_ASAP7_75t_L g2783 ( 
.A1(n_2779),
.A2(n_2781),
.B1(n_2780),
.B2(n_2782),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_SL g2784 ( 
.A1(n_2779),
.A2(n_2773),
.B1(n_2777),
.B2(n_2731),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2778),
.Y(n_2785)
);

AOI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2779),
.A2(n_2750),
.B1(n_2731),
.B2(n_2734),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2785),
.Y(n_2787)
);

OAI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2784),
.A2(n_2769),
.B1(n_2732),
.B2(n_2737),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2783),
.Y(n_2789)
);

OAI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2786),
.A2(n_2732),
.B1(n_2730),
.B2(n_2735),
.Y(n_2790)
);

HB1xp67_ASAP7_75t_L g2791 ( 
.A(n_2785),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2791),
.Y(n_2792)
);

NOR2x1p5_ASAP7_75t_L g2793 ( 
.A(n_2789),
.B(n_2787),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2788),
.Y(n_2794)
);

AOI31xp33_ASAP7_75t_L g2795 ( 
.A1(n_2790),
.A2(n_303),
.A3(n_304),
.B(n_305),
.Y(n_2795)
);

INVx2_ASAP7_75t_SL g2796 ( 
.A(n_2791),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2791),
.Y(n_2797)
);

NOR4xp25_ASAP7_75t_L g2798 ( 
.A(n_2789),
.B(n_304),
.C(n_305),
.D(n_306),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2789),
.A2(n_2738),
.B1(n_2351),
.B2(n_309),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2796),
.Y(n_2800)
);

OR2x2_ASAP7_75t_L g2801 ( 
.A(n_2792),
.B(n_307),
.Y(n_2801)
);

AOI22xp33_ASAP7_75t_L g2802 ( 
.A1(n_2794),
.A2(n_2738),
.B1(n_308),
.B2(n_309),
.Y(n_2802)
);

NOR3xp33_ASAP7_75t_L g2803 ( 
.A(n_2795),
.B(n_307),
.C(n_310),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2793),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2797),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2799),
.Y(n_2806)
);

AOI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2799),
.A2(n_2798),
.B1(n_312),
.B2(n_313),
.Y(n_2807)
);

AO22x2_ASAP7_75t_L g2808 ( 
.A1(n_2804),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_2808)
);

OR3x2_ASAP7_75t_L g2809 ( 
.A(n_2801),
.B(n_311),
.C(n_314),
.Y(n_2809)
);

AOI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2807),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2800),
.B(n_315),
.Y(n_2811)
);

OR3x2_ASAP7_75t_L g2812 ( 
.A(n_2805),
.B(n_316),
.C(n_317),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2806),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2803),
.B(n_317),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2802),
.Y(n_2815)
);

AND2x4_ASAP7_75t_L g2816 ( 
.A(n_2811),
.B(n_318),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2808),
.Y(n_2817)
);

OAI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2812),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2809),
.Y(n_2819)
);

BUFx2_ASAP7_75t_L g2820 ( 
.A(n_2814),
.Y(n_2820)
);

AND2x4_ASAP7_75t_L g2821 ( 
.A(n_2813),
.B(n_319),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2815),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2810),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2816),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2821),
.Y(n_2825)
);

AOI22xp5_ASAP7_75t_L g2826 ( 
.A1(n_2817),
.A2(n_322),
.B1(n_323),
.B2(n_325),
.Y(n_2826)
);

AO22x2_ASAP7_75t_L g2827 ( 
.A1(n_2819),
.A2(n_325),
.B1(n_327),
.B2(n_328),
.Y(n_2827)
);

OAI22x1_ASAP7_75t_L g2828 ( 
.A1(n_2820),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_2828)
);

INVxp33_ASAP7_75t_SL g2829 ( 
.A(n_2818),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2823),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2822),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2827),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2828),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2831),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2824),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2825),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2830),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2826),
.Y(n_2838)
);

AOI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_2833),
.A2(n_2829),
.B1(n_329),
.B2(n_394),
.Y(n_2839)
);

AOI221xp5_ASAP7_75t_L g2840 ( 
.A1(n_2834),
.A2(n_392),
.B1(n_395),
.B2(n_396),
.C(n_403),
.Y(n_2840)
);

AOI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_2837),
.A2(n_408),
.B1(n_417),
.B2(n_419),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2839),
.Y(n_2842)
);

OAI22xp33_ASAP7_75t_L g2843 ( 
.A1(n_2842),
.A2(n_2832),
.B1(n_2836),
.B2(n_2838),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2843),
.Y(n_2844)
);

AOI221xp5_ASAP7_75t_L g2845 ( 
.A1(n_2844),
.A2(n_2835),
.B1(n_2840),
.B2(n_2841),
.C(n_430),
.Y(n_2845)
);

AOI211xp5_ASAP7_75t_L g2846 ( 
.A1(n_2845),
.A2(n_421),
.B(n_422),
.C(n_425),
.Y(n_2846)
);


endmodule