module fake_jpeg_3245_n_618 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_618);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_618;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g18 ( 
.A(n_17),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx12_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_68),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_33),
.Y(n_59)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_61),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_62),
.B(n_75),
.Y(n_126)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_69),
.Y(n_183)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_70),
.B(n_71),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_16),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_73),
.B(n_77),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_0),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_16),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx2_ASAP7_75t_R g83 ( 
.A(n_26),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_15),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_84),
.B(n_88),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_50),
.B(n_14),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_85),
.B(n_93),
.Y(n_129)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_14),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_92),
.B(n_97),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_24),
.B(n_14),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_25),
.B(n_13),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_105),
.Y(n_124)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_106),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_46),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_113),
.B(n_114),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_108),
.Y(n_187)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_46),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_42),
.B1(n_19),
.B2(n_35),
.Y(n_138)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_18),
.B1(n_30),
.B2(n_38),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_120),
.A2(n_122),
.B1(n_134),
.B2(n_139),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_110),
.A2(n_18),
.B1(n_30),
.B2(n_38),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_62),
.A2(n_22),
.B1(n_55),
.B2(n_34),
.Y(n_133)
);

AOI22x1_ASAP7_75t_L g249 ( 
.A1(n_133),
.A2(n_161),
.B1(n_171),
.B2(n_186),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_30),
.B1(n_38),
.B2(n_22),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_138),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_67),
.A2(n_30),
.B1(n_55),
.B2(n_22),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_75),
.A2(n_22),
.B1(n_55),
.B2(n_40),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_60),
.A2(n_41),
.B1(n_55),
.B2(n_40),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_76),
.B1(n_111),
.B2(n_78),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_61),
.A2(n_35),
.B1(n_19),
.B2(n_42),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_144),
.A2(n_188),
.B1(n_28),
.B2(n_102),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_82),
.A2(n_108),
.B1(n_65),
.B2(n_89),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_147),
.A2(n_148),
.B1(n_69),
.B2(n_57),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_66),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_34),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_153),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_81),
.B(n_34),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_41),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_156),
.B(n_157),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_41),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_79),
.B(n_25),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_158),
.B(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_98),
.B(n_40),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_160),
.B(n_166),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_104),
.A2(n_45),
.B1(n_32),
.B2(n_29),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_59),
.A2(n_30),
.B1(n_32),
.B2(n_45),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_163),
.A2(n_175),
.B1(n_179),
.B2(n_0),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_30),
.C(n_29),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_74),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_56),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_106),
.A2(n_56),
.B1(n_53),
.B2(n_36),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_83),
.A2(n_56),
.B1(n_53),
.B2(n_36),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_109),
.B(n_53),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_72),
.A2(n_36),
.B1(n_20),
.B2(n_54),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_80),
.A2(n_20),
.B(n_51),
.C(n_54),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_180),
.A2(n_165),
.B(n_130),
.C(n_173),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_94),
.A2(n_20),
.B1(n_51),
.B2(n_54),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_64),
.A2(n_28),
.B1(n_10),
.B2(n_9),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_137),
.A2(n_95),
.B1(n_113),
.B2(n_87),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_189),
.Y(n_271)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_190),
.Y(n_289)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_191),
.Y(n_285)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_193),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_149),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_195),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_151),
.A2(n_28),
.B1(n_63),
.B2(n_86),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_196),
.A2(n_221),
.B1(n_226),
.B2(n_227),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_197),
.B(n_215),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_198),
.Y(n_287)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_199),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_69),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_200),
.B(n_202),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

INVx4_ASAP7_75t_SL g272 ( 
.A(n_201),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_203),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_204),
.B(n_209),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_205),
.A2(n_234),
.B1(n_237),
.B2(n_251),
.Y(n_259)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_125),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_208),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_57),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_182),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_214),
.Y(n_263)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_212),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_146),
.B(n_9),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_216),
.A2(n_219),
.B(n_241),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_217),
.Y(n_312)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_218),
.Y(n_273)
);

NAND2x1_ASAP7_75t_SL g219 ( 
.A(n_125),
.B(n_0),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_220),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_125),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_1),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_223),
.C(n_256),
.Y(n_261)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_126),
.B(n_1),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_178),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_225),
.B(n_228),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_177),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_127),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_227)
);

NAND2xp33_ASAP7_75t_R g228 ( 
.A(n_129),
.B(n_2),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_230),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_124),
.B(n_5),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_233),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_159),
.B(n_5),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_232),
.B(n_235),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_149),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_147),
.A2(n_7),
.B1(n_8),
.B2(n_160),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_124),
.B(n_8),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_132),
.B(n_8),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_238),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_156),
.A2(n_8),
.B1(n_157),
.B2(n_150),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_162),
.B(n_181),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_239),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_162),
.B(n_123),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_246),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_168),
.A2(n_187),
.B1(n_150),
.B2(n_141),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_253),
.B1(n_155),
.B2(n_119),
.Y(n_276)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_136),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_244),
.Y(n_309)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_167),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_247),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_123),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_255),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_141),
.A2(n_187),
.B1(n_168),
.B2(n_184),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_169),
.A2(n_174),
.B1(n_184),
.B2(n_176),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_176),
.B1(n_174),
.B2(n_169),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_130),
.A2(n_173),
.B1(n_164),
.B2(n_154),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_254),
.Y(n_296)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_152),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_130),
.B(n_185),
.C(n_170),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_152),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_155),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_250),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_258),
.B(n_283),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_260),
.A2(n_280),
.B1(n_286),
.B2(n_308),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_229),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_264),
.B(n_281),
.C(n_295),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_194),
.A2(n_234),
.B1(n_241),
.B2(n_202),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_265),
.A2(n_304),
.B1(n_318),
.B2(n_191),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_276),
.A2(n_207),
.B1(n_201),
.B2(n_230),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_197),
.A2(n_121),
.B(n_154),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_279),
.A2(n_291),
.B(n_248),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_212),
.A2(n_185),
.B1(n_170),
.B2(n_164),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_121),
.C(n_167),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_117),
.Y(n_283)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_194),
.A2(n_119),
.B1(n_135),
.B2(n_249),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_232),
.B(n_135),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_290),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_217),
.A2(n_213),
.B(n_211),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_223),
.B(n_256),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_204),
.B(n_223),
.C(n_189),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_247),
.C(n_279),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_192),
.B(n_235),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_299),
.B(n_306),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_254),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_201),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_205),
.A2(n_237),
.B1(n_249),
.B2(n_227),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_192),
.B(n_203),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_222),
.A2(n_249),
.B1(n_189),
.B2(n_216),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_222),
.B(n_219),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_319),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_190),
.B(n_210),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_315),
.B(n_288),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_189),
.A2(n_216),
.B1(n_225),
.B2(n_199),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_224),
.B1(n_195),
.B2(n_193),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_243),
.A2(n_251),
.B1(n_252),
.B2(n_216),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_219),
.B(n_216),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_287),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_321),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_322),
.A2(n_332),
.B(n_333),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_287),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_324),
.B(n_328),
.Y(n_398)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_275),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g385 ( 
.A(n_325),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_246),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_326),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_282),
.Y(n_328)
);

OAI22x1_ASAP7_75t_L g329 ( 
.A1(n_270),
.A2(n_247),
.B1(n_242),
.B2(n_230),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_360),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_271),
.A2(n_233),
.B(n_239),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_268),
.A2(n_244),
.B(n_218),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_344),
.Y(n_379)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_338),
.A2(n_358),
.B1(n_285),
.B2(n_294),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_258),
.B(n_257),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_341),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_271),
.A2(n_195),
.B(n_255),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_340),
.A2(n_353),
.B(n_305),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_264),
.B(n_245),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_314),
.A2(n_201),
.B1(n_230),
.B2(n_242),
.Y(n_344)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_295),
.B(n_242),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_347),
.C(n_351),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_265),
.B(n_247),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_348),
.B(n_350),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_283),
.B(n_302),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_261),
.B(n_302),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_268),
.A2(n_291),
.B(n_319),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_314),
.A2(n_308),
.B1(n_317),
.B2(n_286),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_363),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_267),
.B(n_261),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_355),
.B(n_357),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_304),
.A2(n_259),
.B1(n_270),
.B2(n_269),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_356),
.A2(n_361),
.B1(n_367),
.B2(n_273),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_277),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_259),
.A2(n_318),
.B1(n_297),
.B2(n_267),
.Y(n_358)
);

AOI32xp33_ASAP7_75t_L g359 ( 
.A1(n_263),
.A2(n_274),
.A3(n_310),
.B1(n_266),
.B2(n_313),
.Y(n_359)
);

AOI21xp33_ASAP7_75t_L g414 ( 
.A1(n_359),
.A2(n_365),
.B(n_374),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_269),
.A2(n_281),
.B1(n_276),
.B2(n_313),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_293),
.B(n_312),
.C(n_280),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_311),
.C(n_320),
.Y(n_397)
);

INVx3_ASAP7_75t_SL g363 ( 
.A(n_272),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_275),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_364),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_288),
.B(n_312),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_292),
.Y(n_366)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_260),
.A2(n_307),
.B1(n_298),
.B2(n_301),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_272),
.A2(n_262),
.B1(n_309),
.B2(n_303),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_368),
.A2(n_369),
.B1(n_373),
.B2(n_370),
.Y(n_410)
);

AOI22x1_ASAP7_75t_SL g369 ( 
.A1(n_307),
.A2(n_298),
.B1(n_301),
.B2(n_292),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_275),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_370),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_309),
.B(n_316),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_278),
.Y(n_405)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_296),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_372),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_272),
.A2(n_262),
.B1(n_309),
.B2(n_303),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g374 ( 
.A(n_307),
.B(n_316),
.CI(n_300),
.CON(n_374),
.SN(n_374)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_375),
.A2(n_377),
.B1(n_408),
.B2(n_416),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_327),
.A2(n_296),
.B1(n_273),
.B2(n_285),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_294),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_378),
.B(n_389),
.C(n_397),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_380),
.A2(n_420),
.B1(n_326),
.B2(n_341),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_371),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_405),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_388),
.A2(n_392),
.B(n_419),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_311),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_353),
.A2(n_320),
.B(n_305),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_343),
.Y(n_395)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_366),
.Y(n_400)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_400),
.Y(n_434)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_402),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_351),
.B(n_346),
.C(n_355),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_411),
.C(n_362),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_338),
.A2(n_278),
.B1(n_305),
.B2(n_358),
.Y(n_408)
);

OAI21xp33_ASAP7_75t_SL g455 ( 
.A1(n_410),
.A2(n_325),
.B(n_344),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_330),
.B(n_347),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_412),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_356),
.A2(n_323),
.B1(n_361),
.B2(n_348),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_417),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_322),
.A2(n_332),
.B(n_333),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_418),
.A2(n_369),
.B(n_359),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_331),
.A2(n_326),
.B(n_340),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_354),
.A2(n_323),
.B1(n_350),
.B2(n_330),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_418),
.A2(n_331),
.B(n_329),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_421),
.B(n_433),
.Y(n_480)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_385),
.Y(n_423)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_423),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_398),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_438),
.Y(n_470)
);

AO21x1_ASAP7_75t_L g469 ( 
.A1(n_425),
.A2(n_436),
.B(n_419),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_426),
.A2(n_392),
.B(n_379),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_378),
.B(n_336),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_427),
.B(n_440),
.C(n_393),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_420),
.A2(n_334),
.B1(n_367),
.B2(n_357),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_429),
.A2(n_390),
.B1(n_417),
.B2(n_407),
.Y(n_466)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_430),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_416),
.A2(n_408),
.B1(n_375),
.B2(n_409),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_431),
.A2(n_456),
.B1(n_459),
.B2(n_443),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_388),
.Y(n_433)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_404),
.Y(n_435)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_401),
.A2(n_328),
.B1(n_365),
.B2(n_336),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_389),
.B(n_360),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_406),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_409),
.B(n_349),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_349),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_439),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_399),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_441),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_399),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_443),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_413),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_447),
.Y(n_481)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_386),
.Y(n_448)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_386),
.Y(n_449)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_449),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_384),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_451),
.B(n_458),
.Y(n_488)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_391),
.Y(n_452)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_391),
.Y(n_453)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_453),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_382),
.B(n_364),
.Y(n_454)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_455),
.A2(n_381),
.B1(n_379),
.B2(n_376),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_412),
.A2(n_374),
.B1(n_324),
.B2(n_321),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_390),
.B(n_363),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_401),
.A2(n_363),
.B1(n_374),
.B2(n_387),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_394),
.Y(n_460)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_413),
.B(n_387),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_464),
.A2(n_444),
.B(n_421),
.Y(n_498)
);

XOR2x2_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_411),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_465),
.B(n_478),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_466),
.A2(n_473),
.B1(n_493),
.B2(n_494),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_467),
.B(n_450),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_469),
.B(n_475),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_SL g471 ( 
.A(n_459),
.B(n_401),
.C(n_393),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_471),
.B(n_446),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_472),
.B(n_482),
.C(n_489),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_425),
.A2(n_380),
.B1(n_379),
.B2(n_407),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_454),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_428),
.B(n_414),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_428),
.B(n_397),
.C(n_383),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_484),
.A2(n_491),
.B1(n_445),
.B2(n_421),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_436),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_486),
.B(n_469),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_487),
.B(n_404),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_440),
.B(n_383),
.C(n_405),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_429),
.A2(n_381),
.B1(n_403),
.B2(n_394),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_441),
.A2(n_426),
.B1(n_445),
.B2(n_433),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_437),
.B(n_395),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_467),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_488),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_497),
.B(n_501),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_498),
.A2(n_524),
.B(n_476),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_461),
.B(n_479),
.Y(n_499)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_499),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_461),
.B(n_446),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_502),
.B(n_503),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_470),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_485),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_504),
.B(n_505),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_490),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_495),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_507),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_508),
.A2(n_511),
.B1(n_493),
.B2(n_494),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_466),
.A2(n_431),
.B1(n_457),
.B2(n_444),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_509),
.A2(n_516),
.B1(n_519),
.B2(n_520),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_510),
.B(n_474),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_472),
.B(n_450),
.C(n_456),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_513),
.B(n_521),
.C(n_523),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_491),
.A2(n_432),
.B1(n_453),
.B2(n_452),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_514),
.A2(n_477),
.B1(n_400),
.B2(n_402),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_464),
.Y(n_528)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_485),
.Y(n_516)
);

XNOR2x1_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_484),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_462),
.B(n_482),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_518),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_473),
.A2(n_432),
.B1(n_449),
.B2(n_448),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_479),
.A2(n_460),
.B1(n_434),
.B2(n_422),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_465),
.B(n_442),
.C(n_422),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_489),
.B(n_396),
.Y(n_522)
);

NOR4xp25_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_480),
.C(n_492),
.D(n_468),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_478),
.B(n_471),
.C(n_481),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_487),
.B(n_442),
.Y(n_524)
);

AO21x1_ASAP7_75t_L g559 ( 
.A1(n_525),
.A2(n_536),
.B(n_519),
.Y(n_559)
);

A2O1A1O1Ixp25_ASAP7_75t_L g526 ( 
.A1(n_500),
.A2(n_498),
.B(n_480),
.C(n_523),
.D(n_513),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_526),
.B(n_532),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_527),
.B(n_504),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_528),
.B(n_540),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_529),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_509),
.A2(n_481),
.B1(n_492),
.B2(n_483),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_463),
.C(n_490),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_534),
.B(n_541),
.C(n_515),
.Y(n_554)
);

XNOR2x1_ASAP7_75t_L g540 ( 
.A(n_517),
.B(n_463),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_483),
.C(n_468),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_503),
.A2(n_477),
.B1(n_476),
.B2(n_434),
.Y(n_543)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_543),
.Y(n_550)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_544),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_505),
.B(n_435),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_502),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_546),
.B(n_547),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_496),
.A2(n_474),
.B1(n_423),
.B2(n_430),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_499),
.Y(n_548)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_548),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_530),
.B(n_521),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_549),
.B(n_554),
.Y(n_585)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_551),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_552),
.B(n_568),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_536),
.A2(n_496),
.B(n_511),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_553),
.A2(n_539),
.B(n_529),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_534),
.B(n_510),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_557),
.B(n_531),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_559),
.A2(n_526),
.B(n_544),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_528),
.B(n_506),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_560),
.B(n_563),
.Y(n_578)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_537),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_562),
.B(n_548),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_533),
.B(n_506),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_546),
.B(n_524),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_565),
.B(n_567),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_531),
.B(n_524),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_541),
.B(n_524),
.C(n_514),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_556),
.A2(n_535),
.B1(n_542),
.B2(n_538),
.Y(n_569)
);

INVxp33_ASAP7_75t_L g597 ( 
.A(n_569),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_570),
.B(n_572),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_554),
.B(n_537),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_567),
.B(n_516),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_573),
.B(n_574),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_568),
.B(n_532),
.C(n_545),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_576),
.C(n_561),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_563),
.B(n_545),
.C(n_540),
.Y(n_576)
);

OAI21xp33_ASAP7_75t_L g595 ( 
.A1(n_577),
.A2(n_579),
.B(n_565),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_551),
.B(n_539),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_559),
.B(n_525),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_582),
.B(n_584),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_583),
.A2(n_566),
.B(n_558),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_553),
.A2(n_520),
.B1(n_547),
.B2(n_385),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_585),
.B(n_575),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_587),
.B(n_588),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_571),
.B(n_550),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_590),
.B(n_595),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_583),
.A2(n_566),
.B(n_551),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_591),
.A2(n_555),
.B(n_581),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_569),
.B(n_564),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_592),
.B(n_593),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_564),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_594),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_580),
.B(n_385),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_576),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_597),
.A2(n_577),
.B1(n_579),
.B2(n_584),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_599),
.B(n_600),
.Y(n_609)
);

NOR3x1_ASAP7_75t_SL g602 ( 
.A(n_597),
.B(n_555),
.C(n_581),
.Y(n_602)
);

AO21x1_ASAP7_75t_L g607 ( 
.A1(n_602),
.A2(n_604),
.B(n_591),
.Y(n_607)
);

MAJx2_ASAP7_75t_L g611 ( 
.A(n_607),
.B(n_605),
.C(n_590),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_603),
.B(n_594),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_608),
.B(n_610),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_606),
.B(n_589),
.C(n_598),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_611),
.B(n_613),
.C(n_586),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_609),
.A2(n_601),
.B(n_605),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_614),
.B(n_615),
.C(n_578),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_612),
.B(n_578),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_595),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_617),
.B(n_560),
.Y(n_618)
);


endmodule