module real_jpeg_33495_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_1),
.B(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_1),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_1),
.B(n_282),
.Y(n_281)
);

NAND2x1_ASAP7_75t_L g377 ( 
.A(n_1),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_1),
.B(n_428),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_2),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_2),
.B(n_32),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_2),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_2),
.B(n_413),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_3),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_4),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_4),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_4),
.B(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_4),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_4),
.B(n_391),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_4),
.Y(n_419)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_5),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_5),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_5),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_5),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_5),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_5),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_5),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_5),
.B(n_396),
.Y(n_395)
);

NAND2xp33_ASAP7_75t_R g48 ( 
.A(n_6),
.B(n_49),
.Y(n_48)
);

AO22x1_ASAP7_75t_L g59 ( 
.A1(n_6),
.A2(n_11),
.B1(n_49),
.B2(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_6),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_6),
.B(n_125),
.Y(n_124)
);

NAND2x1_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_6),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_6),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_6),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_6),
.B(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_7),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_8),
.Y(n_86)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_9),
.Y(n_177)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_10),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_11),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_11),
.B(n_148),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_11),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_11),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_11),
.B(n_415),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_12),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_12),
.B(n_365),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_12),
.B(n_434),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_14),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_14),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_14),
.B(n_83),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_14),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_14),
.Y(n_224)
);

NAND2x1_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_15),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_15),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_15),
.B(n_32),
.Y(n_150)
);

AND2x4_ASAP7_75t_SL g261 ( 
.A(n_15),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_15),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_15),
.B(n_43),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_15),
.B(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_17),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_17),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_17),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_18),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_18),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_18),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_18),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_18),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_18),
.B(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_19),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_401),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_347),
.B(n_399),
.Y(n_23)
);

AOI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_248),
.B(n_344),
.Y(n_24)
);

AO21x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_151),
.B(n_247),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_132),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_27),
.B(n_132),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_79),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_28),
.B(n_342),
.C(n_343),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_46),
.Y(n_28)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_29),
.B(n_47),
.C(n_64),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_37),
.C(n_41),
.Y(n_29)
);

XNOR2x2_ASAP7_75t_L g136 ( 
.A(n_30),
.B(n_137),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_31),
.B(n_33),
.Y(n_139)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_36),
.Y(n_211)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_37),
.B(n_42),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_40),
.Y(n_276)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_45),
.Y(n_260)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_64),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_54),
.B(n_59),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_52),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_53),
.Y(n_319)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_58),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_59),
.B(n_303),
.C(n_309),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_59),
.A2(n_309),
.B1(n_310),
.B2(n_335),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_59),
.Y(n_335)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_63),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_63),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_65),
.B(n_73),
.C(n_78),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_67),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_78),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_71),
.Y(n_413)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_76),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_116),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_80),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_96),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_81),
.B(n_97),
.C(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_82),
.B(n_90),
.C(n_94),
.Y(n_310)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_86),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_86),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_86),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_86),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_105),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_105),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_112),
.Y(n_105)
);

XNOR2x1_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_116),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_131),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_131),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.C(n_127),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_120),
.A2(n_121),
.B1(n_127),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_126),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_126),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_127),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.C(n_138),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_134),
.B(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_136),
.B(n_138),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.C(n_145),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_144),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_145),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_150),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_241),
.B(n_246),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_191),
.B(n_240),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_183),
.Y(n_153)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_154),
.B(n_183),
.Y(n_240)
);

OAI21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_169),
.B(n_182),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_156),
.B(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_166),
.C(n_168),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_173),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_177),
.Y(n_365)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx4f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_185),
.B(n_189),
.C(n_243),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_204),
.B(n_239),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_202),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_202),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.C(n_200),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_195),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_195),
.B(n_219),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_200),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_221),
.B(n_236),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_218),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_208),
.B1(n_212),
.B2(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_207),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_229),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_228),
.Y(n_271)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_228),
.Y(n_435)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_244),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_329),
.B(n_337),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_249),
.B(n_329),
.C(n_345),
.Y(n_344)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_278),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_250),
.B(n_279),
.C(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_266),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2x2_ASAP7_75t_L g330 ( 
.A(n_252),
.B(n_331),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_255),
.A2(n_266),
.B1(n_267),
.B2(n_332),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_255),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_259),
.C(n_264),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_258)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_261),
.Y(n_264)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2x2_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_277),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_301),
.Y(n_278)
);

XOR2x2_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_289),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_280),
.B(n_290),
.C(n_291),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_281),
.B(n_284),
.C(n_287),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_281),
.B(n_284),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_281),
.B(n_284),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g446 ( 
.A1(n_287),
.A2(n_389),
.B(n_395),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_292),
.B(n_297),
.C(n_299),
.Y(n_367)
);

BUFx12f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_L g362 ( 
.A(n_299),
.B(n_363),
.Y(n_362)
);

MAJx2_ASAP7_75t_L g444 ( 
.A(n_299),
.B(n_361),
.C(n_364),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_311),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

XOR2x2_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_313)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_320),
.B1(n_321),
.B2(n_328),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_312),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_315),
.C(n_385),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_317),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_317),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_324),
.B(n_326),
.C(n_327),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_325),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.C(n_336),
.Y(n_329)
);

AOI221xp5_ASAP7_75t_L g337 ( 
.A1(n_330),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.C(n_341),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_338),
.Y(n_346)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_336),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

NOR2x1_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_352),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_358),
.C(n_404),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.C(n_356),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_380),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_366),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_359),
.B(n_367),
.C(n_368),
.Y(n_437)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_363),
.B(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_377),
.C(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_377),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_373),
.Y(n_424)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_380),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_383),
.B2(n_398),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_384),
.C(n_386),
.Y(n_406)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_383),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_389),
.A2(n_390),
.B1(n_394),
.B2(n_395),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_389),
.A2(n_390),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_389),
.B(n_395),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_389),
.B(n_395),
.Y(n_451)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_454),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_405),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_403),
.B(n_405),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_436),
.B1(n_452),
.B2(n_453),
.Y(n_407)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_425),
.Y(n_408)
);

XNOR2x1_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_423),
.Y(n_409)
);

XNOR2x2_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_418),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_431),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_436),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_445),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_444),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_442),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_447),
.B(n_448),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B(n_451),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);


endmodule