module fake_netlist_5_1325_n_1118 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1118);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1118;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_194;
wire n_316;
wire n_785;
wire n_855;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_697;
wire n_376;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_1055;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_864;
wire n_443;
wire n_173;
wire n_859;
wire n_1110;
wire n_951;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_314;
wire n_247;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_516;
wire n_498;
wire n_933;
wire n_385;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_186;
wire n_537;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_171;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_519;
wire n_406;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_167;
wire n_976;
wire n_1096;
wire n_1095;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_1114;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_163;
wire n_339;
wire n_882;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_962;
wire n_181;
wire n_436;
wire n_930;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_922;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_974;
wire n_432;
wire n_164;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_928;
wire n_1064;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_517;
wire n_342;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_736;
wire n_893;
wire n_502;
wire n_892;
wire n_595;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_699;
wire n_632;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_846;
wire n_586;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_170;
wire n_332;
wire n_1053;
wire n_1101;
wire n_161;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_176;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_795;
wire n_695;
wire n_832;
wire n_180;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_205;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_1037;
wire n_202;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_965;
wire n_364;
wire n_319;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_200;
wire n_1056;
wire n_162;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_187;
wire n_348;
wire n_1029;
wire n_166;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_104),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_93),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_20),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_13),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_68),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_59),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_24),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_64),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_13),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_31),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_160),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_9),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_31),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_66),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_98),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_127),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_115),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_0),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_100),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_41),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_25),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_149),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_44),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_81),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_88),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_154),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_28),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_112),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_39),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_67),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_119),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_78),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_123),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_56),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_53),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_110),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_139),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_152),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_14),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_39),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_54),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_84),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_179),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_167),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_182),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_162),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_178),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_197),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_202),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_199),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_169),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_171),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_239),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_212),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_213),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_215),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_216),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_204),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_217),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_173),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_229),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_222),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_230),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_219),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_238),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_238),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_212),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_225),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_242),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_242),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_262),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_256),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_243),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_287),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_278),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_278),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_244),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_251),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_266),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_281),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_281),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_287),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_260),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_282),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_282),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_284),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_277),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_245),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_288),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_289),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_293),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_294),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_293),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_294),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_297),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_295),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_297),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_304),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_312),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_295),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_312),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_305),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_284),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_316),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_316),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_299),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_324),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_322),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_326),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_317),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_317),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_325),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_325),
.B(n_245),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_271),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_328),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_329),
.B(n_246),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_366),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_246),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_337),
.A2(n_276),
.B1(n_275),
.B2(n_247),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_247),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_350),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_341),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_367),
.Y(n_383)
);

BUFx12f_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_344),
.A2(n_320),
.B1(n_272),
.B2(n_268),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_270),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_330),
.B(n_327),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_362),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_332),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_332),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_334),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_339),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_338),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_345),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_348),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

OA21x2_ASAP7_75t_L g408 ( 
.A1(n_353),
.A2(n_318),
.B(n_306),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_320),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_357),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_357),
.B(n_320),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_343),
.B(n_270),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_263),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_346),
.B(n_273),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_368),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_360),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

NOR2x1_ASAP7_75t_L g427 ( 
.A(n_369),
.B(n_273),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_342),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_363),
.B(n_273),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_360),
.A2(n_324),
.B1(n_311),
.B2(n_310),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_350),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_347),
.Y(n_434)
);

BUFx8_ASAP7_75t_L g435 ( 
.A(n_350),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_347),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_347),
.B(n_283),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_330),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_329),
.B(n_263),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_360),
.A2(n_311),
.B1(n_310),
.B2(n_163),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_333),
.A2(n_272),
.B1(n_267),
.B2(n_268),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_333),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_L g444 ( 
.A(n_342),
.B(n_273),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_363),
.B(n_273),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_426),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_402),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_423),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_424),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_372),
.B(n_374),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_411),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_426),
.Y(n_455)
);

CKINVDCx8_ASAP7_75t_R g456 ( 
.A(n_411),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_439),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_425),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_439),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_384),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_402),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_384),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_397),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_429),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_429),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_372),
.B(n_255),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_397),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_397),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_372),
.B(n_327),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_373),
.B(n_258),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_432),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_379),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_441),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_435),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_267),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_435),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_397),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_383),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_379),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_446),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_454),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_454),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_457),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_R g487 ( 
.A(n_457),
.B(n_414),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_478),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_476),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_447),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_478),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

BUFx8_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_450),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_447),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_466),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_459),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_456),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_456),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_449),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_476),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_461),
.Y(n_505)
);

BUFx6f_ASAP7_75t_SL g506 ( 
.A(n_470),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_471),
.B(n_440),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_460),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_463),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_463),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_453),
.B(n_379),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_447),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_475),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_450),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_477),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_470),
.B(n_378),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_464),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_467),
.B(n_375),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_507),
.A2(n_453),
.B1(n_195),
.B2(n_175),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_518),
.B(n_380),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_491),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_517),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_496),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_491),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_495),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_492),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_511),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_483),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_499),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_492),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_487),
.A2(n_392),
.B1(n_438),
.B2(n_419),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_501),
.B(n_464),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_504),
.B(n_455),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_497),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_490),
.B(n_380),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_489),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_R g538 ( 
.A(n_516),
.B(n_468),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_502),
.B(n_468),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_494),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_506),
.A2(n_453),
.B1(n_474),
.B2(n_191),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_486),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_514),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_514),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_483),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_511),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_483),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_511),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_506),
.Y(n_550)
);

NOR2x1p5_ASAP7_75t_L g551 ( 
.A(n_486),
.B(n_396),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_506),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_503),
.A2(n_438),
.B1(n_419),
.B2(n_442),
.Y(n_553)
);

BUFx4f_ASAP7_75t_L g554 ( 
.A(n_484),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_496),
.Y(n_555)
);

OAI22xp33_ASAP7_75t_L g556 ( 
.A1(n_493),
.A2(n_469),
.B1(n_479),
.B2(n_433),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_505),
.B(n_434),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_496),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_485),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_500),
.B(n_433),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_493),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_512),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_498),
.B(n_433),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_498),
.A2(n_191),
.B1(n_388),
.B2(n_374),
.Y(n_564)
);

BUFx4f_ASAP7_75t_L g565 ( 
.A(n_508),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_509),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_510),
.B(n_403),
.Y(n_567)
);

BUFx8_ASAP7_75t_SL g568 ( 
.A(n_515),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_513),
.Y(n_569)
);

BUFx10_ASAP7_75t_L g570 ( 
.A(n_486),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_511),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_507),
.B(n_403),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_517),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_489),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_504),
.B(n_422),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_507),
.B(n_433),
.Y(n_576)
);

AND2x2_ASAP7_75t_SL g577 ( 
.A(n_507),
.B(n_444),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_488),
.Y(n_578)
);

A2O1A1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_507),
.A2(n_383),
.B(n_390),
.C(n_387),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_491),
.Y(n_580)
);

INVx6_ASAP7_75t_L g581 ( 
.A(n_496),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_496),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_507),
.B(n_433),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_483),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_491),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_507),
.B(n_409),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_511),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_507),
.B(n_377),
.C(n_395),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_488),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_488),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_483),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_507),
.B(n_403),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_491),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_511),
.B(n_446),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_507),
.B(n_412),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_507),
.B(n_386),
.Y(n_597)
);

BUFx4f_ASAP7_75t_L g598 ( 
.A(n_516),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_550),
.B(n_469),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_554),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_574),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_598),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_522),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_598),
.B(n_572),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_554),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_576),
.B(n_451),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_576),
.B(n_451),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_537),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_541),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_552),
.B(n_555),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_593),
.B(n_547),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_560),
.B(n_446),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_479),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_565),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_575),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_528),
.B(n_419),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_577),
.B(n_394),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_597),
.B(n_589),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_525),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g620 ( 
.A(n_538),
.B(n_397),
.Y(n_620)
);

AND2x6_ASAP7_75t_L g621 ( 
.A(n_558),
.B(n_446),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_521),
.B(n_569),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_584),
.B(n_452),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_519),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_565),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_520),
.A2(n_191),
.B1(n_207),
.B2(n_164),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

INVx6_ASAP7_75t_L g628 ( 
.A(n_543),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_526),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_531),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_530),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_535),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_578),
.Y(n_633)
);

BUFx4f_ASAP7_75t_L g634 ( 
.A(n_581),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_580),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_520),
.B(n_399),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_584),
.B(n_452),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_577),
.B(n_421),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_587),
.B(n_458),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_543),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_555),
.B(n_446),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_534),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_587),
.B(n_421),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_558),
.B(n_473),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_590),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_591),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_568),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_529),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_544),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_560),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_549),
.B(n_571),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_596),
.B(n_430),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_570),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_571),
.B(n_588),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_561),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_596),
.B(n_458),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_567),
.B(n_418),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_579),
.B(n_462),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_579),
.B(n_394),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_545),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_581),
.B(n_473),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_539),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_539),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_586),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_592),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_592),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_556),
.B(n_404),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_588),
.B(n_422),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_532),
.B(n_399),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_542),
.B(n_399),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_581),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_529),
.Y(n_672)
);

AND2x6_ASAP7_75t_L g673 ( 
.A(n_524),
.B(n_473),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_594),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_594),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_SL g676 ( 
.A(n_556),
.B(n_404),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_624),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_608),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_629),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_618),
.B(n_563),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_608),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_618),
.B(n_542),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_615),
.B(n_534),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_615),
.B(n_536),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_600),
.B(n_523),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_657),
.B(n_559),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_601),
.Y(n_687)
);

BUFx6f_ASAP7_75t_SL g688 ( 
.A(n_625),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_631),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_620),
.B(n_553),
.Y(n_690)
);

NOR2xp67_ASAP7_75t_SL g691 ( 
.A(n_671),
.B(n_399),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_667),
.B(n_564),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_626),
.A2(n_564),
.B1(n_395),
.B2(n_406),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_647),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_628),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_609),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_611),
.B(n_622),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_634),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_633),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_645),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_646),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_604),
.B(n_557),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_649),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_652),
.B(n_546),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_613),
.B(n_548),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_663),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_L g707 ( 
.A(n_605),
.B(n_523),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_667),
.B(n_427),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_606),
.B(n_551),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_660),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_676),
.B(n_398),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_662),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_634),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_606),
.B(n_418),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_628),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_636),
.A2(n_420),
.B(n_418),
.C(n_524),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_664),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_613),
.B(n_533),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_607),
.B(n_623),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_675),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_607),
.B(n_420),
.Y(n_721)
);

NOR2x1_ASAP7_75t_L g722 ( 
.A(n_640),
.B(n_573),
.Y(n_722)
);

NOR2x1p5_ASAP7_75t_L g723 ( 
.A(n_653),
.B(n_582),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_SL g724 ( 
.A(n_602),
.B(n_538),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_628),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_623),
.B(n_420),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_637),
.B(n_413),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_SL g728 ( 
.A(n_671),
.B(n_399),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_617),
.B(n_540),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_643),
.B(n_413),
.Y(n_730)
);

BUFx4_ASAP7_75t_L g731 ( 
.A(n_655),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_610),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_643),
.B(n_573),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_626),
.B(n_407),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_603),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_670),
.A2(n_208),
.B1(n_207),
.B2(n_205),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_610),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_674),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_659),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_602),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_650),
.B(n_582),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_602),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_638),
.B(n_583),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_638),
.B(n_583),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_698),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_719),
.B(n_639),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_682),
.A2(n_669),
.B1(n_671),
.B2(n_472),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_682),
.A2(n_676),
.B1(n_659),
.B2(n_668),
.Y(n_748)
);

BUFx8_ASAP7_75t_L g749 ( 
.A(n_688),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_700),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_697),
.B(n_639),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_677),
.Y(n_752)
);

AO22x2_ASAP7_75t_L g753 ( 
.A1(n_678),
.A2(n_599),
.B1(n_651),
.B2(n_641),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_692),
.A2(n_671),
.B1(n_599),
.B2(n_612),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_700),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_679),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_696),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_703),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_731),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_732),
.B(n_672),
.Y(n_760)
);

BUFx8_ASAP7_75t_L g761 ( 
.A(n_688),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_743),
.B(n_642),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_732),
.B(n_651),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_734),
.B(n_656),
.C(n_406),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_710),
.Y(n_765)
);

AO22x2_ASAP7_75t_L g766 ( 
.A1(n_681),
.A2(n_641),
.B1(n_648),
.B2(n_658),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_684),
.B(n_642),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_689),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_744),
.B(n_614),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_699),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_737),
.B(n_648),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_701),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_687),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_712),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_718),
.B(n_654),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_714),
.B(n_619),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_692),
.A2(n_562),
.B1(n_616),
.B2(n_371),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_721),
.B(n_627),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_736),
.A2(n_612),
.B1(n_417),
.B2(n_405),
.Y(n_779)
);

AOI211xp5_ASAP7_75t_L g780 ( 
.A1(n_690),
.A2(n_208),
.B(n_183),
.C(n_188),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_738),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_733),
.B(n_566),
.Y(n_782)
);

AO22x2_ASAP7_75t_L g783 ( 
.A1(n_739),
.A2(n_658),
.B1(n_654),
.B2(n_632),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_726),
.B(n_630),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_724),
.A2(n_371),
.B1(n_673),
.B2(n_661),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_680),
.A2(n_371),
.B1(n_185),
.B2(n_190),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_706),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_737),
.B(n_661),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_680),
.A2(n_371),
.B1(n_190),
.B2(n_205),
.Y(n_789)
);

NAND2x1p5_ASAP7_75t_L g790 ( 
.A(n_691),
.B(n_665),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_715),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_717),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_720),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_735),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_704),
.B(n_635),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_741),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_695),
.B(n_661),
.Y(n_797)
);

NOR4xp25_ASAP7_75t_SL g798 ( 
.A(n_708),
.B(n_417),
.C(n_405),
.D(n_673),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_683),
.B(n_673),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_709),
.Y(n_800)
);

AO22x2_ASAP7_75t_L g801 ( 
.A1(n_711),
.A2(n_400),
.B1(n_410),
.B2(n_398),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_SL g802 ( 
.A1(n_718),
.A2(n_415),
.B1(n_407),
.B2(n_404),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_705),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_729),
.A2(n_371),
.B1(n_673),
.B2(n_644),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_705),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_698),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_729),
.A2(n_205),
.B1(n_167),
.B2(n_210),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_686),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_727),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_702),
.B(n_570),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_730),
.B(n_673),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_725),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_722),
.Y(n_813)
);

AND2x2_ASAP7_75t_SL g814 ( 
.A(n_748),
.B(n_698),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_L g815 ( 
.A1(n_780),
.A2(n_716),
.B(n_711),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_764),
.A2(n_708),
.B(n_444),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_747),
.A2(n_693),
.B1(n_713),
.B2(n_698),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_745),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_803),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_800),
.B(n_723),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_759),
.B(n_713),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_805),
.B(n_685),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_809),
.A2(n_713),
.B1(n_742),
.B2(n_740),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_751),
.B(n_707),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_749),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_745),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_762),
.B(n_694),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_813),
.B(n_740),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_807),
.A2(n_728),
.B(n_200),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_771),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_754),
.B(n_742),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_808),
.B(n_742),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_749),
.B(n_407),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_796),
.B(n_665),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_777),
.A2(n_210),
.B1(n_167),
.B2(n_201),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_761),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_745),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_757),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_806),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_761),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_767),
.B(n_568),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_750),
.Y(n_842)
);

NOR2x2_ASAP7_75t_L g843 ( 
.A(n_773),
.B(n_400),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_755),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_746),
.B(n_621),
.Y(n_845)
);

NOR3xp33_ASAP7_75t_SL g846 ( 
.A(n_802),
.B(n_181),
.C(n_176),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_810),
.B(n_407),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_790),
.B(n_415),
.Y(n_848)
);

NAND2x2_ASAP7_75t_L g849 ( 
.A(n_791),
.B(n_445),
.Y(n_849)
);

OR2x6_ASAP7_75t_L g850 ( 
.A(n_783),
.B(n_666),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_783),
.B(n_621),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_R g852 ( 
.A(n_806),
.B(n_415),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_758),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_765),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_766),
.B(n_644),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_766),
.B(n_794),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_815),
.A2(n_798),
.B(n_775),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_817),
.A2(n_814),
.B1(n_804),
.B2(n_785),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_824),
.B(n_763),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_816),
.A2(n_779),
.B(n_801),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_848),
.A2(n_801),
.B(n_811),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_831),
.A2(n_753),
.B(n_789),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_829),
.A2(n_753),
.B(n_799),
.Y(n_863)
);

AOI33xp33_ASAP7_75t_L g864 ( 
.A1(n_842),
.A2(n_774),
.A3(n_781),
.B1(n_772),
.B2(n_770),
.B3(n_416),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_829),
.A2(n_786),
.B(n_778),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_840),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_R g867 ( 
.A(n_825),
.B(n_415),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_849),
.A2(n_835),
.B1(n_821),
.B2(n_820),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_821),
.B(n_812),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_856),
.B(n_793),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_833),
.A2(n_784),
.B(n_776),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_844),
.Y(n_872)
);

OR2x2_ASAP7_75t_SL g873 ( 
.A(n_856),
.B(n_795),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_851),
.A2(n_782),
.B(n_769),
.Y(n_874)
);

BUFx8_ASAP7_75t_L g875 ( 
.A(n_818),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_830),
.B(n_760),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_851),
.A2(n_788),
.B(n_756),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_855),
.A2(n_788),
.B(n_768),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_855),
.A2(n_752),
.B(n_797),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_819),
.B(n_787),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_850),
.A2(n_797),
.B(n_792),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_853),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_850),
.A2(n_416),
.B(n_401),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_836),
.Y(n_884)
);

OAI22xp33_ASAP7_75t_L g885 ( 
.A1(n_821),
.A2(n_592),
.B1(n_529),
.B2(n_585),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_850),
.A2(n_389),
.B(n_592),
.Y(n_886)
);

AOI21xp33_ASAP7_75t_L g887 ( 
.A1(n_822),
.A2(n_435),
.B(n_193),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_828),
.A2(n_389),
.B(n_408),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_832),
.A2(n_389),
.B(n_408),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_823),
.B(n_165),
.C(n_161),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_845),
.A2(n_408),
.B(n_529),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_838),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_818),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_846),
.A2(n_192),
.B(n_382),
.C(n_376),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_854),
.Y(n_895)
);

AO21x1_ASAP7_75t_L g896 ( 
.A1(n_839),
.A2(n_841),
.B(n_827),
.Y(n_896)
);

AOI21xp33_ASAP7_75t_L g897 ( 
.A1(n_847),
.A2(n_0),
.B(n_1),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_839),
.B(n_283),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_818),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_852),
.B(n_283),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_834),
.B(n_436),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_830),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_826),
.B(n_381),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_826),
.B(n_2),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_826),
.A2(n_391),
.B(n_388),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_837),
.B(n_2),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_843),
.A2(n_161),
.B(n_165),
.C(n_166),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_896),
.B(n_837),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_857),
.B(n_381),
.Y(n_909)
);

NAND2xp33_ASAP7_75t_SL g910 ( 
.A(n_867),
.B(n_166),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_874),
.B(n_381),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_862),
.B(n_381),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_861),
.B(n_381),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_864),
.B(n_3),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_876),
.B(n_3),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_868),
.B(n_431),
.Y(n_916)
);

NAND2xp33_ASAP7_75t_SL g917 ( 
.A(n_898),
.B(n_187),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_871),
.B(n_4),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_SL g919 ( 
.A(n_900),
.B(n_187),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_863),
.B(n_431),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_SL g921 ( 
.A(n_866),
.B(n_473),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_872),
.B(n_4),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_860),
.B(n_431),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_SL g924 ( 
.A(n_866),
.B(n_473),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_883),
.B(n_431),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_866),
.B(n_431),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_858),
.B(n_443),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_922),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_918),
.B(n_912),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_909),
.B(n_884),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_908),
.B(n_870),
.Y(n_931)
);

AOI21x1_ASAP7_75t_L g932 ( 
.A1(n_908),
.A2(n_869),
.B(n_879),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_915),
.B(n_869),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_927),
.A2(n_894),
.B(n_865),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_914),
.B(n_884),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_911),
.A2(n_873),
.B1(n_907),
.B2(n_890),
.Y(n_936)
);

BUFx12f_ASAP7_75t_L g937 ( 
.A(n_917),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_926),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_923),
.A2(n_891),
.B1(n_888),
.B2(n_889),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_913),
.B(n_882),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_916),
.A2(n_920),
.B(n_925),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_919),
.A2(n_897),
.B1(n_893),
.B2(n_885),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_921),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_924),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_910),
.Y(n_945)
);

NOR2x1_ASAP7_75t_L g946 ( 
.A(n_908),
.B(n_893),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_922),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_908),
.B(n_878),
.Y(n_948)
);

AO32x2_ASAP7_75t_L g949 ( 
.A1(n_908),
.A2(n_877),
.A3(n_892),
.B1(n_880),
.B2(n_859),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_918),
.B(n_895),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_915),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_922),
.Y(n_952)
);

INVx8_ASAP7_75t_L g953 ( 
.A(n_937),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_950),
.B(n_904),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_932),
.A2(n_881),
.B(n_902),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_951),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_946),
.A2(n_931),
.B(n_948),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_935),
.Y(n_958)
);

AND3x2_ASAP7_75t_L g959 ( 
.A(n_945),
.B(n_906),
.C(n_901),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_934),
.A2(n_887),
.B(n_886),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_954),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_953),
.Y(n_962)
);

INVx5_ASAP7_75t_SL g963 ( 
.A(n_953),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_962),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_961),
.A2(n_957),
.B1(n_930),
.B2(n_958),
.Y(n_965)
);

OAI221xp5_ASAP7_75t_L g966 ( 
.A1(n_965),
.A2(n_960),
.B1(n_936),
.B2(n_956),
.C(n_929),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_964),
.A2(n_955),
.B(n_960),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_967),
.Y(n_968)
);

O2A1O1Ixp5_ASAP7_75t_L g969 ( 
.A1(n_966),
.A2(n_936),
.B(n_944),
.C(n_943),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_968),
.B(n_963),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_969),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_971),
.A2(n_963),
.B1(n_950),
.B2(n_938),
.Y(n_972)
);

INVx5_ASAP7_75t_L g973 ( 
.A(n_970),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_973),
.Y(n_974)
);

BUFx12f_ASAP7_75t_L g975 ( 
.A(n_972),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_974),
.B(n_970),
.Y(n_976)
);

NAND2xp33_ASAP7_75t_R g977 ( 
.A(n_974),
.B(n_959),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_R g978 ( 
.A(n_975),
.B(n_5),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_976),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_977),
.B(n_928),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_978),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_981),
.B(n_947),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_979),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_983),
.B(n_980),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_982),
.B(n_949),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_SL g986 ( 
.A1(n_984),
.A2(n_952),
.B(n_942),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_985),
.B(n_933),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_987),
.B(n_941),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_986),
.B(n_940),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_988),
.B(n_942),
.Y(n_990)
);

NOR2x1_ASAP7_75t_L g991 ( 
.A(n_989),
.B(n_940),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_991),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_990),
.B(n_949),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_993),
.B(n_992),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_992),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_993),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_994),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_996),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_995),
.B(n_899),
.Y(n_999)
);

XOR2xp5_ASAP7_75t_L g1000 ( 
.A(n_999),
.B(n_5),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_998),
.B(n_6),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_1001),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_1000),
.Y(n_1003)
);

OAI211xp5_ASAP7_75t_SL g1004 ( 
.A1(n_1003),
.A2(n_997),
.B(n_7),
.C(n_8),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_1002),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_1005),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_1004),
.B(n_6),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1007),
.B(n_7),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1006),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_1009),
.A2(n_875),
.B1(n_939),
.B2(n_899),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1008),
.B(n_8),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1011),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1010),
.Y(n_1013)
);

OAI32xp33_ASAP7_75t_L g1014 ( 
.A1(n_1011),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1012),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1013),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1014),
.B(n_10),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1017),
.Y(n_1018)
);

OAI221xp5_ASAP7_75t_L g1019 ( 
.A1(n_1016),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1018),
.B(n_1015),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1019),
.B(n_15),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_1020),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1021),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1022),
.B(n_949),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_L g1025 ( 
.A(n_1023),
.B(n_875),
.C(n_16),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_1025),
.B(n_17),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_1024),
.Y(n_1027)
);

AOI221xp5_ASAP7_75t_L g1028 ( 
.A1(n_1027),
.A2(n_319),
.B1(n_18),
.B2(n_19),
.C(n_20),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_1026),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_1029),
.B(n_1028),
.Y(n_1030)
);

NAND4xp25_ASAP7_75t_SL g1031 ( 
.A(n_1029),
.B(n_17),
.C(n_18),
.D(n_19),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_1029),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_1032)
);

XOR2xp5_ASAP7_75t_L g1033 ( 
.A(n_1030),
.B(n_21),
.Y(n_1033)
);

OAI221xp5_ASAP7_75t_L g1034 ( 
.A1(n_1032),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.C(n_25),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1031),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1035),
.B(n_26),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1034),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_1037)
);

NOR2x1_ASAP7_75t_L g1038 ( 
.A(n_1037),
.B(n_1033),
.Y(n_1038)
);

NOR2x1_ASAP7_75t_L g1039 ( 
.A(n_1036),
.B(n_27),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_SL g1040 ( 
.A1(n_1038),
.A2(n_29),
.B(n_30),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1039),
.B(n_29),
.Y(n_1041)
);

AOI211x1_ASAP7_75t_L g1042 ( 
.A1(n_1041),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_1040),
.B(n_32),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_R g1044 ( 
.A(n_1043),
.B(n_33),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_1042),
.B(n_319),
.Y(n_1045)
);

INVx3_ASAP7_75t_SL g1046 ( 
.A(n_1045),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_1044),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_1046),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1047),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1047),
.Y(n_1050)
);

AO22x2_ASAP7_75t_L g1051 ( 
.A1(n_1049),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_1048),
.Y(n_1052)
);

AND3x2_ASAP7_75t_L g1053 ( 
.A(n_1050),
.B(n_34),
.C(n_35),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_1052),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1051),
.A2(n_36),
.B(n_37),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1054),
.Y(n_1056)
);

XNOR2xp5_ASAP7_75t_L g1057 ( 
.A(n_1055),
.B(n_1053),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1056),
.A2(n_1057),
.B1(n_899),
.B2(n_37),
.Y(n_1058)
);

NOR2x2_ASAP7_75t_L g1059 ( 
.A(n_1056),
.B(n_38),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_1059),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1058),
.Y(n_1061)
);

XOR2xp5_ASAP7_75t_L g1062 ( 
.A(n_1060),
.B(n_38),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_1061),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1063),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1062),
.A2(n_443),
.B1(n_319),
.B2(n_385),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_319),
.B1(n_443),
.B2(n_385),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1065),
.A2(n_443),
.B1(n_385),
.B2(n_393),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_1064),
.A2(n_443),
.B1(n_393),
.B2(n_43),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_SL g1069 ( 
.A1(n_1067),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_1069)
);

XOR2xp5_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_1066),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1067),
.A2(n_393),
.B1(n_905),
.B2(n_48),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1067),
.Y(n_1072)
);

AO21x2_ASAP7_75t_L g1073 ( 
.A1(n_1072),
.A2(n_46),
.B(n_47),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_1070),
.B(n_49),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1069),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_1075),
.Y(n_1076)
);

OAI222xp33_ASAP7_75t_L g1077 ( 
.A1(n_1074),
.A2(n_1071),
.B1(n_51),
.B2(n_52),
.C1(n_55),
.C2(n_57),
.Y(n_1077)
);

XNOR2xp5_ASAP7_75t_L g1078 ( 
.A(n_1073),
.B(n_50),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1076),
.A2(n_58),
.B(n_60),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1078),
.A2(n_61),
.B(n_62),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1077),
.B(n_63),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1076),
.B(n_65),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1076),
.A2(n_595),
.B1(n_903),
.B2(n_71),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1076),
.B(n_69),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1076),
.B(n_70),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1076),
.A2(n_72),
.B(n_73),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1076),
.A2(n_74),
.B(n_75),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1076),
.A2(n_76),
.B(n_77),
.Y(n_1088)
);

AO21x2_ASAP7_75t_L g1089 ( 
.A1(n_1076),
.A2(n_79),
.B(n_80),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1076),
.A2(n_82),
.B(n_83),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1081),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_SL g1092 ( 
.A1(n_1080),
.A2(n_87),
.B(n_89),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1088),
.Y(n_1093)
);

AOI222xp33_ASAP7_75t_L g1094 ( 
.A1(n_1084),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.C1(n_94),
.C2(n_95),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1085),
.A2(n_96),
.B(n_97),
.Y(n_1095)
);

XNOR2xp5_ASAP7_75t_L g1096 ( 
.A(n_1082),
.B(n_99),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1079),
.A2(n_101),
.B(n_102),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1086),
.A2(n_103),
.B(n_105),
.Y(n_1098)
);

OAI31xp33_ASAP7_75t_SL g1099 ( 
.A1(n_1089),
.A2(n_106),
.A3(n_107),
.B(n_108),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1093),
.A2(n_1087),
.B(n_1083),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_1091),
.A2(n_1090),
.B(n_111),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1097),
.A2(n_595),
.B1(n_113),
.B2(n_114),
.Y(n_1102)
);

AO21x1_ASAP7_75t_L g1103 ( 
.A1(n_1098),
.A2(n_109),
.B(n_116),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_SL g1104 ( 
.A1(n_1092),
.A2(n_117),
.B(n_118),
.Y(n_1104)
);

AO21x2_ASAP7_75t_L g1105 ( 
.A1(n_1096),
.A2(n_120),
.B(n_121),
.Y(n_1105)
);

AO21x2_ASAP7_75t_L g1106 ( 
.A1(n_1099),
.A2(n_122),
.B(n_124),
.Y(n_1106)
);

AOI222xp33_ASAP7_75t_L g1107 ( 
.A1(n_1100),
.A2(n_1106),
.B1(n_1104),
.B2(n_1101),
.C1(n_1103),
.C2(n_1102),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1105),
.A2(n_1095),
.B1(n_1094),
.B2(n_128),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1100),
.A2(n_125),
.B1(n_126),
.B2(n_129),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1100),
.A2(n_595),
.B1(n_482),
.B2(n_481),
.Y(n_1110)
);

OAI211xp5_ASAP7_75t_L g1111 ( 
.A1(n_1107),
.A2(n_130),
.B(n_132),
.C(n_133),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_1108),
.Y(n_1112)
);

OAI321xp33_ASAP7_75t_L g1113 ( 
.A1(n_1112),
.A2(n_1109),
.A3(n_1110),
.B1(n_136),
.B2(n_137),
.C(n_138),
.Y(n_1113)
);

OAI221xp5_ASAP7_75t_R g1114 ( 
.A1(n_1113),
.A2(n_1111),
.B1(n_135),
.B2(n_140),
.C(n_141),
.Y(n_1114)
);

AOI221xp5_ASAP7_75t_L g1115 ( 
.A1(n_1114),
.A2(n_134),
.B1(n_142),
.B2(n_143),
.C(n_144),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_145),
.B(n_146),
.Y(n_1116)
);

AOI211xp5_ASAP7_75t_L g1117 ( 
.A1(n_1116),
.A2(n_147),
.B(n_148),
.C(n_150),
.Y(n_1117)
);

AOI211xp5_ASAP7_75t_L g1118 ( 
.A1(n_1117),
.A2(n_151),
.B(n_155),
.C(n_157),
.Y(n_1118)
);


endmodule