module fake_netlist_6_1684_n_1915 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1915);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1915;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_70),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_50),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_27),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_84),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_28),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_189),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_52),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_80),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_69),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_64),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_49),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_32),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_36),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_100),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_86),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_4),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_0),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_3),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_42),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_39),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_2),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_46),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_58),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_103),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_154),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_92),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_51),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_48),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_109),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_81),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_137),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_90),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_1),
.Y(n_229)
);

BUFx8_ASAP7_75t_SL g230 ( 
.A(n_43),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_117),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_62),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_56),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_146),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_39),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_145),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_51),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_168),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_101),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_54),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_17),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_0),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_77),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_29),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_149),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_188),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_12),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_185),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_2),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_127),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_173),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_74),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_34),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_187),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_152),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_114),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_119),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_11),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_122),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_19),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_158),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_45),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_82),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_45),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_132),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_27),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_11),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_53),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_88),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_87),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_155),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_68),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_163),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_10),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_110),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_28),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_89),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_17),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_26),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_43),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_176),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_9),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_10),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_40),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_112),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_139),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_160),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_46),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_175),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_124),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_31),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_12),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_159),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_174),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_75),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_26),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_178),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_50),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_44),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_186),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_99),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_107),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_1),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_5),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_57),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_115),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_19),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_104),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_66),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_65),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_6),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_140),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_147),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_142),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_35),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_49),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_134),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_136),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_183),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_22),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_166),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_76),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_130),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_78),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_47),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_22),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_16),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_105),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_29),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_116),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_85),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_71),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_13),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_35),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_16),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_121),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_55),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_40),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_182),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_108),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_96),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_170),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_44),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_41),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_177),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_123),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_32),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_164),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_6),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_150),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_14),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_4),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_94),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_60),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_113),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_20),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_20),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_38),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_79),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_73),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_143),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_61),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_24),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_3),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_184),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_128),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_133),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_42),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_59),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_18),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_8),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_30),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_34),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_15),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_365),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_203),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_203),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_230),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_338),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_229),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_234),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_338),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_220),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_226),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_242),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_216),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_242),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_285),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_285),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_293),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_229),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_224),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_192),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_293),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_221),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_250),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_229),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_351),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_228),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_281),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_254),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_265),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_269),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_279),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_231),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_290),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_232),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_320),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_281),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_244),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_246),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_247),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_324),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_249),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_252),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_192),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_235),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_255),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_193),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_258),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_377),
.Y(n_429)
);

BUFx2_ASAP7_75t_SL g430 ( 
.A(n_289),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_282),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_282),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_270),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_257),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_271),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_329),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_329),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_281),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_191),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_200),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_200),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_325),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_325),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_239),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_198),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_206),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_212),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_219),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_273),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_274),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_225),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_251),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_191),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_257),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_301),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_193),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_283),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_227),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_233),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_301),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_257),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_240),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_215),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_266),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_301),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_287),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_288),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_241),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_208),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_223),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_272),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_253),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g473 ( 
.A1(n_434),
.A2(n_264),
.B(n_260),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_289),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_445),
.B(n_223),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_454),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_310),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_454),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_310),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g482 ( 
.A1(n_461),
.A2(n_295),
.B(n_278),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_461),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_440),
.A2(n_303),
.B(n_296),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_430),
.B(n_190),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_346),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_446),
.B(n_346),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_440),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_312),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_421),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_396),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_399),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_441),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_441),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_426),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_396),
.Y(n_500)
);

OA21x2_ASAP7_75t_L g501 ( 
.A1(n_442),
.A2(n_332),
.B(n_321),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_447),
.B(n_335),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_447),
.B(n_341),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_443),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_400),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_443),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_380),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_418),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_430),
.B(n_190),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_387),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_448),
.B(n_451),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_388),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_423),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_384),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_418),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_448),
.B(n_358),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_456),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_451),
.B(n_194),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_463),
.A2(n_309),
.B1(n_375),
.B2(n_298),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_380),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_458),
.B(n_363),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_R g525 ( 
.A(n_456),
.B(n_378),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_458),
.B(n_194),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_404),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_406),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_472),
.A2(n_262),
.B(n_257),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_381),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_406),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_381),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_459),
.B(n_257),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_407),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_459),
.B(n_262),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_462),
.B(n_196),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_383),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_407),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_462),
.B(n_262),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_408),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_383),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_444),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_408),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_386),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_386),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_379),
.B(n_208),
.Y(n_546)
);

BUFx8_ASAP7_75t_L g547 ( 
.A(n_389),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_405),
.B(n_208),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_411),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_468),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_410),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_493),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_550),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_479),
.A2(n_385),
.B1(n_472),
.B2(n_468),
.Y(n_554)
);

AND3x2_ASAP7_75t_L g555 ( 
.A(n_517),
.B(n_243),
.C(n_276),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_479),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_488),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_492),
.A2(n_412),
.B1(n_415),
.B2(n_467),
.Y(n_558)
);

INVx8_ASAP7_75t_L g559 ( 
.A(n_513),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_479),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_495),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_516),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_550),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_550),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_550),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_493),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_514),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_485),
.B(n_416),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_485),
.B(n_417),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_512),
.B(n_419),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_488),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_520),
.B(n_414),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_514),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_481),
.B(n_493),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_515),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_514),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_520),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_535),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_488),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_535),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_475),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_478),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_481),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_480),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_512),
.B(n_420),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_478),
.Y(n_587)
);

BUFx6f_ASAP7_75t_SL g588 ( 
.A(n_476),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_507),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_507),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_535),
.B(n_262),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_480),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_492),
.A2(n_469),
.B1(n_474),
.B2(n_438),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_483),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_527),
.B(n_425),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_533),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_517),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_551),
.B(n_427),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_483),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_488),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_481),
.B(n_433),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_474),
.B(n_435),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_530),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_476),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_507),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_506),
.B(n_449),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_521),
.B(n_450),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_530),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_506),
.B(n_391),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_533),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_477),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_476),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_498),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_530),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_533),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_530),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_498),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_521),
.B(n_457),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_530),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_476),
.B(n_466),
.Y(n_622)
);

AOI21x1_ASAP7_75t_L g623 ( 
.A1(n_529),
.A2(n_482),
.B(n_473),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_533),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_473),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_533),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_539),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_526),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_539),
.Y(n_629)
);

AO21x2_ASAP7_75t_L g630 ( 
.A1(n_529),
.A2(n_359),
.B(n_422),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_542),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_530),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_545),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_476),
.B(n_202),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_539),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_488),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_486),
.B(n_391),
.Y(n_637)
);

OAI21xp33_ASAP7_75t_SL g638 ( 
.A1(n_548),
.A2(n_393),
.B(n_392),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_526),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_545),
.Y(n_640)
);

OAI21xp33_ASAP7_75t_SL g641 ( 
.A1(n_546),
.A2(n_393),
.B(n_392),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_539),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_536),
.B(n_455),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_486),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_545),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_478),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_545),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_488),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_525),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_545),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_536),
.B(n_465),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_489),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_545),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_525),
.A2(n_322),
.B1(n_343),
.B2(n_316),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_539),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_545),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_473),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_478),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_496),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_528),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_489),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_496),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_531),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_496),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_502),
.B(n_237),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_488),
.Y(n_666)
);

INVxp33_ASAP7_75t_L g667 ( 
.A(n_522),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_507),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_486),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_SL g670 ( 
.A(n_522),
.B(n_238),
.Y(n_670)
);

AO21x2_ASAP7_75t_L g671 ( 
.A1(n_529),
.A2(n_424),
.B(n_413),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_507),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_507),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_547),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_531),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_507),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_534),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_547),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_509),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_509),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_534),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_547),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_547),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_538),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_509),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_538),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_540),
.Y(n_687)
);

INVx8_ASAP7_75t_L g688 ( 
.A(n_489),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_509),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_509),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_489),
.B(n_395),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_487),
.Y(n_692)
);

BUFx10_ASAP7_75t_L g693 ( 
.A(n_489),
.Y(n_693)
);

INVx8_ASAP7_75t_L g694 ( 
.A(n_519),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_509),
.Y(n_695)
);

NOR2x1p5_ASAP7_75t_L g696 ( 
.A(n_540),
.B(n_382),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_543),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_509),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_508),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_473),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_502),
.B(n_302),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_628),
.B(n_311),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_556),
.B(n_519),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_556),
.B(n_519),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_560),
.B(n_519),
.Y(n_705)
);

NOR2xp67_ASAP7_75t_L g706 ( 
.A(n_598),
.B(n_401),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_625),
.A2(n_482),
.B(n_473),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_560),
.B(n_519),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_613),
.B(n_460),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_692),
.B(n_487),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_SL g711 ( 
.A(n_576),
.B(n_452),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_552),
.B(n_487),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_584),
.B(n_524),
.Y(n_713)
);

NOR2x2_ASAP7_75t_L g714 ( 
.A(n_670),
.B(n_464),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_628),
.A2(n_471),
.B1(n_524),
.B2(n_503),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_584),
.B(n_524),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_660),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_609),
.B(n_524),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_620),
.B(n_524),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_644),
.B(n_394),
.Y(n_720)
);

OAI21xp33_ASAP7_75t_L g721 ( 
.A1(n_554),
.A2(n_398),
.B(n_394),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_597),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_644),
.B(n_639),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_639),
.B(n_262),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_601),
.B(n_504),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_575),
.B(n_504),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_608),
.B(n_504),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_569),
.B(n_504),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_575),
.B(n_504),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_579),
.B(n_502),
.Y(n_730)
);

INVxp33_ASAP7_75t_SL g731 ( 
.A(n_654),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_552),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_568),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_579),
.B(n_503),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_568),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_649),
.B(n_196),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_581),
.B(n_503),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_566),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_567),
.A2(n_501),
.B1(n_484),
.B2(n_482),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_567),
.A2(n_501),
.B1(n_484),
.B2(n_482),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_649),
.B(n_199),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_597),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_570),
.B(n_199),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_663),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_581),
.B(n_497),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_663),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_691),
.A2(n_497),
.B(n_499),
.C(n_543),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_675),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_566),
.B(n_549),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_661),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_643),
.B(n_402),
.C(n_398),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_582),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_582),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_574),
.B(n_577),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_661),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_574),
.B(n_497),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_577),
.B(n_497),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_586),
.B(n_602),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_622),
.A2(n_308),
.B1(n_327),
.B2(n_323),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_657),
.A2(n_611),
.B1(n_700),
.B2(n_667),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_675),
.B(n_677),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_677),
.B(n_499),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_700),
.B(n_328),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_578),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_613),
.B(n_402),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_578),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_583),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_681),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_596),
.A2(n_499),
.B(n_549),
.C(n_541),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_681),
.B(n_499),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_684),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_583),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_684),
.B(n_484),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_686),
.B(n_484),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_686),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_687),
.B(n_484),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_573),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_619),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_700),
.B(n_328),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_687),
.B(n_501),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_619),
.B(n_403),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_669),
.B(n_201),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_697),
.B(n_501),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_583),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_607),
.B(n_403),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_688),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_611),
.A2(n_501),
.B1(n_482),
.B2(n_245),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_697),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_596),
.B(n_508),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_700),
.B(n_328),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_700),
.B(n_652),
.Y(n_791)
);

AND2x6_ASAP7_75t_L g792 ( 
.A(n_612),
.B(n_328),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_612),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_634),
.A2(n_354),
.B1(n_291),
.B2(n_292),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_652),
.B(n_328),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_617),
.B(n_508),
.Y(n_796)
);

INVxp67_ASAP7_75t_SL g797 ( 
.A(n_666),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_617),
.A2(n_277),
.B1(n_356),
.B2(n_345),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_651),
.B(n_201),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_615),
.B(n_431),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_624),
.B(n_523),
.Y(n_801)
);

OR2x6_ASAP7_75t_L g802 ( 
.A(n_559),
.B(n_431),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_571),
.B(n_207),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_665),
.B(n_207),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_652),
.B(n_345),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_624),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_626),
.A2(n_345),
.B1(n_195),
.B2(n_204),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_558),
.B(n_236),
.C(n_222),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_627),
.A2(n_218),
.B1(n_214),
.B2(n_373),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_627),
.B(n_523),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_587),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_561),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_701),
.B(n_214),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_629),
.B(n_523),
.Y(n_814)
);

BUFx5_ASAP7_75t_L g815 ( 
.A(n_605),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_587),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_629),
.B(n_532),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_635),
.B(n_532),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_693),
.B(n_345),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_635),
.B(n_532),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_637),
.A2(n_411),
.B(n_413),
.C(n_428),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_638),
.B(n_218),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_638),
.B(n_364),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_642),
.B(n_537),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_641),
.B(n_364),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_637),
.Y(n_826)
);

AND2x6_ASAP7_75t_SL g827 ( 
.A(n_561),
.B(n_428),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_655),
.A2(n_588),
.B1(n_641),
.B2(n_593),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_573),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_588),
.A2(n_366),
.B1(n_369),
.B2(n_373),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_559),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_553),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_605),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_588),
.A2(n_350),
.B1(n_297),
.B2(n_307),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_674),
.B(n_366),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_563),
.B(n_541),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_562),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_L g838 ( 
.A(n_688),
.B(n_299),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_563),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_666),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_564),
.B(n_541),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_565),
.B(n_544),
.Y(n_842)
);

BUFx12f_ASAP7_75t_SL g843 ( 
.A(n_559),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_565),
.B(n_544),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_693),
.B(n_345),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_587),
.B(n_544),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_646),
.B(n_490),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_585),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_693),
.B(n_304),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_631),
.B(n_432),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_605),
.B(n_313),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_646),
.B(n_490),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_646),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_614),
.B(n_314),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_614),
.B(n_317),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_658),
.B(n_491),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_614),
.B(n_318),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_595),
.B(n_369),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_658),
.B(n_690),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_592),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_658),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_766),
.B(n_559),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_812),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_760),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_758),
.B(n_725),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_755),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_755),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_793),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_755),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_806),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_758),
.B(n_688),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_832),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_763),
.A2(n_623),
.B(n_668),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_755),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_722),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_778),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_839),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_709),
.B(n_696),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_750),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_743),
.B(n_694),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_743),
.B(n_694),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_848),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_785),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_727),
.B(n_694),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_750),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_727),
.B(n_718),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_719),
.B(n_659),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_710),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_760),
.A2(n_696),
.B1(n_683),
.B2(n_591),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_850),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_860),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_728),
.B(n_815),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_728),
.B(n_576),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_763),
.A2(n_623),
.B(n_668),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_SL g895 ( 
.A(n_798),
.B(n_678),
.C(n_674),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_712),
.B(n_682),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_787),
.A2(n_630),
.B1(n_671),
.B2(n_591),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_777),
.B(n_555),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_800),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_712),
.B(n_682),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_SL g901 ( 
.A1(n_804),
.A2(n_672),
.B(n_698),
.C(n_673),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_764),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_804),
.B(n_659),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_843),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_787),
.A2(n_678),
.B1(n_698),
.B2(n_672),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_813),
.B(n_662),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_765),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_717),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_733),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_735),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_731),
.B(n_248),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_742),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_829),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_815),
.B(n_673),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_826),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_752),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_837),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_702),
.B(n_259),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_813),
.B(n_662),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_767),
.Y(n_920)
);

O2A1O1Ixp5_ASAP7_75t_L g921 ( 
.A1(n_779),
.A2(n_599),
.B(n_594),
.C(n_664),
.Y(n_921)
);

NOR2x1p5_ASAP7_75t_L g922 ( 
.A(n_831),
.B(n_195),
.Y(n_922)
);

AOI21xp33_ASAP7_75t_L g923 ( 
.A1(n_803),
.A2(n_630),
.B(n_263),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_772),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_786),
.B(n_690),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_754),
.B(n_664),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_807),
.A2(n_630),
.B1(n_671),
.B2(n_591),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_702),
.B(n_699),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_753),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_833),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_781),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_802),
.B(n_429),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_784),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_732),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_SL g935 ( 
.A1(n_798),
.A2(n_217),
.B1(n_213),
.B2(n_211),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_744),
.B(n_699),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_746),
.B(n_690),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_811),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_723),
.B(n_261),
.Y(n_939)
);

BUFx8_ASAP7_75t_L g940 ( 
.A(n_720),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_748),
.B(n_695),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_736),
.B(n_267),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_768),
.B(n_695),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_749),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_771),
.B(n_695),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_815),
.B(n_676),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_779),
.A2(n_572),
.B(n_557),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_816),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_775),
.B(n_666),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_833),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_R g951 ( 
.A(n_711),
.B(n_370),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_732),
.Y(n_952)
);

NAND2xp33_ASAP7_75t_L g953 ( 
.A(n_815),
.B(n_591),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_788),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_730),
.B(n_676),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_853),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_815),
.B(n_680),
.Y(n_957)
);

NAND2xp33_ASAP7_75t_SL g958 ( 
.A(n_807),
.B(n_370),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_738),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_782),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_847),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_749),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_815),
.B(n_680),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_802),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_703),
.A2(n_685),
.B1(n_689),
.B2(n_604),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_861),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_852),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_856),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_756),
.Y(n_969)
);

NOR3xp33_ASAP7_75t_SL g970 ( 
.A(n_741),
.B(n_204),
.C(n_197),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_714),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_734),
.B(n_685),
.Y(n_972)
);

O2A1O1Ixp5_ASAP7_75t_L g973 ( 
.A1(n_790),
.A2(n_689),
.B(n_610),
.C(n_618),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_738),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_715),
.B(n_268),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_782),
.B(n_275),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_737),
.B(n_603),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_802),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_827),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_846),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_828),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_757),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_786),
.B(n_557),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_R g984 ( 
.A(n_858),
.B(n_371),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_859),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_799),
.B(n_803),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_704),
.A2(n_705),
.B1(n_713),
.B2(n_708),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_761),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_789),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_792),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_792),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_796),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_724),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_706),
.B(n_371),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_801),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_799),
.B(n_280),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_716),
.B(n_603),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_751),
.B(n_429),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_822),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_858),
.B(n_436),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_762),
.Y(n_1001)
);

AND2x4_ASAP7_75t_SL g1002 ( 
.A(n_834),
.B(n_256),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_759),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_726),
.B(n_604),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_823),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_729),
.B(n_610),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_R g1007 ( 
.A(n_838),
.B(n_326),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_724),
.B(n_284),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_808),
.B(n_286),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_745),
.B(n_616),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_773),
.B(n_616),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_825),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_835),
.B(n_436),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_770),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_792),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_809),
.B(n_294),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_797),
.B(n_618),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_810),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_814),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_774),
.A2(n_671),
.B1(n_591),
.B2(n_197),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_791),
.Y(n_1021)
);

INVxp33_ASAP7_75t_L g1022 ( 
.A(n_721),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_830),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_792),
.Y(n_1024)
);

OR2x6_ASAP7_75t_SL g1025 ( 
.A(n_776),
.B(n_205),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_792),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_840),
.B(n_621),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_817),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_818),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_820),
.Y(n_1030)
);

AND2x2_ASAP7_75t_SL g1031 ( 
.A(n_780),
.B(n_621),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_824),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_821),
.B(n_437),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_R g1034 ( 
.A(n_849),
.B(n_205),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_794),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_L g1036 ( 
.A(n_849),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_790),
.B(n_707),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_747),
.B(n_791),
.Y(n_1038)
);

AND2x4_ASAP7_75t_SL g1039 ( 
.A(n_739),
.B(n_256),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_851),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_783),
.B(n_739),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_868),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_884),
.A2(n_886),
.B(n_871),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_865),
.B(n_857),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_870),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1037),
.A2(n_740),
.B(n_769),
.Y(n_1046)
);

BUFx4_ASAP7_75t_SL g1047 ( 
.A(n_904),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_986),
.B(n_851),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_986),
.A2(n_857),
.B1(n_855),
.B2(n_854),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_960),
.B(n_854),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_863),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_L g1052 ( 
.A1(n_996),
.A2(n_855),
.B(n_845),
.C(n_795),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_883),
.B(n_437),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_917),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_866),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_908),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_864),
.A2(n_740),
.B1(n_845),
.B2(n_819),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_875),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_996),
.A2(n_819),
.B(n_805),
.C(n_795),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_866),
.Y(n_1060)
);

INVx3_ASAP7_75t_SL g1061 ( 
.A(n_971),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_960),
.B(n_836),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1036),
.B(n_841),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_918),
.A2(n_844),
.B(n_842),
.C(n_656),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_918),
.A2(n_632),
.B(n_656),
.C(n_653),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_864),
.A2(n_217),
.B1(n_210),
.B2(n_211),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_911),
.B(n_491),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_988),
.B(n_633),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_976),
.A2(n_633),
.B(n_653),
.C(n_650),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_866),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_976),
.A2(n_640),
.B(n_650),
.C(n_647),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_907),
.B(n_640),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_892),
.A2(n_600),
.B(n_580),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_951),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_866),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_907),
.B(n_1018),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_867),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_954),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_876),
.Y(n_1079)
);

O2A1O1Ixp5_ASAP7_75t_L g1080 ( 
.A1(n_923),
.A2(n_647),
.B(n_645),
.C(n_557),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_911),
.B(n_494),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_877),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1036),
.B(n_334),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_897),
.A2(n_209),
.B1(n_210),
.B2(n_213),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_940),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_872),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_981),
.A2(n_591),
.B1(n_256),
.B2(n_352),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1032),
.B(n_645),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_936),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_880),
.A2(n_600),
.B(n_572),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_896),
.B(n_494),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1008),
.A2(n_349),
.B(n_357),
.C(n_344),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_940),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_1009),
.A2(n_510),
.B(n_511),
.C(n_500),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_888),
.B(n_500),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1040),
.B(n_336),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_881),
.A2(n_580),
.B(n_572),
.Y(n_1097)
);

OAI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_1016),
.A2(n_1022),
.B(n_975),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_887),
.A2(n_600),
.B(n_636),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1016),
.A2(n_510),
.B(n_511),
.C(n_505),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1009),
.A2(n_518),
.B(n_300),
.C(n_305),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_867),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_867),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_888),
.B(n_518),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_989),
.B(n_340),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_953),
.A2(n_636),
.B(n_679),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_992),
.B(n_589),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1023),
.A2(n_348),
.B(n_306),
.C(n_315),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1041),
.A2(n_947),
.B(n_1004),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_931),
.B(n_589),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_890),
.B(n_319),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_995),
.B(n_589),
.Y(n_1112)
);

NAND2x1p5_ASAP7_75t_L g1113 ( 
.A(n_867),
.B(n_636),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_896),
.B(n_589),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_913),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_890),
.B(n_330),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_899),
.B(n_331),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_974),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_869),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_869),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_899),
.B(n_589),
.Y(n_1121)
);

NOR3xp33_ASAP7_75t_L g1122 ( 
.A(n_975),
.B(n_895),
.C(n_1034),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_869),
.B(n_590),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_882),
.Y(n_1124)
);

AO32x2_ASAP7_75t_L g1125 ( 
.A1(n_905),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_909),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1041),
.A2(n_679),
.B(n_606),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_900),
.B(n_590),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_934),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_869),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_874),
.Y(n_1131)
);

NOR2xp67_ASAP7_75t_L g1132 ( 
.A(n_862),
.B(n_63),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_874),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_897),
.A2(n_209),
.B1(n_362),
.B2(n_367),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_983),
.A2(n_679),
.B(n_606),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_874),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_R g1137 ( 
.A(n_1003),
.B(n_362),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_891),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_910),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1019),
.B(n_679),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_927),
.A2(n_367),
.B1(n_368),
.B2(n_372),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_902),
.B(n_360),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1008),
.A2(n_361),
.B(n_339),
.C(n_342),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_902),
.B(n_337),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_969),
.B(n_679),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_874),
.Y(n_1146)
);

CKINVDCx8_ASAP7_75t_R g1147 ( 
.A(n_979),
.Y(n_1147)
);

NOR2x1_ASAP7_75t_L g1148 ( 
.A(n_893),
.B(n_590),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_983),
.A2(n_606),
.B(n_590),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_873),
.A2(n_606),
.B(n_590),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_893),
.A2(n_606),
.B(n_98),
.C(n_148),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_916),
.Y(n_1152)
);

INVx5_ASAP7_75t_L g1153 ( 
.A(n_932),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_912),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_894),
.A2(n_648),
.B(n_97),
.Y(n_1155)
);

INVx6_ASAP7_75t_L g1156 ( 
.A(n_934),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_929),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_927),
.A2(n_378),
.B1(n_372),
.B2(n_368),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_920),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_914),
.A2(n_648),
.B(n_93),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_914),
.A2(n_648),
.B(n_91),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_946),
.A2(n_648),
.B(n_95),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_879),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1020),
.A2(n_355),
.B1(n_353),
.B2(n_347),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_939),
.B(n_1013),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_946),
.A2(n_648),
.B(n_72),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_912),
.B(n_13),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_879),
.Y(n_1168)
);

BUFx8_ASAP7_75t_L g1169 ( 
.A(n_878),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_920),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_957),
.A2(n_648),
.B(n_83),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_952),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_957),
.A2(n_67),
.B(n_180),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_982),
.B(n_14),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_942),
.B(n_15),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_942),
.B(n_18),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_915),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_961),
.B(n_21),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_939),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1020),
.A2(n_23),
.B1(n_25),
.B2(n_30),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_958),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_993),
.A2(n_33),
.B(n_36),
.C(n_37),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_924),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_879),
.B(n_885),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_967),
.B(n_928),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_993),
.A2(n_125),
.B1(n_179),
.B2(n_172),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_879),
.B(n_118),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_963),
.A2(n_111),
.B(n_171),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_968),
.B(n_37),
.Y(n_1189)
);

CKINVDCx16_ASAP7_75t_R g1190 ( 
.A(n_951),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_915),
.B(n_38),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1028),
.B(n_41),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_885),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_999),
.A2(n_129),
.B1(n_167),
.B2(n_162),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_L g1195 ( 
.A1(n_901),
.A2(n_106),
.B(n_157),
.C(n_151),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1165),
.B(n_1000),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1048),
.A2(n_1038),
.B(n_987),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1098),
.A2(n_1012),
.B(n_1005),
.C(n_1035),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1098),
.B(n_952),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_1175),
.B(n_1176),
.C(n_1049),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1043),
.A2(n_1109),
.B(n_1097),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1118),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1090),
.A2(n_903),
.B(n_906),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1127),
.A2(n_973),
.B(n_921),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1079),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1069),
.A2(n_965),
.A3(n_919),
.B(n_901),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1067),
.B(n_959),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1185),
.B(n_1001),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1071),
.A2(n_955),
.A3(n_972),
.B(n_977),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1193),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_SL g1211 ( 
.A(n_1180),
.B(n_935),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1044),
.A2(n_1031),
.B(n_1006),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1065),
.A2(n_1010),
.A3(n_1014),
.B(n_926),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1193),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1059),
.A2(n_950),
.B(n_930),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1073),
.A2(n_963),
.B(n_997),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1081),
.B(n_959),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1052),
.A2(n_997),
.B(n_1006),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1050),
.A2(n_1002),
.B(n_889),
.C(n_1039),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1135),
.A2(n_1011),
.B(n_925),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1193),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1055),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1076),
.A2(n_930),
.B1(n_950),
.B2(n_885),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1101),
.A2(n_898),
.B(n_970),
.C(n_1030),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1064),
.A2(n_1031),
.B(n_985),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1057),
.A2(n_925),
.B(n_990),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1055),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1062),
.B(n_1030),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1179),
.A2(n_994),
.B(n_898),
.C(n_970),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1057),
.A2(n_980),
.A3(n_943),
.B(n_941),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1089),
.A2(n_885),
.B1(n_934),
.B2(n_1021),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1149),
.A2(n_937),
.B(n_945),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1055),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1056),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_SL g1235 ( 
.A1(n_1187),
.A2(n_949),
.B(n_978),
.C(n_964),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1095),
.B(n_1029),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1058),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1155),
.A2(n_1099),
.B(n_1106),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1104),
.B(n_962),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1046),
.A2(n_1017),
.B(n_1027),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1192),
.A2(n_990),
.A3(n_1026),
.B(n_956),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1154),
.B(n_900),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1195),
.A2(n_966),
.B(n_948),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1046),
.A2(n_938),
.B(n_933),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1080),
.A2(n_1015),
.B(n_1024),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1070),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1122),
.A2(n_944),
.B(n_998),
.C(n_1021),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1078),
.B(n_984),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_SL g1249 ( 
.A1(n_1173),
.A2(n_1026),
.B(n_1021),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1063),
.A2(n_1021),
.B(n_1024),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1160),
.A2(n_1015),
.B(n_991),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1082),
.B(n_984),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1124),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1070),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1051),
.Y(n_1255)
);

BUFx8_ASAP7_75t_L g1256 ( 
.A(n_1085),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_SL g1257 ( 
.A1(n_1182),
.A2(n_991),
.B(n_1025),
.C(n_1007),
.Y(n_1257)
);

INVx3_ASAP7_75t_SL g1258 ( 
.A(n_1054),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1161),
.A2(n_922),
.B(n_1007),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1108),
.A2(n_998),
.B(n_934),
.C(n_932),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1181),
.A2(n_932),
.B1(n_1033),
.B2(n_52),
.Y(n_1261)
);

NAND2xp33_ASAP7_75t_L g1262 ( 
.A(n_1174),
.B(n_1033),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1115),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1117),
.B(n_1033),
.Y(n_1264)
);

AOI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1148),
.A2(n_181),
.B(n_102),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1162),
.A2(n_126),
.B(n_135),
.Y(n_1266)
);

AO21x1_ASAP7_75t_L g1267 ( 
.A1(n_1178),
.A2(n_47),
.B(n_48),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1151),
.A2(n_53),
.B(n_1088),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1166),
.A2(n_1171),
.B(n_1145),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1138),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1111),
.B(n_1116),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1068),
.A2(n_1100),
.B(n_1189),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1105),
.A2(n_1072),
.B(n_1140),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1045),
.B(n_1086),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1121),
.A2(n_1083),
.B(n_1110),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1074),
.B(n_1190),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_SL g1277 ( 
.A1(n_1114),
.A2(n_1128),
.B(n_1112),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1156),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1141),
.A2(n_1158),
.A3(n_1164),
.B(n_1092),
.Y(n_1279)
);

NOR2x1_ASAP7_75t_SL g1280 ( 
.A(n_1070),
.B(n_1146),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1107),
.A2(n_1184),
.B(n_1113),
.Y(n_1281)
);

AOI21xp33_ASAP7_75t_L g1282 ( 
.A1(n_1164),
.A2(n_1144),
.B(n_1142),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1188),
.A2(n_1157),
.B(n_1186),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1153),
.B(n_1137),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1172),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1156),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1113),
.A2(n_1128),
.B(n_1114),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_SL g1288 ( 
.A1(n_1186),
.A2(n_1194),
.B(n_1102),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1143),
.A2(n_1132),
.B(n_1194),
.C(n_1191),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1123),
.A2(n_1094),
.B(n_1168),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1123),
.A2(n_1168),
.B(n_1163),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1053),
.B(n_1091),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1126),
.A2(n_1139),
.B(n_1152),
.Y(n_1293)
);

BUFx4_ASAP7_75t_SL g1294 ( 
.A(n_1093),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1159),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_SL g1296 ( 
.A(n_1153),
.B(n_1147),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1060),
.A2(n_1077),
.B(n_1163),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1102),
.A2(n_1130),
.B(n_1120),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1091),
.B(n_1177),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1047),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1119),
.A2(n_1130),
.B(n_1120),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1170),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1167),
.A2(n_1141),
.B1(n_1158),
.B2(n_1134),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1075),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1153),
.B(n_1169),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1183),
.Y(n_1306)
);

NOR4xp25_ASAP7_75t_L g1307 ( 
.A(n_1084),
.B(n_1134),
.C(n_1066),
.D(n_1125),
.Y(n_1307)
);

AND3x1_ASAP7_75t_L g1308 ( 
.A(n_1087),
.B(n_1125),
.C(n_1061),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1066),
.B(n_1096),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1169),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1075),
.A2(n_1103),
.B(n_1131),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1075),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1125),
.A2(n_1103),
.A3(n_1131),
.B(n_1133),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1129),
.B(n_1131),
.Y(n_1314)
);

NOR3xp33_ASAP7_75t_L g1315 ( 
.A(n_1133),
.B(n_1136),
.C(n_1146),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1133),
.Y(n_1316)
);

AOI221xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1136),
.A2(n_1180),
.B1(n_986),
.B2(n_1176),
.C(n_1175),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1136),
.A2(n_986),
.B(n_1048),
.C(n_1098),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1146),
.A2(n_1150),
.B(n_1127),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1193),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1165),
.B(n_986),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1043),
.A2(n_1071),
.A3(n_1069),
.B(n_1065),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1043),
.A2(n_986),
.B(n_865),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1165),
.B(n_986),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1042),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1165),
.B(n_986),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1043),
.A2(n_886),
.B(n_865),
.Y(n_1327)
);

CKINVDCx11_ASAP7_75t_R g1328 ( 
.A(n_1147),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1055),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1048),
.A2(n_986),
.B1(n_865),
.B2(n_864),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1093),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1042),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1043),
.A2(n_1071),
.A3(n_1069),
.B(n_1065),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1150),
.A2(n_1127),
.B(n_1073),
.Y(n_1334)
);

NOR2xp67_ASAP7_75t_SL g1335 ( 
.A(n_1147),
.B(n_831),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1150),
.A2(n_1127),
.B(n_1073),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1043),
.A2(n_1109),
.B(n_1052),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1150),
.A2(n_1127),
.B(n_1073),
.Y(n_1338)
);

O2A1O1Ixp5_ASAP7_75t_L g1339 ( 
.A1(n_1175),
.A2(n_986),
.B(n_996),
.C(n_1176),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_SL g1340 ( 
.A1(n_1180),
.A2(n_1192),
.B(n_1188),
.Y(n_1340)
);

AO32x2_ASAP7_75t_L g1341 ( 
.A1(n_1180),
.A2(n_1057),
.A3(n_1158),
.B1(n_1141),
.B2(n_1134),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_L g1342 ( 
.A(n_1098),
.B(n_831),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1043),
.A2(n_886),
.B(n_865),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1193),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1054),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1048),
.A2(n_986),
.B(n_865),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1042),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1150),
.A2(n_1127),
.B(n_1073),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1043),
.A2(n_886),
.B(n_865),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1234),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1303),
.A2(n_1200),
.B1(n_1308),
.B2(n_1346),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1327),
.A2(n_1349),
.A3(n_1343),
.B(n_1203),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1207),
.B(n_1217),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1348),
.A2(n_1220),
.B(n_1319),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1323),
.A2(n_1197),
.B(n_1240),
.Y(n_1355)
);

AO21x2_ASAP7_75t_L g1356 ( 
.A1(n_1268),
.A2(n_1225),
.B(n_1323),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1232),
.A2(n_1216),
.B(n_1204),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1268),
.A2(n_1225),
.B(n_1215),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1330),
.B(n_1321),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1339),
.A2(n_1282),
.B(n_1200),
.C(n_1289),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1293),
.Y(n_1361)
);

BUFx4f_ASAP7_75t_L g1362 ( 
.A(n_1258),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1318),
.A2(n_1272),
.B(n_1212),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1303),
.A2(n_1308),
.B1(n_1261),
.B2(n_1326),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1269),
.A2(n_1245),
.B(n_1277),
.Y(n_1365)
);

OAI211xp5_ASAP7_75t_L g1366 ( 
.A1(n_1261),
.A2(n_1317),
.B(n_1309),
.C(n_1229),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1281),
.Y(n_1367)
);

NAND2x1p5_ASAP7_75t_L g1368 ( 
.A(n_1233),
.B(n_1329),
.Y(n_1368)
);

NOR2xp67_ASAP7_75t_L g1369 ( 
.A(n_1237),
.B(n_1205),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1324),
.B(n_1263),
.Y(n_1370)
);

OAI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1211),
.A2(n_1208),
.B1(n_1228),
.B2(n_1264),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1292),
.B(n_1196),
.Y(n_1372)
);

OAI221xp5_ASAP7_75t_L g1373 ( 
.A1(n_1211),
.A2(n_1317),
.B1(n_1219),
.B2(n_1198),
.C(n_1224),
.Y(n_1373)
);

AO32x2_ASAP7_75t_L g1374 ( 
.A1(n_1307),
.A2(n_1313),
.A3(n_1341),
.B1(n_1231),
.B2(n_1223),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1316),
.B(n_1242),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1271),
.A2(n_1262),
.B1(n_1342),
.B2(n_1199),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1272),
.A2(n_1340),
.B(n_1290),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1226),
.A2(n_1337),
.B(n_1273),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1345),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1255),
.Y(n_1380)
);

OR2x6_ASAP7_75t_L g1381 ( 
.A(n_1288),
.B(n_1287),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1202),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1267),
.A2(n_1248),
.B1(n_1252),
.B2(n_1284),
.Y(n_1383)
);

CKINVDCx6p67_ASAP7_75t_R g1384 ( 
.A(n_1328),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1276),
.A2(n_1236),
.B1(n_1239),
.B2(n_1285),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1210),
.Y(n_1386)
);

CKINVDCx12_ASAP7_75t_R g1387 ( 
.A(n_1294),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1244),
.A2(n_1249),
.B(n_1250),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1247),
.B(n_1305),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1233),
.B(n_1329),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1285),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1265),
.A2(n_1337),
.B(n_1259),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1260),
.A2(n_1283),
.B(n_1218),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1218),
.A2(n_1275),
.B(n_1297),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1291),
.A2(n_1347),
.B(n_1270),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1300),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1243),
.A2(n_1283),
.B(n_1301),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1299),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1253),
.A2(n_1325),
.B(n_1332),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1243),
.A2(n_1298),
.B(n_1311),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1278),
.B(n_1286),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1274),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1310),
.A2(n_1306),
.B1(n_1302),
.B2(n_1295),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1312),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1221),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1341),
.A2(n_1329),
.B1(n_1233),
.B2(n_1315),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1322),
.A2(n_1333),
.B(n_1213),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1296),
.A2(n_1341),
.B1(n_1279),
.B2(n_1314),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1322),
.A2(n_1333),
.B(n_1213),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1221),
.A2(n_1322),
.B(n_1333),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1210),
.Y(n_1411)
);

NAND2x1p5_ASAP7_75t_L g1412 ( 
.A(n_1335),
.B(n_1246),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1210),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1213),
.A2(n_1209),
.B(n_1206),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1214),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1256),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1214),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1241),
.A2(n_1209),
.B(n_1206),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1296),
.A2(n_1257),
.B1(n_1331),
.B2(n_1256),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1320),
.Y(n_1420)
);

INVx4_ASAP7_75t_L g1421 ( 
.A(n_1320),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1235),
.A2(n_1279),
.B(n_1230),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1344),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1230),
.B(n_1209),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1241),
.A2(n_1206),
.B(n_1230),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1241),
.A2(n_1280),
.B(n_1227),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1222),
.B(n_1227),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1254),
.B(n_1304),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1254),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1304),
.A2(n_1211),
.B1(n_1303),
.B2(n_1261),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1255),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1293),
.Y(n_1432)
);

NAND2x1p5_ASAP7_75t_L g1433 ( 
.A(n_1233),
.B(n_1329),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1321),
.B(n_1324),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1303),
.A2(n_986),
.B1(n_1200),
.B2(n_1308),
.Y(n_1435)
);

AOI222xp33_ASAP7_75t_L g1436 ( 
.A1(n_1211),
.A2(n_1098),
.B1(n_935),
.B2(n_986),
.C1(n_1176),
.C2(n_1175),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1263),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1316),
.B(n_1129),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1334),
.A2(n_1338),
.B(n_1336),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1211),
.A2(n_986),
.B1(n_1098),
.B2(n_1175),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1339),
.A2(n_986),
.B(n_1200),
.Y(n_1441)
);

AOI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1339),
.A2(n_1200),
.B(n_986),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1255),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1316),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1321),
.B(n_1324),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1334),
.A2(n_1338),
.B(n_1336),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1339),
.A2(n_986),
.B(n_1048),
.C(n_1282),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1234),
.Y(n_1448)
);

NAND2x1p5_ASAP7_75t_L g1449 ( 
.A(n_1233),
.B(n_1329),
.Y(n_1449)
);

OAI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1282),
.A2(n_986),
.B1(n_1098),
.B2(n_1339),
.C(n_1200),
.Y(n_1450)
);

NOR2xp67_ASAP7_75t_L g1451 ( 
.A(n_1237),
.B(n_875),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1316),
.B(n_1129),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1303),
.A2(n_986),
.B1(n_1200),
.B2(n_1308),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1346),
.B(n_1330),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1282),
.B(n_399),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1328),
.Y(n_1456)
);

O2A1O1Ixp33_ASAP7_75t_SL g1457 ( 
.A1(n_1289),
.A2(n_986),
.B(n_1282),
.C(n_1200),
.Y(n_1457)
);

BUFx8_ASAP7_75t_L g1458 ( 
.A(n_1331),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_1328),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1200),
.A2(n_986),
.B1(n_1282),
.B2(n_1098),
.Y(n_1460)
);

INVx4_ASAP7_75t_L g1461 ( 
.A(n_1233),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1282),
.B(n_399),
.Y(n_1462)
);

AO31x2_ASAP7_75t_L g1463 ( 
.A1(n_1201),
.A2(n_1238),
.A3(n_1349),
.B(n_1343),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1207),
.B(n_1217),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_SL g1465 ( 
.A(n_1275),
.B(n_1200),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1339),
.A2(n_986),
.B(n_1200),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1233),
.Y(n_1467)
);

AOI222xp33_ASAP7_75t_L g1468 ( 
.A1(n_1211),
.A2(n_1098),
.B1(n_935),
.B2(n_986),
.C1(n_1176),
.C2(n_1175),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1282),
.B(n_399),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1328),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1334),
.A2(n_1338),
.B(n_1336),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1339),
.A2(n_986),
.B(n_1200),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1234),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1210),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1447),
.A2(n_1436),
.B(n_1468),
.C(n_1457),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1399),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1440),
.A2(n_1460),
.B1(n_1435),
.B2(n_1453),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1399),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1359),
.B(n_1454),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1360),
.A2(n_1450),
.B(n_1406),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1391),
.Y(n_1481)
);

NOR2xp67_ASAP7_75t_L g1482 ( 
.A(n_1437),
.B(n_1372),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1393),
.A2(n_1422),
.B(n_1378),
.Y(n_1483)
);

O2A1O1Ixp5_ASAP7_75t_L g1484 ( 
.A1(n_1435),
.A2(n_1453),
.B(n_1351),
.C(n_1441),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1437),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1450),
.A2(n_1406),
.B(n_1390),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1436),
.A2(n_1468),
.B(n_1442),
.C(n_1466),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1430),
.A2(n_1366),
.B1(n_1373),
.B2(n_1351),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1434),
.B(n_1445),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1370),
.B(n_1353),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1398),
.B(n_1364),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1385),
.B(n_1402),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1381),
.B(n_1389),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1393),
.A2(n_1422),
.B(n_1378),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1425),
.A2(n_1418),
.B(n_1397),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1364),
.B(n_1350),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1368),
.A2(n_1449),
.B(n_1390),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1375),
.B(n_1383),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1455),
.B(n_1462),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1459),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1469),
.A2(n_1373),
.B(n_1366),
.C(n_1441),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1371),
.B(n_1466),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1371),
.B(n_1472),
.Y(n_1503)
);

NOR2xp67_ASAP7_75t_L g1504 ( 
.A(n_1382),
.B(n_1380),
.Y(n_1504)
);

O2A1O1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1442),
.A2(n_1472),
.B(n_1430),
.C(n_1363),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1363),
.A2(n_1389),
.B(n_1355),
.C(n_1408),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1424),
.A2(n_1357),
.B(n_1392),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1375),
.B(n_1438),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1376),
.A2(n_1419),
.B1(n_1355),
.B2(n_1389),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1379),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1438),
.B(n_1452),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1444),
.Y(n_1512)
);

O2A1O1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1381),
.A2(n_1356),
.B(n_1448),
.C(n_1473),
.Y(n_1513)
);

CKINVDCx14_ASAP7_75t_R g1514 ( 
.A(n_1384),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1403),
.B(n_1429),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1456),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1404),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1465),
.B(n_1429),
.Y(n_1518)
);

OA22x2_ASAP7_75t_L g1519 ( 
.A1(n_1381),
.A2(n_1415),
.B1(n_1423),
.B2(n_1405),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1431),
.B(n_1369),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1412),
.B(n_1356),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1358),
.A2(n_1362),
.B1(n_1433),
.B2(n_1449),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1412),
.B(n_1420),
.Y(n_1523)
);

O2A1O1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1358),
.A2(n_1377),
.B(n_1401),
.C(n_1416),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1428),
.B(n_1413),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1395),
.B(n_1427),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1368),
.A2(n_1433),
.B(n_1467),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1411),
.B(n_1417),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_SL g1529 ( 
.A1(n_1467),
.A2(n_1461),
.B(n_1443),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1362),
.A2(n_1451),
.B1(n_1432),
.B2(n_1361),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1386),
.B(n_1474),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1407),
.B(n_1409),
.Y(n_1532)
);

A2O1A1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1388),
.A2(n_1410),
.B(n_1365),
.C(n_1367),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1394),
.A2(n_1354),
.B(n_1471),
.Y(n_1534)
);

OR2x6_ASAP7_75t_L g1535 ( 
.A(n_1426),
.B(n_1400),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1396),
.B(n_1470),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1421),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1409),
.B(n_1414),
.Y(n_1538)
);

AOI221x1_ASAP7_75t_SL g1539 ( 
.A1(n_1374),
.A2(n_1387),
.B1(n_1458),
.B2(n_1414),
.C(n_1352),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1374),
.A2(n_1352),
.B1(n_1458),
.B2(n_1463),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1463),
.B(n_1439),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1446),
.B(n_1374),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1434),
.B(n_1445),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1437),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1440),
.A2(n_1303),
.B1(n_986),
.B2(n_1308),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1447),
.A2(n_1339),
.B(n_1282),
.C(n_986),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_L g1547 ( 
.A(n_1440),
.B(n_831),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1467),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1370),
.B(n_1353),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1440),
.A2(n_1303),
.B1(n_986),
.B2(n_1308),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1353),
.B(n_1464),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1456),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1447),
.A2(n_1339),
.B(n_1282),
.C(n_986),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_R g1554 ( 
.A(n_1459),
.B(n_1300),
.Y(n_1554)
);

OA21x2_ASAP7_75t_L g1555 ( 
.A1(n_1393),
.A2(n_1422),
.B(n_1378),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1456),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1353),
.B(n_1464),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1353),
.B(n_1464),
.Y(n_1558)
);

OA22x2_ASAP7_75t_L g1559 ( 
.A1(n_1440),
.A2(n_1303),
.B1(n_1098),
.B2(n_1376),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1389),
.B(n_1438),
.Y(n_1560)
);

NOR2xp67_ASAP7_75t_L g1561 ( 
.A(n_1437),
.B(n_862),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1353),
.B(n_1464),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1434),
.B(n_1445),
.Y(n_1563)
);

OR2x6_ASAP7_75t_L g1564 ( 
.A(n_1381),
.B(n_1389),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1456),
.Y(n_1565)
);

AOI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1457),
.A2(n_1339),
.B1(n_986),
.B2(n_1282),
.C(n_1200),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1362),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1393),
.A2(n_1422),
.B(n_1378),
.Y(n_1568)
);

O2A1O1Ixp5_ASAP7_75t_L g1569 ( 
.A1(n_1435),
.A2(n_1339),
.B(n_986),
.C(n_1200),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1476),
.Y(n_1570)
);

OR2x6_ASAP7_75t_L g1571 ( 
.A(n_1493),
.B(n_1564),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1478),
.Y(n_1572)
);

INVx3_ASAP7_75t_SL g1573 ( 
.A(n_1493),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1519),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1532),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1493),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1538),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1542),
.B(n_1483),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1479),
.B(n_1502),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1483),
.B(n_1494),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1535),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1555),
.B(n_1568),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1495),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1495),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1507),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1559),
.A2(n_1477),
.B1(n_1488),
.B2(n_1550),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1554),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1507),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1526),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1488),
.A2(n_1477),
.B1(n_1550),
.B2(n_1545),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1541),
.Y(n_1591)
);

AO21x1_ASAP7_75t_SL g1592 ( 
.A1(n_1502),
.A2(n_1503),
.B(n_1521),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1534),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1535),
.B(n_1540),
.Y(n_1594)
);

CKINVDCx11_ASAP7_75t_R g1595 ( 
.A(n_1500),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1540),
.B(n_1506),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1517),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1559),
.A2(n_1545),
.B1(n_1499),
.B2(n_1566),
.Y(n_1598)
);

OA21x2_ASAP7_75t_L g1599 ( 
.A1(n_1533),
.A2(n_1484),
.B(n_1569),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1519),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1564),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1480),
.B(n_1479),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1496),
.B(n_1491),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1513),
.Y(n_1604)
);

AOI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1522),
.A2(n_1509),
.B(n_1530),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1539),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1546),
.A2(n_1553),
.B(n_1505),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1524),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1539),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1530),
.Y(n_1610)
);

AO21x2_ASAP7_75t_L g1611 ( 
.A1(n_1509),
.A2(n_1501),
.B(n_1487),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1475),
.B(n_1492),
.Y(n_1612)
);

AO21x2_ASAP7_75t_L g1613 ( 
.A1(n_1518),
.A2(n_1486),
.B(n_1522),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1485),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1544),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1498),
.A2(n_1515),
.B(n_1528),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1560),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1560),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1481),
.Y(n_1619)
);

OAI211xp5_ASAP7_75t_L g1620 ( 
.A1(n_1586),
.A2(n_1482),
.B(n_1481),
.C(n_1561),
.Y(n_1620)
);

NOR2x1_ASAP7_75t_SL g1621 ( 
.A(n_1592),
.B(n_1571),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1578),
.B(n_1557),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1591),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1572),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1570),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1570),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1578),
.B(n_1551),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1578),
.B(n_1562),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1590),
.A2(n_1508),
.B(n_1514),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1579),
.B(n_1489),
.Y(n_1630)
);

INVx4_ASAP7_75t_L g1631 ( 
.A(n_1571),
.Y(n_1631)
);

INVx4_ASAP7_75t_L g1632 ( 
.A(n_1571),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1580),
.B(n_1558),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1579),
.B(n_1543),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1580),
.B(n_1510),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1582),
.B(n_1510),
.Y(n_1636)
);

NOR2x1_ASAP7_75t_L g1637 ( 
.A(n_1613),
.B(n_1497),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1582),
.B(n_1490),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1591),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1612),
.B(n_1563),
.Y(n_1640)
);

AOI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1586),
.A2(n_1547),
.B1(n_1549),
.B2(n_1512),
.C(n_1520),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1575),
.B(n_1523),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1589),
.B(n_1531),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1582),
.B(n_1511),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1575),
.B(n_1537),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1593),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1593),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1589),
.B(n_1525),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1593),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1590),
.B(n_1504),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1581),
.B(n_1548),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1575),
.B(n_1529),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1577),
.B(n_1567),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1638),
.B(n_1589),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1650),
.A2(n_1611),
.B1(n_1598),
.B2(n_1612),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1622),
.B(n_1618),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1638),
.B(n_1615),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_L g1658 ( 
.A1(n_1629),
.A2(n_1598),
.B1(n_1602),
.B2(n_1600),
.C(n_1574),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_SL g1659 ( 
.A(n_1623),
.B(n_1592),
.Y(n_1659)
);

AO21x2_ASAP7_75t_L g1660 ( 
.A1(n_1621),
.A2(n_1585),
.B(n_1588),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1650),
.A2(n_1607),
.B(n_1611),
.Y(n_1661)
);

NAND2xp33_ASAP7_75t_R g1662 ( 
.A(n_1640),
.B(n_1587),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1640),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1620),
.A2(n_1602),
.B(n_1596),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1641),
.A2(n_1602),
.B1(n_1596),
.B2(n_1611),
.C(n_1609),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1641),
.A2(n_1596),
.B1(n_1611),
.B2(n_1606),
.C(n_1609),
.Y(n_1666)
);

OR2x6_ASAP7_75t_L g1667 ( 
.A(n_1637),
.B(n_1571),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1630),
.A2(n_1611),
.B1(n_1606),
.B2(n_1608),
.C(n_1604),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1631),
.A2(n_1607),
.B1(n_1571),
.B2(n_1576),
.Y(n_1669)
);

AO21x2_ASAP7_75t_L g1670 ( 
.A1(n_1621),
.A2(n_1588),
.B(n_1585),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1620),
.A2(n_1600),
.B1(n_1574),
.B2(n_1604),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1637),
.B(n_1608),
.C(n_1604),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1625),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1629),
.A2(n_1610),
.B1(n_1605),
.B2(n_1608),
.C(n_1599),
.Y(n_1674)
);

AOI222xp33_ASAP7_75t_L g1675 ( 
.A1(n_1630),
.A2(n_1595),
.B1(n_1610),
.B2(n_1587),
.C1(n_1603),
.C2(n_1614),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1634),
.A2(n_1574),
.B1(n_1600),
.B2(n_1599),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1634),
.B(n_1595),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1625),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1642),
.A2(n_1597),
.B1(n_1614),
.B2(n_1619),
.C(n_1607),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1635),
.B(n_1615),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1622),
.B(n_1618),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1652),
.A2(n_1605),
.B1(n_1599),
.B2(n_1573),
.C(n_1571),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_L g1683 ( 
.A(n_1652),
.B(n_1613),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1626),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1624),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1648),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1626),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1633),
.B(n_1616),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1633),
.B(n_1616),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1631),
.A2(n_1607),
.B1(n_1571),
.B2(n_1573),
.Y(n_1690)
);

AOI31xp33_ASAP7_75t_L g1691 ( 
.A1(n_1623),
.A2(n_1619),
.A3(n_1617),
.B(n_1594),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1651),
.B(n_1576),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1631),
.A2(n_1573),
.B1(n_1601),
.B2(n_1576),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1653),
.Y(n_1694)
);

AO21x2_ASAP7_75t_L g1695 ( 
.A1(n_1646),
.A2(n_1588),
.B(n_1585),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_SL g1696 ( 
.A(n_1623),
.B(n_1592),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1648),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1660),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1663),
.B(n_1679),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1660),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1673),
.Y(n_1701)
);

OR2x6_ASAP7_75t_L g1702 ( 
.A(n_1661),
.B(n_1631),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1695),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1685),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1678),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1659),
.B(n_1633),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1676),
.A2(n_1583),
.B(n_1584),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1695),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1670),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_1677),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1684),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1670),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1687),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1655),
.B(n_1653),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1692),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1657),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1680),
.Y(n_1717)
);

AOI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1676),
.A2(n_1649),
.B(n_1647),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1688),
.B(n_1639),
.Y(n_1719)
);

INVx4_ASAP7_75t_SL g1720 ( 
.A(n_1667),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1680),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1689),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1654),
.Y(n_1723)
);

INVx4_ASAP7_75t_SL g1724 ( 
.A(n_1667),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1654),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1667),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1697),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1686),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1696),
.B(n_1627),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1694),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1656),
.B(n_1627),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_L g1732 ( 
.A(n_1699),
.B(n_1672),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1698),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1714),
.A2(n_1665),
.B1(n_1666),
.B2(n_1607),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1701),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1723),
.B(n_1725),
.Y(n_1736)
);

AOI222xp33_ASAP7_75t_L g1737 ( 
.A1(n_1699),
.A2(n_1668),
.B1(n_1674),
.B2(n_1658),
.C1(n_1664),
.C2(n_1671),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1720),
.B(n_1683),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1698),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1723),
.B(n_1643),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1704),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1725),
.B(n_1645),
.Y(n_1742)
);

INVx4_ASAP7_75t_L g1743 ( 
.A(n_1720),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1730),
.B(n_1675),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1729),
.B(n_1692),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1729),
.B(n_1681),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1701),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1698),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1720),
.B(n_1631),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1706),
.B(n_1627),
.Y(n_1750)
);

CKINVDCx20_ASAP7_75t_R g1751 ( 
.A(n_1710),
.Y(n_1751)
);

AND3x2_ASAP7_75t_L g1752 ( 
.A(n_1726),
.B(n_1704),
.C(n_1730),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1726),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1706),
.B(n_1628),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1705),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_L g1756 ( 
.A(n_1730),
.B(n_1691),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1705),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1720),
.B(n_1628),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1720),
.B(n_1628),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1724),
.B(n_1632),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1724),
.B(n_1690),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1715),
.A2(n_1674),
.B1(n_1632),
.B2(n_1675),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1724),
.B(n_1635),
.Y(n_1763)
);

NOR2x1_ASAP7_75t_L g1764 ( 
.A(n_1728),
.B(n_1664),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1711),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1724),
.B(n_1636),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1724),
.B(n_1636),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1716),
.B(n_1644),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1711),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1713),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1727),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1744),
.B(n_1728),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1745),
.B(n_1715),
.Y(n_1773)
);

INVx2_ASAP7_75t_SL g1774 ( 
.A(n_1752),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_SL g1775 ( 
.A(n_1764),
.B(n_1671),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1755),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1735),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1732),
.B(n_1717),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1735),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1741),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1753),
.B(n_1768),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1745),
.B(n_1715),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1746),
.B(n_1758),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1747),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1747),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1757),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1737),
.A2(n_1662),
.B1(n_1682),
.B2(n_1669),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1732),
.B(n_1728),
.Y(n_1788)
);

AND2x2_ASAP7_75t_SL g1789 ( 
.A(n_1734),
.B(n_1632),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1751),
.B(n_1516),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1757),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1753),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1743),
.B(n_1552),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1743),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1743),
.B(n_1707),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1765),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_SL g1797 ( 
.A(n_1756),
.B(n_1682),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1736),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1758),
.B(n_1719),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1738),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1765),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1742),
.B(n_1721),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1746),
.B(n_1731),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1769),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1769),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1742),
.B(n_1721),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1771),
.B(n_1713),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1770),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1777),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1779),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1783),
.B(n_1761),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1792),
.B(n_1750),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1788),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1787),
.A2(n_1762),
.B1(n_1761),
.B2(n_1760),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1784),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1799),
.Y(n_1816)
);

CKINVDCx16_ASAP7_75t_R g1817 ( 
.A(n_1775),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1792),
.B(n_1750),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1785),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1774),
.B(n_1759),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1772),
.B(n_1736),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1786),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1778),
.B(n_1770),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1800),
.Y(n_1824)
);

INVxp33_ASAP7_75t_L g1825 ( 
.A(n_1793),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1791),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1773),
.B(n_1782),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1800),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1795),
.A2(n_1739),
.B(n_1733),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1799),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1778),
.B(n_1740),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1803),
.B(n_1759),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1794),
.B(n_1738),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1780),
.B(n_1740),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1814),
.A2(n_1797),
.B1(n_1775),
.B2(n_1789),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1820),
.B(n_1827),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1809),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1809),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1820),
.Y(n_1839)
);

INVxp67_ASAP7_75t_SL g1840 ( 
.A(n_1813),
.Y(n_1840)
);

AOI222xp33_ASAP7_75t_L g1841 ( 
.A1(n_1813),
.A2(n_1797),
.B1(n_1776),
.B2(n_1798),
.C1(n_1738),
.C2(n_1805),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1824),
.B(n_1781),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1817),
.A2(n_1702),
.B1(n_1805),
.B2(n_1807),
.Y(n_1843)
);

INVxp67_ASAP7_75t_SL g1844 ( 
.A(n_1816),
.Y(n_1844)
);

INVxp67_ASAP7_75t_SL g1845 ( 
.A(n_1816),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1812),
.B(n_1807),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1816),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1817),
.A2(n_1749),
.B1(n_1760),
.B2(n_1767),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1828),
.B(n_1796),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1810),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1811),
.A2(n_1749),
.B1(n_1760),
.B2(n_1763),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1827),
.B(n_1754),
.Y(n_1852)
);

INVx2_ASAP7_75t_SL g1853 ( 
.A(n_1830),
.Y(n_1853)
);

OAI21xp33_ASAP7_75t_SL g1854 ( 
.A1(n_1829),
.A2(n_1804),
.B(n_1801),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1836),
.B(n_1830),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1839),
.B(n_1818),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1842),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1847),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_R g1859 ( 
.A(n_1853),
.B(n_1556),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1852),
.B(n_1811),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1847),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1844),
.B(n_1832),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1840),
.B(n_1825),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1845),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1853),
.B(n_1832),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1841),
.B(n_1852),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1848),
.B(n_1833),
.Y(n_1867)
);

NOR3xp33_ASAP7_75t_L g1868 ( 
.A(n_1863),
.B(n_1849),
.C(n_1846),
.Y(n_1868)
);

NAND4xp25_ASAP7_75t_L g1869 ( 
.A(n_1866),
.B(n_1835),
.C(n_1843),
.D(n_1851),
.Y(n_1869)
);

OAI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1857),
.A2(n_1834),
.B1(n_1702),
.B2(n_1821),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1863),
.A2(n_1835),
.B(n_1854),
.Y(n_1871)
);

NAND4xp25_ASAP7_75t_L g1872 ( 
.A(n_1856),
.B(n_1843),
.C(n_1837),
.D(n_1838),
.Y(n_1872)
);

NOR3x1_ASAP7_75t_L g1873 ( 
.A(n_1862),
.B(n_1850),
.C(n_1815),
.Y(n_1873)
);

AOI222xp33_ASAP7_75t_L g1874 ( 
.A1(n_1864),
.A2(n_1826),
.B1(n_1810),
.B2(n_1822),
.C1(n_1815),
.C2(n_1819),
.Y(n_1874)
);

NOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1861),
.B(n_1819),
.Y(n_1875)
);

NAND2xp33_ASAP7_75t_SL g1876 ( 
.A(n_1859),
.B(n_1821),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1865),
.A2(n_1826),
.B1(n_1822),
.B2(n_1833),
.C(n_1834),
.Y(n_1877)
);

AOI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1867),
.A2(n_1823),
.B(n_1829),
.C(n_1831),
.Y(n_1878)
);

OAI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1871),
.A2(n_1855),
.B1(n_1858),
.B2(n_1860),
.C(n_1861),
.Y(n_1879)
);

OAI211xp5_ASAP7_75t_SL g1880 ( 
.A1(n_1878),
.A2(n_1868),
.B(n_1877),
.C(n_1874),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1876),
.A2(n_1749),
.B1(n_1808),
.B2(n_1831),
.Y(n_1881)
);

NOR4xp25_ASAP7_75t_L g1882 ( 
.A(n_1869),
.B(n_1823),
.C(n_1859),
.D(n_1733),
.Y(n_1882)
);

AND4x1_ASAP7_75t_L g1883 ( 
.A(n_1873),
.B(n_1790),
.C(n_1536),
.D(n_1763),
.Y(n_1883)
);

OAI321xp33_ASAP7_75t_L g1884 ( 
.A1(n_1872),
.A2(n_1795),
.A3(n_1702),
.B1(n_1718),
.B2(n_1693),
.C(n_1748),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1875),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1883),
.B(n_1754),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1885),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1882),
.B(n_1766),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1879),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1881),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1880),
.Y(n_1891)
);

NOR2x1_ASAP7_75t_L g1892 ( 
.A(n_1884),
.B(n_1870),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1887),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1888),
.Y(n_1894)
);

AOI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1891),
.A2(n_1702),
.B1(n_1767),
.B2(n_1766),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1891),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1886),
.B(n_1565),
.Y(n_1897)
);

NAND2xp33_ASAP7_75t_R g1898 ( 
.A(n_1890),
.B(n_1806),
.Y(n_1898)
);

NAND4xp75_ASAP7_75t_L g1899 ( 
.A(n_1897),
.B(n_1889),
.C(n_1892),
.D(n_1748),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_SL g1900 ( 
.A1(n_1898),
.A2(n_1895),
.B(n_1894),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1893),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1900),
.Y(n_1902)
);

AOI32xp33_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1901),
.A3(n_1896),
.B1(n_1899),
.B2(n_1893),
.Y(n_1903)
);

NAND4xp25_ASAP7_75t_L g1904 ( 
.A(n_1903),
.B(n_1739),
.C(n_1802),
.D(n_1527),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1903),
.Y(n_1905)
);

XNOR2xp5_ASAP7_75t_L g1906 ( 
.A(n_1905),
.B(n_1702),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1904),
.A2(n_1700),
.B(n_1712),
.Y(n_1907)
);

XNOR2xp5_ASAP7_75t_L g1908 ( 
.A(n_1906),
.B(n_1702),
.Y(n_1908)
);

AO21x1_ASAP7_75t_L g1909 ( 
.A1(n_1907),
.A2(n_1709),
.B(n_1712),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1908),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1910),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1911),
.B(n_1909),
.Y(n_1912)
);

OAI221xp5_ASAP7_75t_R g1913 ( 
.A1(n_1912),
.A2(n_1700),
.B1(n_1709),
.B2(n_1712),
.C(n_1718),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1913),
.A2(n_1700),
.B1(n_1709),
.B2(n_1722),
.Y(n_1914)
);

AOI211xp5_ASAP7_75t_L g1915 ( 
.A1(n_1914),
.A2(n_1707),
.B(n_1708),
.C(n_1703),
.Y(n_1915)
);


endmodule