module fake_aes_12756_n_524 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_524);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_524;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_388;
wire n_139;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g63 ( .A(n_11), .Y(n_63) );
INVx1_ASAP7_75t_L g64 ( .A(n_57), .Y(n_64) );
INVxp67_ASAP7_75t_SL g65 ( .A(n_42), .Y(n_65) );
INVx2_ASAP7_75t_L g66 ( .A(n_31), .Y(n_66) );
CKINVDCx20_ASAP7_75t_R g67 ( .A(n_48), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_27), .Y(n_68) );
INVxp67_ASAP7_75t_L g69 ( .A(n_36), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_11), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_16), .Y(n_71) );
CKINVDCx5p33_ASAP7_75t_R g72 ( .A(n_38), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_39), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_46), .Y(n_74) );
CKINVDCx14_ASAP7_75t_R g75 ( .A(n_45), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_1), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_50), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_22), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_58), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_28), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_51), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_54), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_52), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_30), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_24), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_40), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_5), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_56), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_3), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_4), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_2), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_20), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_35), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_29), .Y(n_95) );
INVxp33_ASAP7_75t_L g96 ( .A(n_12), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_43), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_4), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_10), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_8), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_32), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_41), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_7), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_66), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_64), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_66), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_102), .B(n_0), .Y(n_107) );
NOR2xp33_ASAP7_75t_R g108 ( .A(n_75), .B(n_18), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_63), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_63), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_64), .Y(n_111) );
INVx4_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_67), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_71), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_96), .B(n_0), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_101), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_83), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_101), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_71), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_92), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_73), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_73), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_74), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_74), .B(n_1), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_68), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_77), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_79), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_78), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_85), .B(n_2), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_70), .B(n_3), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_70), .B(n_5), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_93), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_94), .B(n_6), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_97), .Y(n_136) );
BUFx2_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_116), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_109), .Y(n_140) );
INVx2_ASAP7_75t_SL g141 ( .A(n_112), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_112), .B(n_89), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
BUFx4f_ASAP7_75t_L g145 ( .A(n_105), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_137), .B(n_100), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_137), .B(n_76), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_132), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_112), .B(n_76), .Y(n_149) );
BUFx4f_ASAP7_75t_L g150 ( .A(n_105), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_132), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
BUFx4f_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
NOR2xp33_ASAP7_75t_SL g154 ( .A(n_112), .B(n_95), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_110), .Y(n_155) );
AO22x2_ASAP7_75t_L g156 ( .A1(n_129), .A2(n_114), .B1(n_119), .B2(n_134), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_119), .B(n_100), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_133), .B(n_80), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_133), .B(n_80), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_111), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_116), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_111), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_129), .B(n_72), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_111), .B(n_103), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_111), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_116), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_116), .Y(n_167) );
INVxp67_ASAP7_75t_L g168 ( .A(n_127), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_134), .B(n_95), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_121), .A2(n_98), .B1(n_91), .B2(n_90), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_122), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_122), .Y(n_172) );
NAND3xp33_ASAP7_75t_L g173 ( .A(n_107), .B(n_87), .C(n_82), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_125), .B(n_69), .Y(n_174) );
INVxp33_ASAP7_75t_L g175 ( .A(n_115), .Y(n_175) );
INVx4_ASAP7_75t_SL g176 ( .A(n_130), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_126), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_155), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_160), .Y(n_180) );
INVx5_ASAP7_75t_L g181 ( .A(n_171), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_143), .B(n_125), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_142), .B(n_135), .Y(n_184) );
BUFx12f_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_155), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_163), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_146), .B(n_175), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_156), .A2(n_117), .B1(n_113), .B2(n_120), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_176), .Y(n_191) );
NOR2xp33_ASAP7_75t_R g192 ( .A(n_140), .B(n_82), .Y(n_192) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_145), .B(n_124), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_144), .A2(n_123), .B(n_136), .C(n_99), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_156), .A2(n_121), .B1(n_123), .B2(n_136), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_146), .B(n_121), .Y(n_196) );
CKINVDCx12_ASAP7_75t_R g197 ( .A(n_147), .Y(n_197) );
INVxp67_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_168), .Y(n_199) );
INVx5_ASAP7_75t_L g200 ( .A(n_171), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_159), .B(n_169), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_149), .B(n_130), .Y(n_202) );
BUFx12f_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_149), .B(n_130), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_148), .B(n_136), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_151), .B(n_106), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_164), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
CKINVDCx6p67_ASAP7_75t_R g210 ( .A(n_147), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_164), .Y(n_211) );
NOR2xp33_ASAP7_75t_R g212 ( .A(n_154), .B(n_6), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_157), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_145), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_145), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_173), .B(n_106), .Y(n_220) );
NOR3xp33_ASAP7_75t_SL g221 ( .A(n_174), .B(n_65), .C(n_81), .Y(n_221) );
INVx5_ASAP7_75t_L g222 ( .A(n_171), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_182), .A2(n_150), .B1(n_153), .B2(n_174), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_203), .Y(n_224) );
INVxp67_ASAP7_75t_L g225 ( .A(n_189), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_180), .Y(n_226) );
INVx3_ASAP7_75t_SL g227 ( .A(n_210), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_191), .B(n_153), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_180), .Y(n_229) );
OR2x2_ASAP7_75t_L g230 ( .A(n_187), .B(n_170), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g231 ( .A1(n_185), .A2(n_99), .B1(n_141), .B2(n_104), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_201), .A2(n_202), .B(n_204), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_209), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_203), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_185), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_198), .B(n_196), .Y(n_236) );
INVx5_ASAP7_75t_L g237 ( .A(n_191), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g238 ( .A1(n_199), .A2(n_141), .B1(n_104), .B2(n_106), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_188), .B(n_176), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_191), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_209), .Y(n_241) );
INVx5_ASAP7_75t_L g242 ( .A(n_218), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_213), .B(n_176), .Y(n_243) );
BUFx2_ASAP7_75t_L g244 ( .A(n_212), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_197), .B(n_176), .Y(n_245) );
INVx8_ASAP7_75t_L g246 ( .A(n_205), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g247 ( .A1(n_216), .A2(n_84), .B(n_172), .C(n_161), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_215), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_215), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_218), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_184), .B(n_104), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_195), .B(n_118), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_184), .B(n_108), .Y(n_253) );
NOR2x1_ASAP7_75t_SL g254 ( .A(n_214), .B(n_126), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_212), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_179), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_207), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_227), .B(n_179), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_252), .A2(n_184), .B1(n_195), .B2(n_220), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_246), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_227), .B(n_190), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_227), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
OAI22xp5_ASAP7_75t_SL g264 ( .A1(n_256), .A2(n_186), .B1(n_199), .B2(n_192), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_246), .Y(n_265) );
NOR2x1p5_ASAP7_75t_L g266 ( .A(n_230), .B(n_186), .Y(n_266) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_229), .A2(n_166), .B(n_161), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_236), .Y(n_268) );
INVx4_ASAP7_75t_L g269 ( .A(n_246), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_SL g270 ( .A1(n_223), .A2(n_183), .B(n_194), .C(n_219), .Y(n_270) );
AOI221xp5_ASAP7_75t_L g271 ( .A1(n_225), .A2(n_221), .B1(n_205), .B2(n_192), .C(n_206), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_236), .B(n_205), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_238), .A2(n_211), .B1(n_208), .B2(n_183), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_232), .A2(n_220), .B(n_206), .C(n_118), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_230), .B(n_206), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_235), .B(n_193), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_229), .A2(n_217), .B1(n_220), .B2(n_193), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_234), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_252), .A2(n_128), .B1(n_126), .B2(n_122), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_251), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_251), .Y(n_281) );
OA21x2_ASAP7_75t_L g282 ( .A1(n_274), .A2(n_233), .B(n_249), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_272), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_267), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_261), .A2(n_246), .B1(n_244), .B2(n_255), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_268), .B(n_235), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_267), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_271), .A2(n_231), .B1(n_251), .B2(n_253), .C(n_224), .Y(n_288) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_267), .A2(n_248), .B(n_241), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_260), .Y(n_290) );
CKINVDCx14_ASAP7_75t_R g291 ( .A(n_264), .Y(n_291) );
AOI222xp33_ASAP7_75t_L g292 ( .A1(n_266), .A2(n_244), .B1(n_224), .B2(n_257), .C1(n_233), .C2(n_249), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_274), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_260), .Y(n_294) );
AOI22xp33_ASAP7_75t_SL g295 ( .A1(n_265), .A2(n_254), .B1(n_248), .B2(n_226), .Y(n_295) );
OAI21x1_ASAP7_75t_SL g296 ( .A1(n_277), .A2(n_254), .B(n_241), .Y(n_296) );
AOI22xp33_ASAP7_75t_SL g297 ( .A1(n_269), .A2(n_239), .B1(n_245), .B2(n_237), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_259), .B(n_239), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_263), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_275), .A2(n_250), .B1(n_242), .B2(n_243), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_259), .A2(n_250), .B1(n_242), .B2(n_240), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_298), .B(n_281), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_284), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_284), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_288), .A2(n_273), .B(n_270), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_298), .B(n_280), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_291), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_288), .A2(n_278), .B1(n_270), .B2(n_279), .C(n_258), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_284), .Y(n_309) );
OAI211xp5_ASAP7_75t_L g310 ( .A1(n_292), .A2(n_276), .B(n_279), .C(n_262), .Y(n_310) );
NOR2xp33_ASAP7_75t_R g311 ( .A(n_290), .B(n_237), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_294), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_299), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_299), .Y(n_315) );
AOI21x1_ASAP7_75t_L g316 ( .A1(n_287), .A2(n_118), .B(n_166), .Y(n_316) );
AND4x1_ASAP7_75t_L g317 ( .A(n_292), .B(n_7), .C(n_8), .D(n_9), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_286), .A2(n_247), .B1(n_122), .B2(n_126), .C(n_128), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_287), .Y(n_319) );
AO221x2_ASAP7_75t_L g320 ( .A1(n_285), .A2(n_9), .B1(n_10), .B2(n_12), .C(n_13), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_290), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_296), .B(n_228), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_283), .A2(n_242), .B1(n_250), .B2(n_126), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_289), .Y(n_325) );
NAND4xp25_ASAP7_75t_L g326 ( .A(n_293), .B(n_178), .C(n_177), .D(n_13), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_283), .B(n_122), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_290), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_289), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_302), .B(n_293), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_302), .B(n_282), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_322), .B(n_289), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_306), .B(n_282), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_303), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_306), .B(n_282), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_319), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_319), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_311), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_313), .B(n_282), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_322), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_313), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_312), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_315), .B(n_295), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_315), .B(n_295), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_312), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_304), .B(n_301), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_304), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_309), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_322), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_322), .B(n_300), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_323), .B(n_122), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_328), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_323), .B(n_128), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_322), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_314), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_314), .B(n_297), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_329), .B(n_128), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_325), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_305), .B(n_297), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_321), .B(n_128), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_316), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_321), .Y(n_365) );
AND2x4_ASAP7_75t_SL g366 ( .A(n_324), .B(n_240), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_316), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_327), .B(n_14), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_330), .B(n_320), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_330), .B(n_320), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_338), .B(n_317), .Y(n_372) );
NOR4xp25_ASAP7_75t_SL g373 ( .A(n_338), .B(n_307), .C(n_308), .D(n_320), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_345), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_367), .A2(n_317), .B(n_310), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_342), .B(n_320), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_353), .B(n_327), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_353), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_369), .B(n_237), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_341), .B(n_307), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_341), .B(n_318), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_331), .B(n_250), .Y(n_382) );
INVxp33_ASAP7_75t_SL g383 ( .A(n_365), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_332), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_331), .B(n_15), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_355), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_363), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_336), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_369), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_369), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_335), .B(n_17), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_340), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_356), .B(n_237), .Y(n_393) );
AOI211xp5_ASAP7_75t_SL g394 ( .A1(n_356), .A2(n_240), .B(n_21), .C(n_23), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_355), .B(n_19), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_337), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_337), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_369), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_335), .B(n_138), .Y(n_399) );
NOR3xp33_ASAP7_75t_L g400 ( .A(n_361), .B(n_172), .C(n_178), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_334), .B(n_25), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_354), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_334), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_361), .A2(n_228), .B(n_242), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_339), .B(n_333), .Y(n_405) );
INVx4_ASAP7_75t_L g406 ( .A(n_363), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_354), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_334), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_343), .B(n_26), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_346), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_356), .B(n_33), .Y(n_411) );
NOR3xp33_ASAP7_75t_SL g412 ( .A(n_358), .B(n_34), .C(n_37), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_346), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_364), .A2(n_237), .B(n_228), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_343), .B(n_47), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_346), .Y(n_416) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_359), .B(n_172), .C(n_177), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_383), .B(n_344), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_396), .Y(n_419) );
NOR4xp25_ASAP7_75t_L g420 ( .A(n_375), .B(n_358), .C(n_344), .D(n_356), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_372), .A2(n_351), .B1(n_340), .B2(n_350), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_378), .B(n_351), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_397), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_375), .A2(n_359), .B(n_339), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_386), .Y(n_427) );
INVxp33_ASAP7_75t_L g428 ( .A(n_380), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_370), .A2(n_351), .B1(n_350), .B2(n_332), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_376), .A2(n_351), .B(n_347), .Y(n_430) );
OAI32xp33_ASAP7_75t_L g431 ( .A1(n_379), .A2(n_347), .A3(n_364), .B1(n_357), .B2(n_348), .Y(n_431) );
NOR2xp67_ASAP7_75t_L g432 ( .A(n_384), .B(n_364), .Y(n_432) );
NAND4xp25_ASAP7_75t_L g433 ( .A(n_370), .B(n_332), .C(n_352), .D(n_360), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_408), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_374), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_402), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_389), .A2(n_366), .B1(n_348), .B2(n_357), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_407), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
AOI322xp5_ASAP7_75t_L g440 ( .A1(n_371), .A2(n_348), .A3(n_349), .B1(n_357), .B2(n_362), .C1(n_364), .C2(n_368), .Y(n_440) );
AO22x1_ASAP7_75t_L g441 ( .A1(n_392), .A2(n_349), .B1(n_368), .B2(n_362), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_405), .B(n_349), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_394), .A2(n_368), .B(n_366), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_410), .Y(n_444) );
OAI32xp33_ASAP7_75t_L g445 ( .A1(n_406), .A2(n_49), .A3(n_53), .B1(n_55), .B2(n_59), .Y(n_445) );
INVxp33_ASAP7_75t_L g446 ( .A(n_385), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_394), .A2(n_152), .B(n_167), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_390), .A2(n_222), .B1(n_200), .B2(n_181), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_406), .B(n_60), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_414), .A2(n_222), .B(n_200), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_398), .A2(n_400), .B1(n_415), .B2(n_409), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_416), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_413), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_399), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_405), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_417), .A2(n_152), .B1(n_167), .B2(n_138), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_382), .A2(n_167), .B1(n_138), .B2(n_139), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_455), .B(n_387), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_423), .Y(n_459) );
NOR3xp33_ASAP7_75t_SL g460 ( .A(n_447), .B(n_404), .C(n_411), .Y(n_460) );
XNOR2xp5_ASAP7_75t_L g461 ( .A(n_435), .B(n_391), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_426), .B(n_387), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_428), .B(n_381), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_423), .B(n_399), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_436), .B(n_373), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_438), .B(n_404), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_422), .B(n_393), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_419), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_424), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_427), .Y(n_470) );
OAI221xp5_ASAP7_75t_SL g471 ( .A1(n_420), .A2(n_395), .B1(n_401), .B2(n_412), .C(n_393), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_442), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_418), .B(n_61), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_434), .Y(n_474) );
NOR2xp33_ASAP7_75t_SL g475 ( .A(n_433), .B(n_167), .Y(n_475) );
OAI21xp33_ASAP7_75t_L g476 ( .A1(n_425), .A2(n_138), .B(n_139), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_454), .B(n_139), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_444), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_453), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_454), .B(n_139), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_446), .B(n_62), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g482 ( .A(n_449), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_439), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_452), .Y(n_484) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_429), .A2(n_152), .B(n_171), .Y(n_485) );
XOR2xp5_ASAP7_75t_L g486 ( .A(n_461), .B(n_421), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_475), .B(n_432), .Y(n_487) );
AOI31xp33_ASAP7_75t_L g488 ( .A1(n_465), .A2(n_430), .A3(n_451), .B(n_443), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_459), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_462), .B(n_437), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_482), .B(n_443), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_460), .B(n_440), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_474), .B(n_441), .Y(n_493) );
XOR2x2_ASAP7_75t_L g494 ( .A(n_463), .B(n_448), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_472), .B(n_431), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_478), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_479), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_458), .Y(n_498) );
OAI22xp33_ASAP7_75t_SL g499 ( .A1(n_471), .A2(n_457), .B1(n_450), .B2(n_445), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_464), .B(n_456), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_464), .Y(n_501) );
NAND2xp33_ASAP7_75t_SL g502 ( .A(n_491), .B(n_460), .Y(n_502) );
NOR2xp33_ASAP7_75t_R g503 ( .A(n_489), .B(n_481), .Y(n_503) );
OAI21xp33_ASAP7_75t_L g504 ( .A1(n_492), .A2(n_466), .B(n_485), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_501), .B(n_470), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_492), .B(n_468), .Y(n_506) );
NOR2xp33_ASAP7_75t_R g507 ( .A(n_500), .B(n_481), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_491), .A2(n_473), .B(n_476), .C(n_469), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_488), .A2(n_473), .B1(n_484), .B2(n_483), .C(n_467), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_499), .A2(n_477), .B(n_480), .C(n_450), .Y(n_510) );
XNOR2x1_ASAP7_75t_L g511 ( .A(n_494), .B(n_222), .Y(n_511) );
XNOR2xp5_ASAP7_75t_L g512 ( .A(n_486), .B(n_181), .Y(n_512) );
NAND4xp25_ASAP7_75t_SL g513 ( .A(n_493), .B(n_200), .C(n_495), .D(n_494), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_487), .A2(n_490), .B(n_498), .C(n_496), .Y(n_514) );
NAND5xp2_ASAP7_75t_L g515 ( .A(n_497), .B(n_375), .C(n_475), .D(n_460), .E(n_447), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_502), .A2(n_509), .B1(n_504), .B2(n_513), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_506), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_505), .Y(n_518) );
INVxp67_ASAP7_75t_L g519 ( .A(n_517), .Y(n_519) );
AOI211xp5_ASAP7_75t_L g520 ( .A1(n_516), .A2(n_515), .B(n_514), .C(n_510), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_519), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_521), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_522), .A2(n_520), .B1(n_511), .B2(n_518), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g524 ( .A1(n_523), .A2(n_503), .B1(n_508), .B2(n_507), .C(n_512), .Y(n_524) );
endmodule