module fake_jpeg_28989_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_52),
.Y(n_55)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_0),
.CON(n_47),
.SN(n_47)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_42),
.B1(n_36),
.B2(n_6),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_2),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_5),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_38),
.B1(n_45),
.B2(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_67),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_82),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_36),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_15),
.C(n_16),
.Y(n_91)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_81),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_5),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_31),
.Y(n_86)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_8),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_56),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_86),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_91),
.B(n_78),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_17),
.B(n_18),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_99),
.A2(n_100),
.B1(n_92),
.B2(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_72),
.C(n_73),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_71),
.B1(n_86),
.B2(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_68),
.B1(n_97),
.B2(n_84),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_104),
.A2(n_105),
.B(n_103),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_102),
.C(n_21),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_30),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_20),
.C(n_22),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_26),
.Y(n_110)
);


endmodule