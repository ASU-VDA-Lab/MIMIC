module fake_jpeg_31457_n_232 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_165;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_11),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_49),
.Y(n_64)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_57),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_15),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_1),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_36),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_28),
.B1(n_37),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_77),
.B1(n_81),
.B2(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_61),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_36),
.B1(n_38),
.B2(n_29),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_27),
.B1(n_37),
.B2(n_35),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_79),
.B1(n_86),
.B2(n_90),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_83),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_30),
.B1(n_17),
.B2(n_35),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_36),
.B1(n_20),
.B2(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_34),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_33),
.B1(n_32),
.B2(n_22),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_33),
.B1(n_22),
.B2(n_19),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_19),
.B1(n_26),
.B2(n_4),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_65),
.B(n_12),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_98),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_106),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_26),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_26),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_69),
.A2(n_44),
.B1(n_52),
.B2(n_58),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_71),
.B1(n_89),
.B2(n_74),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_53),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_119),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_47),
.B1(n_42),
.B2(n_39),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_98),
.B1(n_116),
.B2(n_108),
.Y(n_136)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_11),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_2),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_132),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_134),
.B(n_120),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_90),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_86),
.C(n_75),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_73),
.B1(n_82),
.B2(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_71),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_117),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_62),
.C(n_73),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_103),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_74),
.B(n_4),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_3),
.B(n_5),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_82),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_95),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_168),
.C(n_146),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_100),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_153),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_97),
.B1(n_109),
.B2(n_104),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_151),
.B1(n_156),
.B2(n_167),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_97),
.B(n_117),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_119),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_165),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_114),
.B1(n_118),
.B2(n_105),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_160),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_78),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_39),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_135),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_142),
.B1(n_133),
.B2(n_138),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_141),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_153),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_183),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_168),
.C(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_188),
.C(n_192),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_149),
.C(n_143),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_159),
.B(n_149),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_170),
.B(n_169),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_157),
.B1(n_151),
.B2(n_159),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_173),
.B1(n_170),
.B2(n_169),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_174),
.C(n_172),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_128),
.C(n_161),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_197),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_SL g194 ( 
.A1(n_178),
.A2(n_161),
.A3(n_128),
.B1(n_137),
.B2(n_163),
.C1(n_147),
.C2(n_9),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_194),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_144),
.B(n_145),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_195),
.A2(n_171),
.B(n_179),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_205),
.B(n_189),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_181),
.A3(n_175),
.B1(n_182),
.B2(n_179),
.C1(n_176),
.C2(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_204),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_188),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_208),
.C(n_203),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_144),
.C(n_140),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_147),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_198),
.B(n_190),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_213),
.B(n_214),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_208),
.A2(n_198),
.B(n_196),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_191),
.B(n_193),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_206),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_200),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_SL g225 ( 
.A1(n_216),
.A2(n_130),
.B(n_6),
.C(n_7),
.Y(n_225)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_130),
.B1(n_5),
.B2(n_6),
.Y(n_224)
);

OAI221xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_147),
.C(n_130),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_145),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_221),
.A2(n_218),
.B(n_220),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_224),
.C(n_3),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_3),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_216),
.B(n_39),
.Y(n_230)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_228),
.B(n_8),
.CI(n_9),
.CON(n_229),
.SN(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_230),
.C(n_226),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_39),
.Y(n_232)
);


endmodule