module fake_jpeg_3710_n_440 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_2),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_53),
.Y(n_98)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_47),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_21),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_48),
.B(n_79),
.Y(n_137)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_64),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_68),
.Y(n_136)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_15),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_82),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_12),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx2_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_81),
.Y(n_127)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_85),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_14),
.Y(n_123)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_87),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_33),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_92),
.A2(n_81),
.B(n_80),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_22),
.B1(n_41),
.B2(n_32),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_93),
.A2(n_96),
.B1(n_102),
.B2(n_105),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_36),
.B1(n_30),
.B2(n_32),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_95),
.A2(n_107),
.B1(n_116),
.B2(n_121),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_59),
.A2(n_22),
.B1(n_32),
.B2(n_36),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_51),
.A2(n_22),
.B1(n_36),
.B2(n_43),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_31),
.B1(n_37),
.B2(n_30),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_46),
.A2(n_37),
.B1(n_34),
.B2(n_38),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_67),
.A2(n_34),
.B1(n_37),
.B2(n_28),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_71),
.A2(n_37),
.B1(n_34),
.B2(n_38),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_68),
.B1(n_2),
.B2(n_3),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_72),
.A2(n_50),
.B1(n_58),
.B2(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_131),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_69),
.A2(n_38),
.B1(n_33),
.B2(n_34),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_128),
.A2(n_68),
.B1(n_3),
.B2(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_12),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_83),
.A2(n_34),
.B1(n_33),
.B2(n_11),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_54),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_133),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_87),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_138),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_86),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_141),
.A2(n_146),
.B(n_149),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_142),
.B(n_152),
.Y(n_207)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_100),
.B(n_76),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_171),
.C(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_74),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_115),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_106),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_85),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_82),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_156),
.B(n_157),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_89),
.B(n_56),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_91),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_161),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

BUFx2_ASAP7_75t_SL g213 ( 
.A(n_160),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_88),
.B(n_0),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_173),
.B1(n_127),
.B2(n_136),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_98),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_167),
.Y(n_189)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_91),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_121),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_10),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_89),
.B(n_4),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_5),
.B(n_6),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_6),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_120),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_176),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_107),
.A2(n_6),
.B(n_7),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_125),
.B(n_97),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_126),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_179),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_129),
.B1(n_130),
.B2(n_110),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_183),
.B(n_192),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_184),
.B(n_149),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_145),
.A2(n_125),
.B1(n_132),
.B2(n_103),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_196),
.B1(n_201),
.B2(n_204),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_145),
.A2(n_103),
.B1(n_108),
.B2(n_104),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_147),
.A2(n_104),
.B1(n_108),
.B2(n_130),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_138),
.B1(n_178),
.B2(n_162),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_171),
.C(n_141),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_138),
.C(n_170),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_147),
.A2(n_110),
.B1(n_114),
.B2(n_129),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_241),
.C(n_245),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_154),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_220),
.B(n_227),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_192),
.A2(n_180),
.B1(n_158),
.B2(n_170),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_161),
.B1(n_111),
.B2(n_117),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_197),
.A2(n_155),
.B1(n_140),
.B2(n_148),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_150),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_165),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_228),
.B(n_229),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_155),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_216),
.B(n_199),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_152),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_231),
.B(n_232),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_187),
.B(n_163),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_208),
.A2(n_117),
.B1(n_111),
.B2(n_177),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_233),
.A2(n_214),
.B1(n_209),
.B2(n_198),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_184),
.B(n_179),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_234),
.B(n_235),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_143),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_237),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_194),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_215),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_149),
.B(n_153),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_247),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_151),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

OAI22x1_ASAP7_75t_L g243 ( 
.A1(n_183),
.A2(n_206),
.B1(n_185),
.B2(n_212),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_97),
.B1(n_168),
.B2(n_198),
.Y(n_279)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_126),
.C(n_151),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_196),
.A2(n_112),
.B1(n_144),
.B2(n_176),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_176),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_188),
.B(n_210),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_255),
.B(n_264),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_188),
.C(n_206),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_261),
.C(n_269),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_210),
.C(n_182),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_218),
.B(n_204),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_243),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_235),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_212),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_240),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_182),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_248),
.A2(n_201),
.B1(n_214),
.B2(n_209),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_270),
.A2(n_164),
.B1(n_181),
.B2(n_139),
.Y(n_307)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_279),
.B1(n_242),
.B2(n_245),
.Y(n_283)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_280),
.A2(n_285),
.B(n_293),
.Y(n_310)
);

BUFx4f_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_227),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_295),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_286),
.B1(n_297),
.B2(n_300),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_248),
.B(n_240),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_248),
.B1(n_219),
.B2(n_222),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_287),
.B(n_289),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_238),
.Y(n_290)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_291),
.B(n_271),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_229),
.C(n_231),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_302),
.C(n_305),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_268),
.A2(n_244),
.B(n_232),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_223),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_262),
.A2(n_219),
.B1(n_221),
.B2(n_243),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_299),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_271),
.A2(n_236),
.B1(n_224),
.B2(n_249),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_252),
.A2(n_247),
.B1(n_205),
.B2(n_233),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_239),
.C(n_99),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_266),
.B(n_247),
.Y(n_304)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_213),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_211),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_261),
.C(n_251),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_307),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_285),
.A2(n_252),
.B(n_268),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_309),
.A2(n_298),
.B(n_295),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_293),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_311),
.B(n_320),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_325),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_315),
.Y(n_336)
);

XOR2x2_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_267),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_250),
.C(n_278),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_323),
.C(n_324),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_256),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_253),
.C(n_277),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_257),
.C(n_253),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_257),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_294),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_333),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_250),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_331),
.C(n_303),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_252),
.C(n_272),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_SL g332 ( 
.A(n_286),
.B(n_258),
.C(n_270),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_301),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_290),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_321),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_338),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_328),
.A2(n_326),
.B1(n_313),
.B2(n_309),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_335),
.A2(n_341),
.B1(n_317),
.B2(n_312),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_314),
.B(n_306),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_296),
.C(n_275),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_319),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_281),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_344),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_328),
.A2(n_298),
.B1(n_304),
.B2(n_279),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_343),
.A2(n_354),
.B(n_322),
.Y(n_361)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_316),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_351),
.Y(n_369)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_330),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_349),
.Y(n_364)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_350),
.A2(n_343),
.B1(n_342),
.B2(n_347),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_281),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_284),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_352),
.B(n_296),
.Y(n_370)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_274),
.Y(n_374)
);

OAI211xp5_ASAP7_75t_SL g354 ( 
.A1(n_315),
.A2(n_327),
.B(n_332),
.C(n_322),
.Y(n_354)
);

AND2x2_ASAP7_75t_SL g355 ( 
.A(n_331),
.B(n_303),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_355),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_356),
.B(n_308),
.Y(n_365)
);

INVx13_ASAP7_75t_L g357 ( 
.A(n_334),
.Y(n_357)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_358),
.A2(n_338),
.B1(n_339),
.B2(n_344),
.Y(n_383)
);

AO21x1_ASAP7_75t_L g384 ( 
.A1(n_360),
.A2(n_361),
.B(n_366),
.Y(n_384)
);

BUFx12_ASAP7_75t_L g362 ( 
.A(n_351),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_362),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_368),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_335),
.A2(n_350),
.B(n_354),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_341),
.A2(n_324),
.B1(n_308),
.B2(n_307),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_367),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_336),
.B(n_258),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_371),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_346),
.B(n_345),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_336),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_340),
.B(n_356),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_340),
.C(n_355),
.Y(n_386)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_374),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_373),
.B(n_346),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_382),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_359),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_383),
.A2(n_369),
.B1(n_363),
.B2(n_357),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_355),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_389),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_386),
.B(n_375),
.Y(n_395)
);

AOI21x1_ASAP7_75t_L g397 ( 
.A1(n_388),
.A2(n_372),
.B(n_369),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_337),
.C(n_181),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_205),
.Y(n_390)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_390),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_134),
.C(n_136),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_378),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_360),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_393),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_359),
.C(n_364),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_399),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_366),
.B(n_361),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_390),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_397),
.A2(n_405),
.B(n_391),
.Y(n_413)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_398),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_368),
.C(n_362),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_362),
.C(n_134),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_404),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_176),
.Y(n_402)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_402),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_119),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_384),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_412),
.C(n_417),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_396),
.A2(n_381),
.B1(n_383),
.B2(n_377),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_411),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_400),
.B(n_403),
.C(n_393),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_378),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_413),
.B(n_416),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_211),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_398),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_418),
.A2(n_426),
.B(n_406),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_411),
.B(n_401),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_421),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_99),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_423),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_8),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_410),
.A2(n_211),
.B1(n_112),
.B2(n_94),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_425),
.A2(n_417),
.B(n_416),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_9),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_427),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_430),
.A2(n_431),
.B(n_432),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_424),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_SL g432 ( 
.A(n_419),
.B(n_412),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_428),
.B(n_420),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_435),
.A2(n_211),
.B1(n_9),
.B2(n_94),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_434),
.A2(n_426),
.B(n_429),
.Y(n_436)
);

BUFx24_ASAP7_75t_SL g438 ( 
.A(n_436),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_438),
.A2(n_433),
.B1(n_437),
.B2(n_9),
.Y(n_439)
);

BUFx24_ASAP7_75t_SL g440 ( 
.A(n_439),
.Y(n_440)
);


endmodule