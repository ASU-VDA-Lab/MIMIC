module fake_ariane_144_n_2343 (n_295, n_356, n_556, n_170, n_190, n_695, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_2343);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_695;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_2343;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_1174;
wire n_1469;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_1298;
wire n_737;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2233;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_2332;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_1819;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_1442;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2087;
wire n_931;
wire n_1491;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_2312;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2059;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1608;
wire n_1304;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_2075;
wire n_1726;
wire n_1945;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_951;
wire n_862;
wire n_1700;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_791;
wire n_876;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_1118;
wire n_943;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_819;
wire n_1971;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_911;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_1630;
wire n_1720;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_1393;
wire n_723;
wire n_2240;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx1_ASAP7_75t_L g697 ( 
.A(n_610),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_591),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_166),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_685),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_267),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_240),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_20),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_381),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_626),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_149),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_38),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_682),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_659),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_632),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_345),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_623),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_546),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_571),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_472),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_602),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_200),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_612),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_61),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_490),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_511),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_196),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_554),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_675),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_184),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_380),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_651),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_679),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_284),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_542),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_605),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_544),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_164),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_689),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_662),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_11),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_665),
.Y(n_737)
);

BUFx2_ASAP7_75t_SL g738 ( 
.A(n_424),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_695),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_684),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_151),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_535),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_582),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_155),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_619),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_581),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_310),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_638),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_598),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_377),
.Y(n_750)
);

BUFx10_ASAP7_75t_L g751 ( 
.A(n_495),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_256),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_280),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_693),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_529),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_423),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_661),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_69),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_173),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_119),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_419),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_222),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_629),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_164),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_22),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_47),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_635),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_322),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_586),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_232),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_522),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_60),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_337),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_247),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_170),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_631),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_116),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_11),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_126),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_523),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_393),
.Y(n_781)
);

BUFx10_ASAP7_75t_L g782 ( 
.A(n_7),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_676),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_374),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_540),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_108),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_482),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_95),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_174),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_485),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_408),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_663),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_493),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_594),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_156),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_539),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_525),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_609),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_668),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_297),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_42),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_628),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_413),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_620),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_611),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_205),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_75),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_669),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_690),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_28),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_18),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_578),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_468),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_607),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_6),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_677),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_124),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_647),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_146),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_670),
.Y(n_820)
);

CKINVDCx14_ASAP7_75t_R g821 ( 
.A(n_484),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_379),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_657),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_246),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_7),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_681),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_687),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_340),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_121),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_432),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_678),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_387),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_596),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_579),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_383),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_655),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_688),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_507),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_106),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_399),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_335),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_396),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_618),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_595),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_532),
.Y(n_845)
);

CKINVDCx16_ASAP7_75t_R g846 ( 
.A(n_403),
.Y(n_846)
);

CKINVDCx16_ASAP7_75t_R g847 ( 
.A(n_538),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_90),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_597),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_641),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_692),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_189),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_145),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_664),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_683),
.Y(n_855)
);

BUFx5_ASAP7_75t_L g856 ( 
.A(n_630),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_238),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_278),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_674),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_397),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_72),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_543),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_241),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_497),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_615),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_606),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_624),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_534),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_573),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_74),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_633),
.Y(n_871)
);

CKINVDCx16_ASAP7_75t_R g872 ( 
.A(n_653),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_167),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_572),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_518),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_364),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_374),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_479),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_272),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_414),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_395),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_308),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_622),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_85),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_658),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_95),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_437),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_645),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_672),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_239),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_29),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_302),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_666),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_694),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_296),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_634),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_671),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_382),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_648),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_639),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_509),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_646),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_691),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_356),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_299),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_660),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_643),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_621),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_262),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_12),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_563),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_642),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_644),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_526),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_640),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_404),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_82),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_617),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_288),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_503),
.Y(n_920)
);

CKINVDCx16_ASAP7_75t_R g921 ( 
.A(n_349),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_128),
.Y(n_922)
);

CKINVDCx14_ASAP7_75t_R g923 ( 
.A(n_105),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_94),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_114),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_608),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_62),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_452),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_189),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_177),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_393),
.Y(n_931)
);

BUFx10_ASAP7_75t_L g932 ( 
.A(n_604),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_41),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_652),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_467),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_21),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_149),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_625),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_680),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_656),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_404),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_545),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_367),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_472),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_116),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_577),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_461),
.Y(n_947)
);

CKINVDCx16_ASAP7_75t_R g948 ( 
.A(n_166),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_76),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_221),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_478),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_165),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_121),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_74),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_654),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_215),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_90),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_576),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_463),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_348),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_614),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_627),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_377),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_636),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_82),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_468),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_92),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_686),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_567),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_696),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_256),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_673),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_361),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_15),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_650),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_649),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_365),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_32),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_616),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_33),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_323),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_481),
.Y(n_982)
);

BUFx10_ASAP7_75t_L g983 ( 
.A(n_224),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_231),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_387),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_637),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_667),
.Y(n_987)
);

BUFx10_ASAP7_75t_L g988 ( 
.A(n_613),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_108),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_599),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_553),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_779),
.B(n_1),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_869),
.B(n_0),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_707),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_751),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_923),
.B(n_0),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_711),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_861),
.B(n_1),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_880),
.B(n_971),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_762),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_846),
.B(n_2),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_840),
.Y(n_1002)
);

AND2x6_ASAP7_75t_L g1003 ( 
.A(n_769),
.B(n_480),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_886),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_762),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_779),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_707),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_901),
.B(n_3),
.Y(n_1008)
);

BUFx12f_ASAP7_75t_L g1009 ( 
.A(n_751),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_707),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_744),
.B(n_2),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_782),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_786),
.B(n_3),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_925),
.Y(n_1014)
);

INVx5_ASAP7_75t_L g1015 ( 
.A(n_809),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_925),
.Y(n_1016)
);

BUFx12f_ASAP7_75t_L g1017 ( 
.A(n_809),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_925),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_909),
.B(n_4),
.Y(n_1019)
);

BUFx8_ASAP7_75t_SL g1020 ( 
.A(n_791),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_966),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_921),
.B(n_948),
.Y(n_1022)
);

INVx5_ASAP7_75t_L g1023 ( 
.A(n_920),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_920),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_697),
.B(n_4),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_1022),
.A2(n_996),
.B1(n_1001),
.B2(n_997),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_1004),
.B(n_701),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1006),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_994),
.Y(n_1029)
);

NOR2x1p5_ASAP7_75t_L g1030 ( 
.A(n_995),
.B(n_924),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_994),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1015),
.B(n_847),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1015),
.B(n_821),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1007),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_1023),
.B(n_872),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1010),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_996),
.A2(n_917),
.B1(n_937),
.B2(n_890),
.Y(n_1037)
);

OR2x6_ASAP7_75t_L g1038 ( 
.A(n_1009),
.B(n_738),
.Y(n_1038)
);

AO22x2_ASAP7_75t_L g1039 ( 
.A1(n_1001),
.A2(n_941),
.B1(n_729),
.B2(n_752),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1016),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1008),
.A2(n_954),
.B1(n_745),
.B2(n_754),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_1014),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_992),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1023),
.B(n_932),
.Y(n_1044)
);

AO22x2_ASAP7_75t_L g1045 ( 
.A1(n_999),
.A2(n_768),
.B1(n_817),
.B2(n_704),
.Y(n_1045)
);

AND2x2_ASAP7_75t_SL g1046 ( 
.A(n_998),
.B(n_736),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1014),
.Y(n_1047)
);

AND2x4_ASAP7_75t_SL g1048 ( 
.A(n_998),
.B(n_988),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1018),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1002),
.B(n_932),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_993),
.B(n_1017),
.Y(n_1051)
);

INVx8_ASAP7_75t_L g1052 ( 
.A(n_1024),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1018),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1021),
.B(n_955),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1025),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_1020),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1000),
.A2(n_793),
.B1(n_805),
.B2(n_700),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1048),
.B(n_1019),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1028),
.Y(n_1059)
);

XNOR2xp5_ASAP7_75t_L g1060 ( 
.A(n_1037),
.B(n_845),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1034),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1036),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_1043),
.B(n_1005),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1032),
.B(n_1012),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1040),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1055),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1029),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1047),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1049),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1033),
.B(n_1011),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1044),
.B(n_1013),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1031),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1042),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1050),
.B(n_782),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1046),
.A2(n_885),
.B(n_802),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1027),
.B(n_910),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1053),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1054),
.B(n_983),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1035),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1026),
.B(n_983),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1039),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1039),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1051),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1045),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1045),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1038),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1038),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_1052),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1057),
.B(n_957),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1052),
.Y(n_1090)
);

XOR2xp5_ASAP7_75t_L g1091 ( 
.A(n_1056),
.B(n_1041),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_1032),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_1027),
.B(n_967),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1028),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_1030),
.B(n_718),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1043),
.B(n_698),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1028),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1028),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1028),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_1056),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1048),
.B(n_815),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_SL g1102 ( 
.A(n_1052),
.B(n_911),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1098),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_1100),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1074),
.B(n_907),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1066),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1092),
.B(n_749),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1061),
.Y(n_1108)
);

AND2x6_ASAP7_75t_L g1109 ( 
.A(n_1058),
.B(n_705),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1059),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1096),
.B(n_794),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1078),
.B(n_876),
.Y(n_1112)
);

INVx3_ASAP7_75t_SL g1113 ( 
.A(n_1088),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1076),
.B(n_884),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1094),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_1093),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1097),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_1101),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1101),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1099),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1090),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1062),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1083),
.B(n_699),
.Y(n_1123)
);

AND2x2_ASAP7_75t_SL g1124 ( 
.A(n_1080),
.B(n_760),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_1058),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1065),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1072),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_1060),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1086),
.B(n_702),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_1095),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_1068),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1089),
.B(n_706),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1079),
.B(n_703),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1067),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1075),
.A2(n_728),
.B(n_714),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1063),
.B(n_719),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1064),
.B(n_715),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1073),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1087),
.B(n_726),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1069),
.Y(n_1140)
);

BUFx12f_ASAP7_75t_SL g1141 ( 
.A(n_1091),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1077),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1071),
.B(n_804),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1070),
.B(n_747),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1081),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1081),
.Y(n_1146)
);

INVx4_ASAP7_75t_L g1147 ( 
.A(n_1082),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1084),
.B(n_753),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1085),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1092),
.B(n_936),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_1058),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1092),
.B(n_936),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1098),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1058),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1088),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1083),
.B(n_984),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_1058),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1076),
.B(n_825),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1088),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1092),
.B(n_936),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1074),
.B(n_766),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1058),
.B(n_773),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1098),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1074),
.B(n_775),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1098),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1083),
.B(n_717),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1098),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1100),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1058),
.B(n_778),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1074),
.B(n_784),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1101),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1100),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1066),
.Y(n_1173)
);

NOR2xp67_ASAP7_75t_L g1174 ( 
.A(n_1088),
.B(n_730),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1058),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1096),
.A2(n_757),
.B(n_748),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1092),
.B(n_722),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1100),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1058),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1100),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1074),
.B(n_807),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_1058),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_1100),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1092),
.B(n_725),
.Y(n_1184)
);

NOR2xp67_ASAP7_75t_L g1185 ( 
.A(n_1088),
.B(n_982),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_1088),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1083),
.B(n_733),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1074),
.B(n_830),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1074),
.B(n_835),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1088),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1100),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1074),
.B(n_839),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1058),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1098),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1102),
.B(n_955),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1066),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1092),
.B(n_741),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1145),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1153),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1165),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1111),
.B(n_841),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1167),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1183),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1104),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1191),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1119),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1168),
.B(n_848),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_1151),
.B(n_781),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1106),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1116),
.B(n_1114),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1194),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1105),
.B(n_852),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1106),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1125),
.B(n_750),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1113),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1112),
.B(n_873),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1180),
.B(n_882),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_SL g1218 ( 
.A(n_1195),
.B(n_988),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1137),
.B(n_891),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1173),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1107),
.B(n_1136),
.Y(n_1221)
);

INVx6_ASAP7_75t_L g1222 ( 
.A(n_1172),
.Y(n_1222)
);

INVx6_ASAP7_75t_L g1223 ( 
.A(n_1178),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1173),
.Y(n_1224)
);

BUFx2_ASAP7_75t_SL g1225 ( 
.A(n_1154),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1190),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1157),
.B(n_904),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1123),
.B(n_922),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1175),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1176),
.B(n_935),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1179),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1196),
.B(n_947),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1196),
.B(n_949),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1182),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1161),
.B(n_953),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1144),
.B(n_960),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1171),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1118),
.B(n_756),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1193),
.B(n_973),
.Y(n_1239)
);

AND2x6_ASAP7_75t_L g1240 ( 
.A(n_1146),
.B(n_771),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1108),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1143),
.B(n_974),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1141),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_L g1244 ( 
.A(n_1121),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1110),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1130),
.B(n_977),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1121),
.B(n_985),
.Y(n_1247)
);

NAND2x1_ASAP7_75t_SL g1248 ( 
.A(n_1132),
.B(n_783),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1164),
.B(n_758),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1170),
.B(n_759),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1158),
.B(n_761),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1117),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_1181),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1186),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1131),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1124),
.B(n_764),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1155),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1128),
.B(n_765),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1120),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1188),
.B(n_770),
.Y(n_1260)
);

AND2x2_ASAP7_75t_SL g1261 ( 
.A(n_1147),
.B(n_801),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1159),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1115),
.Y(n_1263)
);

AND2x4_ASAP7_75t_SL g1264 ( 
.A(n_1162),
.B(n_832),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1189),
.B(n_772),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1169),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1169),
.B(n_898),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1177),
.B(n_774),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1129),
.Y(n_1269)
);

BUFx2_ASAP7_75t_SL g1270 ( 
.A(n_1109),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1126),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1122),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1109),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1134),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1192),
.B(n_777),
.Y(n_1275)
);

OR2x6_ASAP7_75t_L g1276 ( 
.A(n_1149),
.B(n_944),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1129),
.B(n_959),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1139),
.B(n_1148),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1127),
.Y(n_1279)
);

BUFx4f_ASAP7_75t_L g1280 ( 
.A(n_1109),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1184),
.B(n_788),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1139),
.B(n_1103),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1163),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1134),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1140),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1142),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1133),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1174),
.B(n_980),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1138),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1150),
.Y(n_1290)
);

BUFx8_ASAP7_75t_SL g1291 ( 
.A(n_1197),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1152),
.Y(n_1292)
);

OR2x6_ASAP7_75t_L g1293 ( 
.A(n_1185),
.B(n_989),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1135),
.B(n_789),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1156),
.B(n_1166),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1187),
.B(n_798),
.Y(n_1296)
);

NOR2x1_ASAP7_75t_L g1297 ( 
.A(n_1160),
.B(n_818),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1111),
.B(n_795),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_SL g1299 ( 
.A(n_1191),
.B(n_800),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1111),
.B(n_803),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1153),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1183),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1145),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1153),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1125),
.B(n_866),
.Y(n_1305)
);

BUFx12f_ASAP7_75t_L g1306 ( 
.A(n_1191),
.Y(n_1306)
);

INVx5_ASAP7_75t_L g1307 ( 
.A(n_1190),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1145),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1116),
.B(n_806),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1104),
.B(n_833),
.Y(n_1310)
);

OR2x6_ASAP7_75t_L g1311 ( 
.A(n_1151),
.B(n_938),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1104),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1183),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1111),
.B(n_810),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_SL g1315 ( 
.A(n_1191),
.B(n_811),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1153),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1104),
.B(n_837),
.Y(n_1317)
);

NOR2x1_ASAP7_75t_L g1318 ( 
.A(n_1130),
.B(n_843),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1153),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1180),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1104),
.B(n_851),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1116),
.B(n_813),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1153),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1119),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1111),
.B(n_819),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_SL g1326 ( 
.A(n_1191),
.B(n_822),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1104),
.B(n_844),
.Y(n_1327)
);

BUFx8_ASAP7_75t_SL g1328 ( 
.A(n_1183),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1111),
.B(n_824),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1145),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1153),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1111),
.B(n_828),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1111),
.B(n_829),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1210),
.B(n_1278),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1320),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1241),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1209),
.Y(n_1337)
);

INVx3_ASAP7_75t_SL g1338 ( 
.A(n_1222),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1328),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1223),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1204),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1204),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1213),
.Y(n_1343)
);

NAND2x1p5_ASAP7_75t_L g1344 ( 
.A(n_1307),
.B(n_942),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1220),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1221),
.B(n_842),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1203),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1312),
.Y(n_1348)
);

BUFx2_ASAP7_75t_SL g1349 ( 
.A(n_1243),
.Y(n_1349)
);

NAND2x1p5_ASAP7_75t_L g1350 ( 
.A(n_1244),
.B(n_961),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1313),
.Y(n_1351)
);

BUFx12f_ASAP7_75t_L g1352 ( 
.A(n_1306),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1224),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1215),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1266),
.B(n_855),
.Y(n_1355)
);

NAND2x1p5_ASAP7_75t_L g1356 ( 
.A(n_1312),
.B(n_859),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1245),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1226),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1226),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_SL g1360 ( 
.A(n_1207),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1263),
.Y(n_1361)
);

CKINVDCx16_ASAP7_75t_R g1362 ( 
.A(n_1299),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1302),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1237),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1205),
.Y(n_1365)
);

BUFx24_ASAP7_75t_L g1366 ( 
.A(n_1310),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_R g1367 ( 
.A(n_1315),
.B(n_1326),
.Y(n_1367)
);

INVx5_ASAP7_75t_L g1368 ( 
.A(n_1255),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1279),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1253),
.B(n_853),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1198),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1256),
.A2(n_858),
.B1(n_860),
.B2(n_857),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1229),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1283),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1229),
.Y(n_1375)
);

INVx6_ASAP7_75t_SL g1376 ( 
.A(n_1208),
.Y(n_1376)
);

INVx6_ASAP7_75t_SL g1377 ( 
.A(n_1267),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1287),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1303),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1309),
.B(n_863),
.Y(n_1380)
);

INVx3_ASAP7_75t_SL g1381 ( 
.A(n_1317),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1257),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1280),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1262),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1231),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1284),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1308),
.Y(n_1387)
);

BUFx4_ASAP7_75t_SL g1388 ( 
.A(n_1293),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1330),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1219),
.B(n_978),
.Y(n_1390)
);

OR2x6_ASAP7_75t_L g1391 ( 
.A(n_1270),
.B(n_867),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1291),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1285),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1234),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1286),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1212),
.B(n_870),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1234),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1225),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1269),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1252),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1322),
.B(n_1251),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1274),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1259),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1254),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1282),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1272),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1261),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1271),
.Y(n_1408)
);

INVx5_ASAP7_75t_L g1409 ( 
.A(n_1240),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1199),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1200),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1247),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1202),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1311),
.Y(n_1414)
);

INVx5_ASAP7_75t_L g1415 ( 
.A(n_1240),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1264),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1324),
.B(n_868),
.Y(n_1417)
);

INVx8_ASAP7_75t_L g1418 ( 
.A(n_1276),
.Y(n_1418)
);

BUFx5_ASAP7_75t_L g1419 ( 
.A(n_1240),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1258),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1321),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1217),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1246),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1211),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1268),
.A2(n_878),
.B1(n_879),
.B2(n_877),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1327),
.Y(n_1426)
);

BUFx2_ASAP7_75t_SL g1427 ( 
.A(n_1273),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1305),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1277),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1281),
.B(n_881),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1248),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1206),
.B(n_883),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1395),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1364),
.Y(n_1434)
);

INVx4_ASAP7_75t_SL g1435 ( 
.A(n_1338),
.Y(n_1435)
);

BUFx12f_ASAP7_75t_L g1436 ( 
.A(n_1378),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1412),
.A2(n_1238),
.B1(n_1218),
.B2(n_1214),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1400),
.Y(n_1438)
);

AOI22x1_ASAP7_75t_SL g1439 ( 
.A1(n_1392),
.A2(n_892),
.B1(n_895),
.B2(n_887),
.Y(n_1439)
);

INVx3_ASAP7_75t_SL g1440 ( 
.A(n_1398),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1352),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1422),
.A2(n_1239),
.B1(n_1227),
.B2(n_1294),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1403),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1374),
.Y(n_1444)
);

BUFx4f_ASAP7_75t_SL g1445 ( 
.A(n_1351),
.Y(n_1445)
);

INVx5_ASAP7_75t_L g1446 ( 
.A(n_1339),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1430),
.A2(n_1228),
.B1(n_1333),
.B2(n_1332),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1406),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1407),
.A2(n_1296),
.B1(n_1304),
.B2(n_1301),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1408),
.Y(n_1450)
);

BUFx10_ASAP7_75t_L g1451 ( 
.A(n_1340),
.Y(n_1451)
);

INVx6_ASAP7_75t_L g1452 ( 
.A(n_1368),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1375),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1357),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1368),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1425),
.A2(n_1300),
.B(n_1298),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1390),
.A2(n_1325),
.B1(n_1329),
.B2(n_1314),
.Y(n_1457)
);

BUFx8_ASAP7_75t_L g1458 ( 
.A(n_1360),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1367),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1401),
.A2(n_1230),
.B1(n_1275),
.B2(n_1289),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1407),
.A2(n_1319),
.B1(n_1323),
.B2(n_1316),
.Y(n_1461)
);

INVxp67_ASAP7_75t_SL g1462 ( 
.A(n_1405),
.Y(n_1462)
);

OAI21xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1336),
.A2(n_1343),
.B(n_1337),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1365),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1342),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1361),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1348),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1345),
.Y(n_1468)
);

CKINVDCx11_ASAP7_75t_R g1469 ( 
.A(n_1381),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1396),
.A2(n_1331),
.B1(n_1216),
.B2(n_1235),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_R g1471 ( 
.A1(n_1380),
.A2(n_956),
.B1(n_981),
.B2(n_927),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1362),
.Y(n_1472)
);

CKINVDCx6p67_ASAP7_75t_R g1473 ( 
.A(n_1366),
.Y(n_1473)
);

CKINVDCx11_ASAP7_75t_R g1474 ( 
.A(n_1426),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1373),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1420),
.A2(n_1250),
.B1(n_1260),
.B2(n_1249),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1353),
.Y(n_1477)
);

INVx8_ASAP7_75t_L g1478 ( 
.A(n_1418),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1341),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1346),
.A2(n_1265),
.B1(n_1201),
.B2(n_1295),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1373),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1377),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1334),
.B(n_1236),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1355),
.A2(n_1288),
.B1(n_1318),
.B2(n_1290),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1382),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1369),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1335),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1405),
.B(n_1242),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1372),
.A2(n_1233),
.B1(n_1232),
.B2(n_1297),
.Y(n_1489)
);

BUFx8_ASAP7_75t_SL g1490 ( 
.A(n_1363),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1385),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1384),
.Y(n_1492)
);

BUFx10_ASAP7_75t_L g1493 ( 
.A(n_1417),
.Y(n_1493)
);

CKINVDCx6p67_ASAP7_75t_R g1494 ( 
.A(n_1421),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1359),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1371),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1349),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1409),
.A2(n_1292),
.B1(n_930),
.B2(n_916),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1409),
.A2(n_951),
.B1(n_933),
.B2(n_919),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1376),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1415),
.A2(n_928),
.B1(n_929),
.B2(n_905),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1393),
.Y(n_1502)
);

CKINVDCx14_ASAP7_75t_R g1503 ( 
.A(n_1414),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1388),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1347),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1402),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1399),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1432),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1423),
.A2(n_943),
.B1(n_945),
.B2(n_931),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1410),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1411),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1397),
.Y(n_1512)
);

BUFx8_ASAP7_75t_SL g1513 ( 
.A(n_1354),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1415),
.A2(n_952),
.B1(n_963),
.B2(n_950),
.Y(n_1514)
);

NAND2x1p5_ASAP7_75t_L g1515 ( 
.A(n_1358),
.B(n_888),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1429),
.A2(n_965),
.B1(n_1003),
.B2(n_899),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1379),
.A2(n_964),
.B1(n_889),
.B2(n_913),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1387),
.Y(n_1518)
);

INVx6_ASAP7_75t_L g1519 ( 
.A(n_1399),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1389),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1394),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1404),
.A2(n_1370),
.B1(n_1391),
.B2(n_1356),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1419),
.A2(n_918),
.B1(n_934),
.B2(n_900),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1386),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1416),
.B(n_1003),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1428),
.Y(n_1526)
);

OAI21xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1424),
.A2(n_940),
.B(n_939),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1431),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1383),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1413),
.B(n_958),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1427),
.A2(n_976),
.B1(n_979),
.B2(n_975),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1419),
.A2(n_716),
.B1(n_735),
.B2(n_727),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1344),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1350),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1419),
.A2(n_755),
.B1(n_767),
.B2(n_739),
.Y(n_1535)
);

INVx5_ASAP7_75t_L g1536 ( 
.A(n_1352),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1400),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1338),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1459),
.B(n_1473),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1471),
.A2(n_962),
.B1(n_769),
.B2(n_856),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1448),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1456),
.A2(n_709),
.B1(n_710),
.B2(n_708),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1434),
.B(n_5),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1480),
.A2(n_962),
.B1(n_856),
.B2(n_713),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1460),
.A2(n_856),
.B1(n_720),
.B2(n_721),
.Y(n_1545)
);

OAI21xp33_ASAP7_75t_L g1546 ( 
.A1(n_1447),
.A2(n_723),
.B(n_712),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1433),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1483),
.A2(n_731),
.B1(n_732),
.B2(n_724),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1476),
.A2(n_737),
.B1(n_740),
.B2(n_734),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1467),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1437),
.A2(n_743),
.B1(n_746),
.B2(n_742),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1496),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1442),
.A2(n_856),
.B1(n_776),
.B2(n_780),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1502),
.B(n_5),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1452),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1470),
.B(n_6),
.Y(n_1556)
);

AOI222xp33_ASAP7_75t_L g1557 ( 
.A1(n_1457),
.A2(n_790),
.B1(n_785),
.B2(n_792),
.C1(n_787),
.C2(n_763),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1538),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1465),
.B(n_8),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1489),
.A2(n_856),
.B1(n_797),
.B2(n_799),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1484),
.A2(n_808),
.B1(n_812),
.B2(n_796),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1493),
.A2(n_816),
.B1(n_820),
.B2(n_814),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1535),
.A2(n_826),
.B1(n_827),
.B2(n_823),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1508),
.A2(n_834),
.B1(n_836),
.B2(n_831),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1518),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1499),
.A2(n_8),
.B(n_9),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1454),
.A2(n_849),
.B1(n_850),
.B2(n_838),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1444),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1523),
.A2(n_864),
.B1(n_865),
.B2(n_854),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1488),
.B(n_9),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1522),
.B(n_862),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1467),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1507),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1466),
.A2(n_874),
.B1(n_875),
.B2(n_871),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1520),
.Y(n_1575)
);

BUFx12f_ASAP7_75t_L g1576 ( 
.A(n_1441),
.Y(n_1576)
);

INVx2_ASAP7_75t_SL g1577 ( 
.A(n_1478),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1505),
.A2(n_1497),
.B1(n_1531),
.B2(n_1464),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1527),
.A2(n_894),
.B1(n_896),
.B2(n_893),
.Y(n_1579)
);

INVx4_ASAP7_75t_L g1580 ( 
.A(n_1435),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1517),
.A2(n_902),
.B1(n_903),
.B2(n_897),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1510),
.A2(n_908),
.B1(n_912),
.B2(n_906),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1511),
.A2(n_915),
.B1(n_926),
.B2(n_914),
.Y(n_1583)
);

AOI222xp33_ASAP7_75t_L g1584 ( 
.A1(n_1438),
.A2(n_970),
.B1(n_968),
.B2(n_972),
.C1(n_969),
.C2(n_946),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1443),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1450),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1537),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1515),
.A2(n_987),
.B1(n_991),
.B2(n_986),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1490),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1455),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1468),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1528),
.A2(n_990),
.B1(n_13),
.B2(n_10),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1477),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1487),
.B(n_10),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_L g1595 ( 
.A(n_1463),
.B(n_12),
.C(n_13),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1449),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1486),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1538),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1501),
.A2(n_17),
.B(n_18),
.Y(n_1599)
);

BUFx4f_ASAP7_75t_SL g1600 ( 
.A(n_1436),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1478),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1530),
.Y(n_1602)
);

AOI222xp33_ASAP7_75t_L g1603 ( 
.A1(n_1472),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.C1(n_20),
.C2(n_22),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1446),
.A2(n_24),
.B1(n_19),
.B2(n_23),
.Y(n_1604)
);

OAI222xp33_ASAP7_75t_L g1605 ( 
.A1(n_1439),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.C1(n_25),
.C2(n_27),
.Y(n_1605)
);

OAI21xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1516),
.A2(n_25),
.B(n_26),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1461),
.A2(n_31),
.B1(n_27),
.B2(n_30),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1462),
.B(n_34),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1512),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1532),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1533),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1533),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1492),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1524),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1521),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1526),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1509),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1506),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1609),
.Y(n_1619)
);

AOI211xp5_ASAP7_75t_L g1620 ( 
.A1(n_1605),
.A2(n_1514),
.B(n_1440),
.C(n_1529),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1552),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1599),
.A2(n_1445),
.B1(n_1536),
.B2(n_1498),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1566),
.A2(n_1504),
.B1(n_1494),
.B2(n_1534),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1540),
.A2(n_1458),
.B1(n_1479),
.B2(n_1495),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1602),
.A2(n_1546),
.B1(n_1557),
.B2(n_1556),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1565),
.Y(n_1626)
);

AOI222xp33_ASAP7_75t_L g1627 ( 
.A1(n_1617),
.A2(n_1474),
.B1(n_1469),
.B2(n_1500),
.C1(n_1482),
.C2(n_1453),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1597),
.Y(n_1628)
);

OAI222xp33_ASAP7_75t_L g1629 ( 
.A1(n_1545),
.A2(n_1503),
.B1(n_1525),
.B2(n_1481),
.C1(n_1491),
.C2(n_1475),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1616),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1560),
.A2(n_1479),
.B1(n_1519),
.B2(n_1485),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1570),
.B(n_1615),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1575),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1595),
.A2(n_1513),
.B1(n_1451),
.B2(n_46),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1603),
.A2(n_1544),
.B1(n_1568),
.B2(n_1547),
.Y(n_1635)
);

OAI222xp33_ASAP7_75t_L g1636 ( 
.A1(n_1613),
.A2(n_50),
.B1(n_52),
.B2(n_48),
.C1(n_49),
.C2(n_51),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1541),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1571),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1638)
);

OA222x2_ASAP7_75t_L g1639 ( 
.A1(n_1543),
.A2(n_1554),
.B1(n_1558),
.B2(n_1586),
.C1(n_1587),
.C2(n_1585),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1606),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1640)
);

OA21x2_ASAP7_75t_L g1641 ( 
.A1(n_1591),
.A2(n_56),
.B(n_57),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1610),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1553),
.A2(n_61),
.B1(n_58),
.B2(n_59),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1593),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1584),
.A2(n_1542),
.B1(n_1578),
.B2(n_1592),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1608),
.A2(n_63),
.B1(n_59),
.B2(n_62),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1611),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1559),
.B(n_67),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1612),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1596),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1604),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1607),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1579),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1653)
);

OAI222xp33_ASAP7_75t_L g1654 ( 
.A1(n_1594),
.A2(n_79),
.B1(n_81),
.B2(n_77),
.C1(n_78),
.C2(n_80),
.Y(n_1654)
);

OAI222xp33_ASAP7_75t_L g1655 ( 
.A1(n_1551),
.A2(n_83),
.B1(n_85),
.B2(n_80),
.C1(n_81),
.C2(n_84),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_SL g1656 ( 
.A1(n_1588),
.A2(n_93),
.B1(n_102),
.B2(n_83),
.Y(n_1656)
);

OAI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1581),
.A2(n_1563),
.B1(n_1561),
.B2(n_1564),
.C(n_1562),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1548),
.A2(n_87),
.B1(n_84),
.B2(n_86),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1549),
.A2(n_89),
.B1(n_86),
.B2(n_88),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1569),
.A2(n_91),
.B1(n_88),
.B2(n_89),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1618),
.B(n_91),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1576),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_1662)
);

NAND3xp33_ASAP7_75t_L g1663 ( 
.A(n_1567),
.B(n_96),
.C(n_97),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1574),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1664)
);

OAI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1539),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1573),
.B(n_99),
.Y(n_1666)
);

OAI222xp33_ASAP7_75t_L g1667 ( 
.A1(n_1580),
.A2(n_104),
.B1(n_106),
.B2(n_101),
.C1(n_103),
.C2(n_105),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1580),
.A2(n_107),
.B1(n_103),
.B2(n_104),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1582),
.A2(n_110),
.B1(n_107),
.B2(n_109),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1583),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1598),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1550),
.Y(n_1672)
);

OAI21xp33_ASAP7_75t_SL g1673 ( 
.A1(n_1577),
.A2(n_1601),
.B(n_1590),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1614),
.A2(n_118),
.B1(n_115),
.B2(n_117),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1573),
.A2(n_125),
.B1(n_133),
.B2(n_115),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1555),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.C(n_120),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1550),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1550),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1572),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1572),
.A2(n_1600),
.B1(n_1589),
.B2(n_127),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1572),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1556),
.A2(n_133),
.B1(n_141),
.B2(n_125),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1556),
.A2(n_135),
.B1(n_143),
.B2(n_126),
.Y(n_1683)
);

AND2x2_ASAP7_75t_SL g1684 ( 
.A(n_1639),
.B(n_127),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1630),
.B(n_128),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1619),
.B(n_129),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_R g1687 ( 
.A(n_1648),
.B(n_1672),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_L g1688 ( 
.A(n_1676),
.B(n_130),
.C(n_131),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1621),
.B(n_1626),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1632),
.B(n_130),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1633),
.B(n_131),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1644),
.B(n_132),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1645),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1662),
.A2(n_137),
.B1(n_134),
.B2(n_136),
.C(n_138),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1677),
.B(n_137),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1661),
.B(n_138),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1679),
.B(n_139),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1625),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1628),
.B(n_140),
.Y(n_1699)
);

OAI221xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1620),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.C(n_145),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_1663),
.B(n_1646),
.C(n_1656),
.Y(n_1701)
);

NOR3xp33_ASAP7_75t_SL g1702 ( 
.A(n_1674),
.B(n_144),
.C(n_146),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1654),
.A2(n_150),
.B1(n_147),
.B2(n_148),
.C(n_151),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1681),
.B(n_147),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1682),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1641),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1683),
.B(n_152),
.Y(n_1707)
);

NAND3xp33_ASAP7_75t_L g1708 ( 
.A(n_1668),
.B(n_153),
.C(n_154),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1623),
.B(n_1635),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1627),
.B(n_155),
.Y(n_1710)
);

AOI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1667),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.C(n_159),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1671),
.B(n_157),
.C(n_158),
.Y(n_1712)
);

NOR3xp33_ASAP7_75t_L g1713 ( 
.A(n_1655),
.B(n_159),
.C(n_160),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1675),
.B(n_160),
.C(n_161),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1665),
.B(n_161),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1622),
.B(n_1627),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1680),
.B(n_162),
.Y(n_1717)
);

OA21x2_ASAP7_75t_L g1718 ( 
.A1(n_1636),
.A2(n_162),
.B(n_163),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_L g1719 ( 
.A(n_1660),
.B(n_165),
.C(n_168),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_R g1720 ( 
.A(n_1631),
.B(n_168),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1634),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_1721)
);

NAND2xp33_ASAP7_75t_SL g1722 ( 
.A(n_1651),
.B(n_169),
.Y(n_1722)
);

OAI22xp33_ASAP7_75t_SL g1723 ( 
.A1(n_1653),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1640),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1637),
.B(n_178),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1659),
.B(n_178),
.C(n_179),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1678),
.B(n_179),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1642),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1658),
.B(n_180),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1664),
.B(n_181),
.Y(n_1730)
);

NOR2xp67_ASAP7_75t_L g1731 ( 
.A(n_1624),
.B(n_1647),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1638),
.B(n_183),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1669),
.B(n_183),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1670),
.B(n_184),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1650),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1643),
.B(n_186),
.C(n_187),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1652),
.B(n_188),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1649),
.B(n_188),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1629),
.B(n_190),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1657),
.B(n_190),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1627),
.A2(n_191),
.B(n_192),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1673),
.B(n_191),
.Y(n_1742)
);

OAI21xp33_ASAP7_75t_L g1743 ( 
.A1(n_1668),
.A2(n_193),
.B(n_194),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1676),
.B(n_193),
.C(n_194),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1630),
.B(n_195),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1620),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1673),
.B(n_197),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1632),
.B(n_198),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1630),
.B(n_198),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1673),
.B(n_199),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1645),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_1751)
);

OAI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1620),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.C(n_204),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1627),
.A2(n_202),
.B(n_203),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1673),
.B(n_204),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1673),
.B(n_206),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1632),
.B(n_206),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1630),
.B(n_207),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1673),
.B(n_208),
.Y(n_1758)
);

NAND3xp33_ASAP7_75t_L g1759 ( 
.A(n_1676),
.B(n_208),
.C(n_209),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_SL g1760 ( 
.A1(n_1641),
.A2(n_209),
.B(n_210),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_SL g1761 ( 
.A(n_1700),
.B(n_210),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1687),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1689),
.B(n_211),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1690),
.B(n_212),
.Y(n_1764)
);

OA211x2_ASAP7_75t_L g1765 ( 
.A1(n_1716),
.A2(n_223),
.B(n_231),
.C(n_213),
.Y(n_1765)
);

AOI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1740),
.A2(n_217),
.B1(n_214),
.B2(n_216),
.C(n_218),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1713),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1685),
.Y(n_1768)
);

NOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1745),
.B(n_219),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1692),
.Y(n_1770)
);

NAND3xp33_ASAP7_75t_L g1771 ( 
.A(n_1746),
.B(n_220),
.C(n_221),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1749),
.B(n_220),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1757),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1696),
.B(n_223),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1699),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1748),
.B(n_224),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1752),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1741),
.B(n_225),
.C(n_226),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_SL g1779 ( 
.A(n_1753),
.B(n_227),
.C(n_228),
.Y(n_1779)
);

NAND4xp75_ASAP7_75t_L g1780 ( 
.A(n_1710),
.B(n_230),
.C(n_228),
.D(n_229),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1708),
.B(n_230),
.C(n_232),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1691),
.B(n_233),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1756),
.B(n_233),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1709),
.B(n_234),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1704),
.B(n_1695),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1720),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1697),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1701),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1739),
.B(n_1718),
.Y(n_1789)
);

NAND4xp75_ASAP7_75t_L g1790 ( 
.A(n_1731),
.B(n_237),
.C(n_235),
.D(n_236),
.Y(n_1790)
);

AND2x4_ASAP7_75t_SL g1791 ( 
.A(n_1717),
.B(n_1702),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1742),
.B(n_239),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1747),
.B(n_240),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1712),
.B(n_241),
.C(n_242),
.Y(n_1794)
);

AOI211xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1723),
.A2(n_244),
.B(n_242),
.C(n_243),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1750),
.B(n_243),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1718),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1760),
.B(n_245),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1754),
.B(n_247),
.Y(n_1799)
);

NAND3xp33_ASAP7_75t_L g1800 ( 
.A(n_1703),
.B(n_248),
.C(n_249),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1711),
.B(n_248),
.C(n_249),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1722),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_1802)
);

NAND4xp75_ASAP7_75t_L g1803 ( 
.A(n_1755),
.B(n_252),
.C(n_250),
.D(n_251),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1758),
.B(n_1715),
.Y(n_1804)
);

NAND4xp75_ASAP7_75t_L g1805 ( 
.A(n_1707),
.B(n_255),
.C(n_253),
.D(n_254),
.Y(n_1805)
);

AOI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1723),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1725),
.Y(n_1807)
);

OA211x2_ASAP7_75t_L g1808 ( 
.A1(n_1743),
.A2(n_265),
.B(n_274),
.C(n_257),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1751),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_1809)
);

NOR3xp33_ASAP7_75t_L g1810 ( 
.A(n_1694),
.B(n_258),
.C(n_259),
.Y(n_1810)
);

NAND4xp25_ASAP7_75t_L g1811 ( 
.A(n_1721),
.B(n_262),
.C(n_260),
.D(n_261),
.Y(n_1811)
);

NOR2x1_ASAP7_75t_L g1812 ( 
.A(n_1714),
.B(n_261),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1698),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.C(n_266),
.Y(n_1813)
);

NAND3xp33_ASAP7_75t_L g1814 ( 
.A(n_1688),
.B(n_264),
.C(n_266),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1729),
.B(n_268),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1737),
.B(n_1730),
.Y(n_1816)
);

NAND3xp33_ASAP7_75t_L g1817 ( 
.A(n_1744),
.B(n_268),
.C(n_269),
.Y(n_1817)
);

OAI211xp5_ASAP7_75t_L g1818 ( 
.A1(n_1728),
.A2(n_1735),
.B(n_1738),
.C(n_1759),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_L g1819 ( 
.A(n_1719),
.B(n_269),
.C(n_270),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1734),
.B(n_271),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1727),
.B(n_272),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1733),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1693),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_1823)
);

NAND3xp33_ASAP7_75t_L g1824 ( 
.A(n_1726),
.B(n_275),
.C(n_276),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1736),
.B(n_276),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1705),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1724),
.B(n_277),
.Y(n_1827)
);

NAND3xp33_ASAP7_75t_L g1828 ( 
.A(n_1732),
.B(n_278),
.C(n_279),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1689),
.B(n_279),
.Y(n_1829)
);

AO21x2_ASAP7_75t_L g1830 ( 
.A1(n_1706),
.A2(n_280),
.B(n_281),
.Y(n_1830)
);

XOR2x2_ASAP7_75t_L g1831 ( 
.A(n_1684),
.B(n_282),
.Y(n_1831)
);

AO21x2_ASAP7_75t_L g1832 ( 
.A1(n_1706),
.A2(n_283),
.B(n_284),
.Y(n_1832)
);

NOR2x1_ASAP7_75t_L g1833 ( 
.A(n_1686),
.B(n_283),
.Y(n_1833)
);

NAND4xp75_ASAP7_75t_L g1834 ( 
.A(n_1684),
.B(n_287),
.C(n_285),
.D(n_286),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1687),
.B(n_285),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1689),
.B(n_287),
.Y(n_1836)
);

NOR3xp33_ASAP7_75t_L g1837 ( 
.A(n_1741),
.B(n_288),
.C(n_289),
.Y(n_1837)
);

NOR3xp33_ASAP7_75t_L g1838 ( 
.A(n_1741),
.B(n_289),
.C(n_290),
.Y(n_1838)
);

INVxp67_ASAP7_75t_SL g1839 ( 
.A(n_1773),
.Y(n_1839)
);

XOR2x2_ASAP7_75t_L g1840 ( 
.A(n_1831),
.B(n_290),
.Y(n_1840)
);

NOR3xp33_ASAP7_75t_SL g1841 ( 
.A(n_1779),
.B(n_1778),
.C(n_1818),
.Y(n_1841)
);

NOR4xp25_ASAP7_75t_L g1842 ( 
.A(n_1789),
.B(n_293),
.C(n_291),
.D(n_292),
.Y(n_1842)
);

BUFx2_ASAP7_75t_L g1843 ( 
.A(n_1768),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1787),
.B(n_292),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1837),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_1845)
);

NAND4xp75_ASAP7_75t_L g1846 ( 
.A(n_1765),
.B(n_1812),
.C(n_1808),
.D(n_1769),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1822),
.Y(n_1847)
);

NAND2x1p5_ASAP7_75t_L g1848 ( 
.A(n_1835),
.B(n_1786),
.Y(n_1848)
);

NAND4xp75_ASAP7_75t_L g1849 ( 
.A(n_1833),
.B(n_298),
.C(n_295),
.D(n_297),
.Y(n_1849)
);

NAND4xp75_ASAP7_75t_L g1850 ( 
.A(n_1774),
.B(n_300),
.C(n_298),
.D(n_299),
.Y(n_1850)
);

INVx2_ASAP7_75t_SL g1851 ( 
.A(n_1785),
.Y(n_1851)
);

XNOR2x2_ASAP7_75t_L g1852 ( 
.A(n_1834),
.B(n_300),
.Y(n_1852)
);

INVx2_ASAP7_75t_SL g1853 ( 
.A(n_1829),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1764),
.B(n_301),
.Y(n_1854)
);

XNOR2xp5_ASAP7_75t_L g1855 ( 
.A(n_1838),
.B(n_301),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1830),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1807),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1836),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1763),
.B(n_303),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1761),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1816),
.B(n_305),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1832),
.B(n_306),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1776),
.B(n_307),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1772),
.Y(n_1864)
);

XOR2x2_ASAP7_75t_L g1865 ( 
.A(n_1780),
.B(n_307),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1784),
.Y(n_1866)
);

XNOR2xp5_ASAP7_75t_L g1867 ( 
.A(n_1790),
.B(n_308),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1771),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1804),
.Y(n_1869)
);

NAND4xp75_ASAP7_75t_SL g1870 ( 
.A(n_1796),
.B(n_312),
.C(n_309),
.D(n_311),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1815),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1798),
.Y(n_1872)
);

NAND4xp75_ASAP7_75t_SL g1873 ( 
.A(n_1783),
.B(n_314),
.C(n_312),
.D(n_313),
.Y(n_1873)
);

INVx2_ASAP7_75t_SL g1874 ( 
.A(n_1782),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1825),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1826),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1791),
.B(n_313),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1820),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1821),
.B(n_314),
.Y(n_1879)
);

OAI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1795),
.A2(n_317),
.B1(n_315),
.B2(n_316),
.Y(n_1880)
);

NAND4xp75_ASAP7_75t_L g1881 ( 
.A(n_1766),
.B(n_317),
.C(n_315),
.D(n_316),
.Y(n_1881)
);

AND2x4_ASAP7_75t_L g1882 ( 
.A(n_1792),
.B(n_318),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1793),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1799),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1806),
.A2(n_319),
.B(n_320),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1781),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1805),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1794),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1810),
.A2(n_324),
.B1(n_321),
.B2(n_323),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1819),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1802),
.B(n_1797),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1788),
.B(n_1827),
.Y(n_1892)
);

NAND4xp75_ASAP7_75t_L g1893 ( 
.A(n_1813),
.B(n_326),
.C(n_324),
.D(n_325),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1777),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1824),
.Y(n_1895)
);

XNOR2xp5_ASAP7_75t_L g1896 ( 
.A(n_1803),
.B(n_327),
.Y(n_1896)
);

NOR3xp33_ASAP7_75t_L g1897 ( 
.A(n_1814),
.B(n_1817),
.C(n_1801),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1828),
.Y(n_1898)
);

NOR2x1_ASAP7_75t_L g1899 ( 
.A(n_1811),
.B(n_328),
.Y(n_1899)
);

NAND4xp75_ASAP7_75t_SL g1900 ( 
.A(n_1800),
.B(n_330),
.C(n_328),
.D(n_329),
.Y(n_1900)
);

INVx3_ASAP7_75t_L g1901 ( 
.A(n_1767),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1809),
.B(n_329),
.Y(n_1902)
);

NAND4xp75_ASAP7_75t_L g1903 ( 
.A(n_1823),
.B(n_332),
.C(n_330),
.D(n_331),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1770),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1770),
.Y(n_1905)
);

XOR2x2_ASAP7_75t_L g1906 ( 
.A(n_1831),
.B(n_333),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1770),
.Y(n_1907)
);

XNOR2xp5_ASAP7_75t_L g1908 ( 
.A(n_1831),
.B(n_334),
.Y(n_1908)
);

XNOR2xp5_ASAP7_75t_L g1909 ( 
.A(n_1831),
.B(n_336),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1770),
.Y(n_1910)
);

XOR2x2_ASAP7_75t_L g1911 ( 
.A(n_1831),
.B(n_336),
.Y(n_1911)
);

NAND4xp75_ASAP7_75t_L g1912 ( 
.A(n_1765),
.B(n_339),
.C(n_337),
.D(n_338),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1773),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1775),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1762),
.B(n_338),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1770),
.B(n_339),
.Y(n_1916)
);

NOR4xp25_ASAP7_75t_L g1917 ( 
.A(n_1779),
.B(n_342),
.C(n_340),
.D(n_341),
.Y(n_1917)
);

XOR2x2_ASAP7_75t_L g1918 ( 
.A(n_1831),
.B(n_341),
.Y(n_1918)
);

NAND4xp75_ASAP7_75t_SL g1919 ( 
.A(n_1774),
.B(n_345),
.C(n_343),
.D(n_344),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1847),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_R g1921 ( 
.A(n_1877),
.B(n_343),
.Y(n_1921)
);

XOR2x2_ASAP7_75t_L g1922 ( 
.A(n_1840),
.B(n_344),
.Y(n_1922)
);

XNOR2x2_ASAP7_75t_L g1923 ( 
.A(n_1906),
.B(n_346),
.Y(n_1923)
);

XOR2x2_ASAP7_75t_L g1924 ( 
.A(n_1911),
.B(n_346),
.Y(n_1924)
);

INVx4_ASAP7_75t_L g1925 ( 
.A(n_1915),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1869),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1913),
.Y(n_1927)
);

CKINVDCx8_ASAP7_75t_R g1928 ( 
.A(n_1882),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1878),
.B(n_347),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1857),
.Y(n_1930)
);

XOR2x2_ASAP7_75t_L g1931 ( 
.A(n_1918),
.B(n_347),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1875),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1848),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1839),
.B(n_349),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1890),
.Y(n_1935)
);

XOR2xp5_ASAP7_75t_L g1936 ( 
.A(n_1908),
.B(n_350),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1904),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1864),
.Y(n_1938)
);

XOR2x2_ASAP7_75t_L g1939 ( 
.A(n_1908),
.B(n_1909),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1905),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1907),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1910),
.Y(n_1942)
);

INVxp67_ASAP7_75t_L g1943 ( 
.A(n_1895),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1876),
.Y(n_1944)
);

XOR2x2_ASAP7_75t_L g1945 ( 
.A(n_1855),
.B(n_351),
.Y(n_1945)
);

XNOR2x1_ASAP7_75t_L g1946 ( 
.A(n_1865),
.B(n_352),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1843),
.B(n_353),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1856),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1871),
.B(n_354),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1884),
.Y(n_1950)
);

XOR2x2_ASAP7_75t_L g1951 ( 
.A(n_1899),
.B(n_1852),
.Y(n_1951)
);

XNOR2xp5_ASAP7_75t_L g1952 ( 
.A(n_1867),
.B(n_355),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1866),
.B(n_355),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1851),
.B(n_1853),
.Y(n_1954)
);

INVxp67_ASAP7_75t_L g1955 ( 
.A(n_1886),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1861),
.Y(n_1956)
);

XNOR2x1_ASAP7_75t_L g1957 ( 
.A(n_1863),
.B(n_357),
.Y(n_1957)
);

XNOR2xp5_ASAP7_75t_L g1958 ( 
.A(n_1854),
.B(n_357),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1888),
.Y(n_1959)
);

OA22x2_ASAP7_75t_L g1960 ( 
.A1(n_1898),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_1960)
);

XNOR2x2_ASAP7_75t_L g1961 ( 
.A(n_1846),
.B(n_360),
.Y(n_1961)
);

XNOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1896),
.B(n_361),
.Y(n_1962)
);

XOR2x2_ASAP7_75t_L g1963 ( 
.A(n_1879),
.B(n_362),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1883),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1858),
.B(n_363),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1874),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1862),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1842),
.B(n_363),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1844),
.Y(n_1969)
);

XNOR2xp5_ASAP7_75t_L g1970 ( 
.A(n_1873),
.B(n_364),
.Y(n_1970)
);

INVxp67_ASAP7_75t_L g1971 ( 
.A(n_1916),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1914),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1897),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_1973)
);

XOR2x2_ASAP7_75t_L g1974 ( 
.A(n_1850),
.B(n_366),
.Y(n_1974)
);

XOR2x2_ASAP7_75t_L g1975 ( 
.A(n_1849),
.B(n_368),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1841),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1859),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1901),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1892),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1891),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1887),
.Y(n_1981)
);

INVx1_ASAP7_75t_SL g1982 ( 
.A(n_1919),
.Y(n_1982)
);

AO22x2_ASAP7_75t_L g1983 ( 
.A1(n_1845),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.Y(n_1983)
);

INVxp67_ASAP7_75t_L g1984 ( 
.A(n_1912),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1868),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1917),
.B(n_370),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1885),
.B(n_371),
.Y(n_1987)
);

INVxp67_ASAP7_75t_L g1988 ( 
.A(n_1889),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1902),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1870),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1880),
.B(n_372),
.Y(n_1991)
);

CKINVDCx16_ASAP7_75t_R g1992 ( 
.A(n_1894),
.Y(n_1992)
);

CKINVDCx16_ASAP7_75t_R g1993 ( 
.A(n_1900),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1881),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1903),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1893),
.Y(n_1996)
);

XOR2xp5_ASAP7_75t_L g1997 ( 
.A(n_1860),
.B(n_372),
.Y(n_1997)
);

AO22x2_ASAP7_75t_L g1998 ( 
.A1(n_1872),
.A2(n_376),
.B1(n_373),
.B2(n_375),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1899),
.A2(n_376),
.B1(n_373),
.B2(n_375),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1847),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1847),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1913),
.Y(n_2002)
);

NOR2x1_ASAP7_75t_R g2003 ( 
.A(n_1877),
.B(n_378),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1847),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1938),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_SL g2006 ( 
.A1(n_1992),
.A2(n_1961),
.B1(n_1978),
.B2(n_1960),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1944),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1930),
.Y(n_2008)
);

OA22x2_ASAP7_75t_L g2009 ( 
.A1(n_1935),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_2009)
);

OAI22x1_ASAP7_75t_L g2010 ( 
.A1(n_1943),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1981),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1932),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1937),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1940),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1941),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1942),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1951),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_2017)
);

OA22x2_ASAP7_75t_L g2018 ( 
.A1(n_1933),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_2018)
);

XNOR2x1_ASAP7_75t_L g2019 ( 
.A(n_1923),
.B(n_391),
.Y(n_2019)
);

OA22x2_ASAP7_75t_L g2020 ( 
.A1(n_1980),
.A2(n_1959),
.B1(n_1955),
.B2(n_1979),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1964),
.Y(n_2021)
);

OA22x2_ASAP7_75t_L g2022 ( 
.A1(n_1956),
.A2(n_395),
.B1(n_392),
.B2(n_394),
.Y(n_2022)
);

XNOR2xp5_ASAP7_75t_L g2023 ( 
.A(n_1939),
.B(n_1922),
.Y(n_2023)
);

XNOR2x1_ASAP7_75t_L g2024 ( 
.A(n_1924),
.B(n_398),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1926),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1967),
.Y(n_2026)
);

OA22x2_ASAP7_75t_L g2027 ( 
.A1(n_1988),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_1957),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1950),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1954),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1920),
.Y(n_2031)
);

XNOR2xp5_ASAP7_75t_L g2032 ( 
.A(n_1931),
.B(n_1945),
.Y(n_2032)
);

INVx1_ASAP7_75t_SL g2033 ( 
.A(n_1969),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2000),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2001),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2004),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1927),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1977),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1985),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_2039)
);

OA22x2_ASAP7_75t_L g2040 ( 
.A1(n_1999),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_2040)
);

OA22x2_ASAP7_75t_L g2041 ( 
.A1(n_1952),
.A2(n_1958),
.B1(n_1989),
.B2(n_1936),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1968),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_2042)
);

INVx5_ASAP7_75t_L g2043 ( 
.A(n_1974),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1966),
.Y(n_2044)
);

OA22x2_ASAP7_75t_L g2045 ( 
.A1(n_1971),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1948),
.Y(n_2046)
);

INVxp67_ASAP7_75t_L g2047 ( 
.A(n_2003),
.Y(n_2047)
);

BUFx3_ASAP7_75t_L g2048 ( 
.A(n_1928),
.Y(n_2048)
);

XNOR2x2_ASAP7_75t_L g2049 ( 
.A(n_1963),
.B(n_415),
.Y(n_2049)
);

AO22x2_ASAP7_75t_L g2050 ( 
.A1(n_1946),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_2050)
);

INVx2_ASAP7_75t_SL g2051 ( 
.A(n_1947),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1949),
.Y(n_2052)
);

OA22x2_ASAP7_75t_L g2053 ( 
.A1(n_1994),
.A2(n_1996),
.B1(n_1973),
.B2(n_1984),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1934),
.B(n_418),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1953),
.Y(n_2055)
);

OA22x2_ASAP7_75t_L g2056 ( 
.A1(n_1995),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_2056)
);

OA22x2_ASAP7_75t_L g2057 ( 
.A1(n_1929),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1965),
.Y(n_2058)
);

XOR2x2_ASAP7_75t_L g2059 ( 
.A(n_1962),
.B(n_423),
.Y(n_2059)
);

XOR2x2_ASAP7_75t_L g2060 ( 
.A(n_1975),
.B(n_424),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1998),
.Y(n_2061)
);

OA22x2_ASAP7_75t_L g2062 ( 
.A1(n_1986),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1998),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1983),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_2064)
);

OA22x2_ASAP7_75t_L g2065 ( 
.A1(n_1991),
.A2(n_1997),
.B1(n_1987),
.B2(n_1990),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1972),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1983),
.Y(n_2067)
);

XNOR2xp5_ASAP7_75t_L g2068 ( 
.A(n_1970),
.B(n_428),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1982),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1976),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1938),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1938),
.Y(n_2072)
);

INVx3_ASAP7_75t_SL g2073 ( 
.A(n_1963),
.Y(n_2073)
);

INVx4_ASAP7_75t_L g2074 ( 
.A(n_1947),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1981),
.Y(n_2075)
);

INVxp67_ASAP7_75t_L g2076 ( 
.A(n_1961),
.Y(n_2076)
);

OAI22x1_ASAP7_75t_L g2077 ( 
.A1(n_1978),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_2077)
);

OA22x2_ASAP7_75t_L g2078 ( 
.A1(n_1978),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_2078)
);

OA22x2_ASAP7_75t_L g2079 ( 
.A1(n_1978),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1938),
.Y(n_2080)
);

OAI22x1_ASAP7_75t_SL g2081 ( 
.A1(n_1976),
.A2(n_439),
.B1(n_436),
.B2(n_438),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_1961),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_1992),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_2083)
);

OA22x2_ASAP7_75t_L g2084 ( 
.A1(n_1978),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1981),
.Y(n_2085)
);

OA22x2_ASAP7_75t_L g2086 ( 
.A1(n_1978),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1976),
.B(n_446),
.Y(n_2087)
);

XOR2x2_ASAP7_75t_L g2088 ( 
.A(n_1923),
.B(n_447),
.Y(n_2088)
);

INVxp67_ASAP7_75t_L g2089 ( 
.A(n_1961),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1928),
.Y(n_2090)
);

INVx2_ASAP7_75t_SL g2091 ( 
.A(n_1925),
.Y(n_2091)
);

INVxp33_ASAP7_75t_SL g2092 ( 
.A(n_1921),
.Y(n_2092)
);

INVxp67_ASAP7_75t_R g2093 ( 
.A(n_1947),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_2002),
.Y(n_2094)
);

INVxp33_ASAP7_75t_L g2095 ( 
.A(n_1921),
.Y(n_2095)
);

AO22x2_ASAP7_75t_L g2096 ( 
.A1(n_1978),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_2096)
);

AO22x2_ASAP7_75t_L g2097 ( 
.A1(n_1978),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_2097)
);

AO22x2_ASAP7_75t_L g2098 ( 
.A1(n_1978),
.A2(n_453),
.B1(n_450),
.B2(n_451),
.Y(n_2098)
);

INVxp67_ASAP7_75t_L g2099 ( 
.A(n_1961),
.Y(n_2099)
);

OA22x2_ASAP7_75t_L g2100 ( 
.A1(n_1978),
.A2(n_454),
.B1(n_451),
.B2(n_453),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1992),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_2101)
);

OAI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1935),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1938),
.Y(n_2103)
);

XNOR2x2_ASAP7_75t_L g2104 ( 
.A(n_1951),
.B(n_457),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_1961),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1938),
.Y(n_2106)
);

AOI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_1992),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_2107)
);

AOI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_1992),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.Y(n_2108)
);

XNOR2x1_ASAP7_75t_L g2109 ( 
.A(n_1923),
.B(n_462),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1981),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2002),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1981),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1938),
.Y(n_2113)
);

BUFx2_ASAP7_75t_SL g2114 ( 
.A(n_1928),
.Y(n_2114)
);

OA22x2_ASAP7_75t_L g2115 ( 
.A1(n_1978),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1981),
.Y(n_2116)
);

OA22x2_ASAP7_75t_L g2117 ( 
.A1(n_1978),
.A2(n_470),
.B1(n_467),
.B2(n_469),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1938),
.Y(n_2118)
);

INVxp33_ASAP7_75t_SL g2119 ( 
.A(n_1921),
.Y(n_2119)
);

BUFx3_ASAP7_75t_L g2120 ( 
.A(n_1928),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1981),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1938),
.Y(n_2122)
);

AOI22x1_ASAP7_75t_L g2123 ( 
.A1(n_1993),
.A2(n_474),
.B1(n_471),
.B2(n_473),
.Y(n_2123)
);

XOR2xp5_ASAP7_75t_L g2124 ( 
.A(n_1939),
.B(n_475),
.Y(n_2124)
);

OA22x2_ASAP7_75t_L g2125 ( 
.A1(n_1978),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_1935),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1938),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1981),
.Y(n_2128)
);

OA22x2_ASAP7_75t_L g2129 ( 
.A1(n_1978),
.A2(n_487),
.B1(n_483),
.B2(n_486),
.Y(n_2129)
);

AOI322xp5_ASAP7_75t_L g2130 ( 
.A1(n_2006),
.A2(n_2099),
.A3(n_2076),
.B1(n_2105),
.B2(n_2089),
.C1(n_2082),
.C2(n_2028),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2026),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2038),
.Y(n_2132)
);

INVx1_ASAP7_75t_SL g2133 ( 
.A(n_2114),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2007),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2048),
.Y(n_2135)
);

INVx2_ASAP7_75t_SL g2136 ( 
.A(n_2090),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2008),
.Y(n_2137)
);

OAI322xp33_ASAP7_75t_L g2138 ( 
.A1(n_2104),
.A2(n_496),
.A3(n_494),
.B1(n_491),
.B2(n_488),
.C1(n_489),
.C2(n_492),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2120),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2051),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2011),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2013),
.Y(n_2142)
);

HB1xp67_ASAP7_75t_L g2143 ( 
.A(n_2094),
.Y(n_2143)
);

XOR2x2_ASAP7_75t_L g2144 ( 
.A(n_2023),
.B(n_2032),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2014),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2015),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2016),
.Y(n_2147)
);

INVxp67_ASAP7_75t_L g2148 ( 
.A(n_2069),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2075),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_2111),
.Y(n_2150)
);

AOI22xp5_ASAP7_75t_SL g2151 ( 
.A1(n_2092),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.Y(n_2151)
);

BUFx2_ASAP7_75t_R g2152 ( 
.A(n_2070),
.Y(n_2152)
);

OAI322xp33_ASAP7_75t_L g2153 ( 
.A1(n_2020),
.A2(n_508),
.A3(n_506),
.B1(n_504),
.B2(n_501),
.C1(n_502),
.C2(n_505),
.Y(n_2153)
);

INVx1_ASAP7_75t_SL g2154 ( 
.A(n_2073),
.Y(n_2154)
);

INVx3_ASAP7_75t_L g2155 ( 
.A(n_2074),
.Y(n_2155)
);

INVx2_ASAP7_75t_SL g2156 ( 
.A(n_2091),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_2044),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2025),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2021),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2085),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2037),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2031),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2034),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2110),
.Y(n_2164)
);

INVx8_ASAP7_75t_L g2165 ( 
.A(n_2043),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2035),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2036),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_2119),
.Y(n_2168)
);

CKINVDCx20_ASAP7_75t_R g2169 ( 
.A(n_2059),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2029),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2067),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2112),
.Y(n_2172)
);

XOR2x2_ASAP7_75t_L g2173 ( 
.A(n_2049),
.B(n_510),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_2088),
.Y(n_2174)
);

HB1xp67_ASAP7_75t_L g2175 ( 
.A(n_2033),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2066),
.Y(n_2176)
);

OA22x2_ASAP7_75t_L g2177 ( 
.A1(n_2017),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2005),
.Y(n_2178)
);

AOI322xp5_ASAP7_75t_L g2179 ( 
.A1(n_2042),
.A2(n_515),
.A3(n_516),
.B1(n_517),
.B2(n_519),
.C1(n_520),
.C2(n_521),
.Y(n_2179)
);

OAI322xp33_ASAP7_75t_L g2180 ( 
.A1(n_2053),
.A2(n_524),
.A3(n_527),
.B1(n_528),
.B2(n_530),
.C1(n_531),
.C2(n_533),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2071),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2072),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2116),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2080),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2121),
.Y(n_2185)
);

OAI322xp33_ASAP7_75t_L g2186 ( 
.A1(n_2019),
.A2(n_2109),
.A3(n_2062),
.B1(n_2009),
.B2(n_2079),
.C1(n_2084),
.C2(n_2078),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2103),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2106),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2113),
.Y(n_2189)
);

INVx1_ASAP7_75t_SL g2190 ( 
.A(n_2024),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2118),
.Y(n_2191)
);

INVx1_ASAP7_75t_SL g2192 ( 
.A(n_2081),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2122),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2127),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2046),
.Y(n_2195)
);

HB1xp67_ASAP7_75t_L g2196 ( 
.A(n_2030),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2055),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2058),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2052),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2061),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2063),
.Y(n_2201)
);

INVxp33_ASAP7_75t_L g2202 ( 
.A(n_2124),
.Y(n_2202)
);

INVxp67_ASAP7_75t_SL g2203 ( 
.A(n_2041),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2096),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2097),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2097),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2128),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2098),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2012),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2098),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2056),
.A2(n_541),
.B1(n_536),
.B2(n_537),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2022),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2064),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_2095),
.B(n_2043),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_2060),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2018),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2054),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_2068),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2086),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2100),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2065),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2115),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2117),
.Y(n_2223)
);

NAND4xp75_ASAP7_75t_L g2224 ( 
.A(n_2221),
.B(n_2101),
.C(n_2107),
.D(n_2083),
.Y(n_2224)
);

OA22x2_ASAP7_75t_L g2225 ( 
.A1(n_2203),
.A2(n_2108),
.B1(n_2010),
.B2(n_2047),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2175),
.B(n_2077),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2143),
.Y(n_2227)
);

A2O1A1Ixp33_ASAP7_75t_SL g2228 ( 
.A1(n_2214),
.A2(n_2126),
.B(n_2102),
.C(n_2087),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2136),
.Y(n_2229)
);

BUFx4f_ASAP7_75t_SL g2230 ( 
.A(n_2133),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2169),
.A2(n_2050),
.B1(n_2040),
.B2(n_2027),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2150),
.Y(n_2232)
);

CKINVDCx14_ASAP7_75t_R g2233 ( 
.A(n_2218),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2171),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2157),
.Y(n_2235)
);

AOI22xp33_ASAP7_75t_L g2236 ( 
.A1(n_2222),
.A2(n_2129),
.B1(n_2045),
.B2(n_2125),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2200),
.Y(n_2237)
);

AOI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_2211),
.A2(n_2057),
.B1(n_2039),
.B2(n_2093),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2201),
.Y(n_2239)
);

AOI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_2219),
.A2(n_2123),
.B1(n_549),
.B2(n_547),
.Y(n_2240)
);

AOI221xp5_ASAP7_75t_L g2241 ( 
.A1(n_2186),
.A2(n_551),
.B1(n_548),
.B2(n_550),
.C(n_552),
.Y(n_2241)
);

HB1xp67_ASAP7_75t_L g2242 ( 
.A(n_2148),
.Y(n_2242)
);

AOI311xp33_ASAP7_75t_L g2243 ( 
.A1(n_2178),
.A2(n_557),
.A3(n_555),
.B(n_556),
.C(n_558),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2197),
.Y(n_2244)
);

NOR2x1_ASAP7_75t_L g2245 ( 
.A(n_2135),
.B(n_559),
.Y(n_2245)
);

A2O1A1Ixp33_ASAP7_75t_L g2246 ( 
.A1(n_2130),
.A2(n_562),
.B(n_560),
.C(n_561),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2139),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2220),
.A2(n_566),
.B1(n_564),
.B2(n_565),
.Y(n_2248)
);

NAND4xp25_ASAP7_75t_L g2249 ( 
.A(n_2168),
.B(n_570),
.C(n_568),
.D(n_569),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2134),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2137),
.Y(n_2251)
);

AOI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_2223),
.A2(n_580),
.B1(n_574),
.B2(n_575),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2142),
.Y(n_2253)
);

AOI221xp5_ASAP7_75t_L g2254 ( 
.A1(n_2204),
.A2(n_2208),
.B1(n_2210),
.B2(n_2206),
.C(n_2205),
.Y(n_2254)
);

AO22x1_ASAP7_75t_L g2255 ( 
.A1(n_2174),
.A2(n_585),
.B1(n_583),
.B2(n_584),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2145),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2212),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2146),
.Y(n_2258)
);

AOI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_2216),
.A2(n_2213),
.B1(n_2144),
.B2(n_2174),
.Y(n_2259)
);

OA22x2_ASAP7_75t_L g2260 ( 
.A1(n_2154),
.A2(n_593),
.B1(n_590),
.B2(n_592),
.Y(n_2260)
);

INVx1_ASAP7_75t_SL g2261 ( 
.A(n_2152),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2147),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2158),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2177),
.A2(n_603),
.B1(n_600),
.B2(n_601),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2159),
.Y(n_2265)
);

INVxp67_ASAP7_75t_SL g2266 ( 
.A(n_2155),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2199),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2198),
.Y(n_2268)
);

A2O1A1Ixp33_ASAP7_75t_L g2269 ( 
.A1(n_2246),
.A2(n_2241),
.B(n_2231),
.C(n_2238),
.Y(n_2269)
);

HB1xp67_ASAP7_75t_L g2270 ( 
.A(n_2229),
.Y(n_2270)
);

AOI221xp5_ASAP7_75t_L g2271 ( 
.A1(n_2254),
.A2(n_2165),
.B1(n_2190),
.B2(n_2192),
.C(n_2196),
.Y(n_2271)
);

INVx2_ASAP7_75t_SL g2272 ( 
.A(n_2230),
.Y(n_2272)
);

AOI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2225),
.A2(n_2173),
.B1(n_2215),
.B2(n_2202),
.Y(n_2273)
);

AOI22x1_ASAP7_75t_SL g2274 ( 
.A1(n_2261),
.A2(n_2140),
.B1(n_2217),
.B2(n_2165),
.Y(n_2274)
);

INVxp33_ASAP7_75t_SL g2275 ( 
.A(n_2242),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2227),
.Y(n_2276)
);

OA22x2_ASAP7_75t_L g2277 ( 
.A1(n_2259),
.A2(n_2156),
.B1(n_2182),
.B2(n_2181),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2232),
.Y(n_2278)
);

AOI22x1_ASAP7_75t_SL g2279 ( 
.A1(n_2266),
.A2(n_2132),
.B1(n_2131),
.B2(n_2184),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2235),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2234),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2237),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2226),
.A2(n_2188),
.B1(n_2189),
.B2(n_2187),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2239),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2250),
.Y(n_2285)
);

O2A1O1Ixp33_ASAP7_75t_L g2286 ( 
.A1(n_2228),
.A2(n_2138),
.B(n_2153),
.C(n_2180),
.Y(n_2286)
);

NOR4xp25_ASAP7_75t_L g2287 ( 
.A(n_2247),
.B(n_2193),
.C(n_2194),
.D(n_2191),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2251),
.Y(n_2288)
);

AO22x2_ASAP7_75t_L g2289 ( 
.A1(n_2224),
.A2(n_2162),
.B1(n_2163),
.B2(n_2161),
.Y(n_2289)
);

OAI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_2236),
.A2(n_2167),
.B1(n_2170),
.B2(n_2166),
.Y(n_2290)
);

AOI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2240),
.A2(n_2149),
.B1(n_2160),
.B2(n_2141),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2233),
.Y(n_2292)
);

A2O1A1Ixp33_ASAP7_75t_L g2293 ( 
.A1(n_2245),
.A2(n_2151),
.B(n_2179),
.C(n_2176),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2270),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2289),
.A2(n_2264),
.B1(n_2260),
.B2(n_2249),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2276),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2272),
.Y(n_2297)
);

NOR2x1_ASAP7_75t_L g2298 ( 
.A(n_2278),
.B(n_2253),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2280),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2281),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2292),
.B(n_2244),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2282),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2273),
.A2(n_2252),
.B1(n_2248),
.B2(n_2257),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2284),
.Y(n_2304)
);

AOI221xp5_ASAP7_75t_L g2305 ( 
.A1(n_2290),
.A2(n_2268),
.B1(n_2267),
.B2(n_2256),
.C(n_2263),
.Y(n_2305)
);

AOI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2291),
.A2(n_2172),
.B1(n_2183),
.B2(n_2164),
.Y(n_2306)
);

NOR2x1_ASAP7_75t_L g2307 ( 
.A(n_2285),
.B(n_2258),
.Y(n_2307)
);

AOI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_2277),
.A2(n_2185),
.B1(n_2209),
.B2(n_2207),
.Y(n_2308)
);

INVxp67_ASAP7_75t_SL g2309 ( 
.A(n_2275),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2288),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2309),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2294),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2301),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2298),
.Y(n_2314)
);

AOI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2295),
.A2(n_2271),
.B1(n_2269),
.B2(n_2293),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2307),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2297),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2296),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2299),
.Y(n_2319)
);

AND4x1_ASAP7_75t_L g2320 ( 
.A(n_2317),
.B(n_2286),
.C(n_2287),
.D(n_2305),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2313),
.Y(n_2321)
);

AND4x1_ASAP7_75t_L g2322 ( 
.A(n_2311),
.B(n_2243),
.C(n_2302),
.D(n_2300),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2312),
.Y(n_2323)
);

INVx2_ASAP7_75t_SL g2324 ( 
.A(n_2314),
.Y(n_2324)
);

AND4x1_ASAP7_75t_L g2325 ( 
.A(n_2315),
.B(n_2310),
.C(n_2304),
.D(n_2303),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2316),
.Y(n_2326)
);

AO22x2_ASAP7_75t_L g2327 ( 
.A1(n_2318),
.A2(n_2279),
.B1(n_2274),
.B2(n_2283),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2322),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2321),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2326),
.Y(n_2330)
);

NOR2xp67_ASAP7_75t_L g2331 ( 
.A(n_2324),
.B(n_2323),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2325),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2320),
.Y(n_2333)
);

CKINVDCx20_ASAP7_75t_R g2334 ( 
.A(n_2332),
.Y(n_2334)
);

INVx1_ASAP7_75t_SL g2335 ( 
.A(n_2330),
.Y(n_2335)
);

BUFx2_ASAP7_75t_L g2336 ( 
.A(n_2329),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2336),
.Y(n_2337)
);

OAI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2337),
.A2(n_2335),
.B1(n_2333),
.B2(n_2334),
.Y(n_2338)
);

BUFx3_ASAP7_75t_L g2339 ( 
.A(n_2338),
.Y(n_2339)
);

OAI22xp33_ASAP7_75t_L g2340 ( 
.A1(n_2339),
.A2(n_2328),
.B1(n_2331),
.B2(n_2319),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2340),
.Y(n_2341)
);

AOI221xp5_ASAP7_75t_L g2342 ( 
.A1(n_2341),
.A2(n_2327),
.B1(n_2308),
.B2(n_2265),
.C(n_2262),
.Y(n_2342)
);

AOI211xp5_ASAP7_75t_L g2343 ( 
.A1(n_2342),
.A2(n_2306),
.B(n_2195),
.C(n_2255),
.Y(n_2343)
);


endmodule