module fake_jpeg_24975_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_38),
.Y(n_65)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_59),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_31),
.B1(n_22),
.B2(n_33),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_56),
.B1(n_37),
.B2(n_18),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_31),
.B1(n_22),
.B2(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_25),
.C(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_66),
.Y(n_72)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_16),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_16),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_23),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_43),
.B1(n_45),
.B2(n_31),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_47),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_45),
.B1(n_43),
.B2(n_34),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_43),
.B1(n_34),
.B2(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_82),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_42),
.B1(n_41),
.B2(n_39),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_90),
.B1(n_52),
.B2(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_18),
.Y(n_109)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_89),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_41),
.B1(n_39),
.B2(n_36),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_109),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_59),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_108),
.B1(n_71),
.B2(n_74),
.Y(n_119)
);

XOR2x2_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_52),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_104),
.C(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_19),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_32),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_106),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_29),
.A3(n_25),
.B1(n_20),
.B2(n_32),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_20),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_47),
.B1(n_51),
.B2(n_53),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_18),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_86),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_122),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_121),
.B1(n_127),
.B2(n_130),
.Y(n_146)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_110),
.A2(n_75),
.B1(n_74),
.B2(n_80),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_70),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_80),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_109),
.C(n_114),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_85),
.B1(n_84),
.B2(n_73),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_85),
.B1(n_49),
.B2(n_84),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_76),
.B1(n_87),
.B2(n_28),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_103),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_49),
.B1(n_57),
.B2(n_81),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_96),
.B(n_115),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_160),
.B(n_133),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_99),
.C(n_94),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_157),
.C(n_29),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_141),
.B(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_144),
.B(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_95),
.B1(n_104),
.B2(n_92),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_161),
.Y(n_170)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_155),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_102),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_113),
.C(n_106),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_97),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_114),
.B(n_28),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_126),
.B1(n_128),
.B2(n_138),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_138),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_165),
.Y(n_184)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_168),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_119),
.A3(n_118),
.B1(n_127),
.B2(n_135),
.C1(n_134),
.C2(n_29),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_23),
.B1(n_24),
.B2(n_81),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_149),
.B1(n_160),
.B2(n_146),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_1),
.B(n_2),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_142),
.B1(n_4),
.B2(n_5),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_23),
.B1(n_24),
.B2(n_57),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_173),
.A2(n_174),
.B1(n_158),
.B2(n_161),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_24),
.B1(n_57),
.B2(n_55),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_175),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_55),
.B1(n_41),
.B2(n_27),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_142),
.B1(n_155),
.B2(n_55),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_185),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_195),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_178),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_186),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_196),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_144),
.C(n_147),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_191),
.C(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_148),
.C(n_163),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_3),
.B(n_5),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_27),
.C(n_21),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_14),
.C(n_4),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_8),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_176),
.C(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_195),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_179),
.B1(n_172),
.B2(n_166),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_203),
.A2(n_204),
.B1(n_194),
.B2(n_190),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_167),
.B1(n_174),
.B2(n_171),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_173),
.B1(n_5),
.B2(n_6),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_3),
.B(n_6),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_8),
.B(n_10),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_193),
.A2(n_3),
.B(n_6),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_219),
.B1(n_222),
.B2(n_212),
.Y(n_227)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_201),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_206),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_207),
.A2(n_191),
.B1(n_189),
.B2(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_205),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_227),
.B(n_203),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_202),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_230),
.C(n_210),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_205),
.C(n_202),
.Y(n_230)
);

AOI21x1_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_218),
.B(n_216),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_236),
.B(n_224),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_209),
.B1(n_207),
.B2(n_189),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_235),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_239),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_232),
.B1(n_236),
.B2(n_228),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_221),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_231),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_230),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_243),
.B(n_242),
.C(n_12),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_244),
.A2(n_245),
.B(n_12),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_241),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_13),
.Y(n_247)
);


endmodule