module fake_jpeg_9808_n_66 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_66);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_66;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_1),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_31),
.B1(n_5),
.B2(n_6),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_15),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_3),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_30),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_48),
.C(n_49),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_51),
.B(n_52),
.Y(n_57)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

FAx1_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_26),
.CI(n_16),
.CON(n_48),
.SN(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_4),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_4),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_18),
.C(n_23),
.Y(n_53)
);

XNOR2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_54),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_5),
.C(n_6),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_55),
.B1(n_48),
.B2(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_60),
.B(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_57),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_58),
.B1(n_56),
.B2(n_46),
.Y(n_63)
);

AOI322xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_58),
.A3(n_55),
.B1(n_45),
.B2(n_44),
.C1(n_47),
.C2(n_53),
.Y(n_64)
);

AOI322xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_44),
.A3(n_13),
.B1(n_14),
.B2(n_19),
.C1(n_21),
.C2(n_11),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_65),
.B(n_22),
.Y(n_66)
);


endmodule