module real_jpeg_14093_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_65),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_65),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_4),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_6),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_42),
.B1(n_83),
.B2(n_84),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_10),
.B(n_30),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_49),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_12),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_12),
.A2(n_34),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_40),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_13),
.A2(n_24),
.B(n_29),
.C(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_13),
.B(n_83),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_73),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_13),
.B(n_47),
.C(n_60),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_13),
.B(n_23),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_13),
.A2(n_50),
.B(n_131),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_73),
.Y(n_157)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_112),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_110),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_77),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_18),
.B(n_77),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_56),
.C(n_69),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_19),
.A2(n_20),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_38),
.C(n_44),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_28),
.B(n_32),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_22),
.A2(n_28),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_23),
.B(n_33),
.Y(n_158)
);

AO22x1_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_25),
.A2(n_26),
.B(n_73),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_26),
.A2(n_27),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_27),
.B(n_121),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_29),
.A2(n_42),
.A3(n_84),
.B1(n_87),
.B2(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_41),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_50),
.B1(n_53),
.B2(n_55),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_55),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_52),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_46),
.B(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_53),
.B1(n_55),
.B2(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_50),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_51),
.A2(n_52),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_52),
.B(n_76),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_55),
.A2(n_75),
.B(n_136),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_55),
.B(n_73),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_56),
.A2(n_69),
.B1(n_70),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_56),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_63),
.B(n_66),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_57),
.A2(n_66),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_68),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_58),
.A2(n_64),
.B1(n_67),
.B2(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_95),
.B(n_97),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_62),
.A2(n_97),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_62),
.B(n_73),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_71),
.B(n_74),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_84),
.B(n_86),
.C(n_88),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_99),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_90),
.B2(n_98),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_92),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_164),
.B(n_170),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_151),
.B(n_163),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_132),
.B(n_150),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_116),
.B(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_127),
.C(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_140),
.B(n_149),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_138),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_144),
.B(n_148),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_142),
.B(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_153),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_159),
.C(n_162),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_165),
.B(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);


endmodule